PK3  c w^S�S���'  � H  d5d9210ef49c6780016536b0863cc50f6de03f73e70c2af46cc3cff0e2bf9353.unknown�  AE ���P�Ӑ����>e��1���� P<ax8k䛜�,JF��K؜a,�E���`�����&Wr�O���{���H��ɀ�5˹�[�naH��h��ҪG�ӆ�=�[?���}Tt�^��k۝���Q�
{ �̸���/�zх�z�W�:�W��d@d+���7t�o���h����V�q��0֪)�"<C��^�vA>._M���,�8r%�������x&��`���@Z�}[��Ǝ8/�� �T�'�)��y�P�u���˟�ش��)ָ[����Ѐ������zB�VP���&��1sZ�ˇ�떊�Kݭ�Gd��v%�54��b�J�Q��OCNZM��`����G/�kmz��z��۸����&�pD���⠘կ[w(���D��J�2V����J.~��J��n�p��$^���~I�ώ���)�8�ځ;c�܀��n���e!�lH���@��6�2�a�H�31�bU��BA�K�N=�>��(��tX2���ŎKQ2���� ���+r�m�MV�s���E'��{��t}F/.2k�D�e���܎���b��;qs���{������Ա^z���G��C�ہQ�o.����I ���6�c��:zԸ���o���Ӏ��@�q{ʦk(��ITq@��/��v 䜟1[��ͬ�|�z�}T��@�7��F�=P��<���� X���,�(1X�L�7�z����V9/��S*�9�|c��)3�A�5E�Ij�K�I<����ReWB<��q��{�𦗲§,�ۋ�dA��a�7P���:)fFM�6�'>Q�#,O��y8��L��e��]p羒{)Uc��rJNQ��7\��OJEX�)ŰV!;��r�����Vx�Ma���i[�6֍;�L��:�]W-�U�*-�޷�{��4T�;��
q �=�D��W5=�e�2ՄzIM2��w\������btλ�v2čDGH�����e ||WՈ6��}5*.$�D=mH���_a{đЫ+�7����-E�e �jvS�3G���1�p.`6ڽ�wo��.hY�f�S��vzel�#�P�Y�QՊ/^)�m�SQ%%p�א���m%ZsQ#����o3t�ѫ�.z����,q����8Z��Z�S���	Ur�<g������`��V��5׷���v��#��A5���ٕx��0�qj�����[�z��S��W�k5\ Dw;�k:-ve���E�O��֋�}cx�\�r[�?�(q*�,�_�WӼ8��`�v��*����.:�O�����~��"6���7��B'xҶVH�j�=�Ŷ$��KJ7NFOE5������-�Y[�`��X���t���eH}�M ����B���(t;'���y<�XD-7o`.���j��f_L�逼R-�.���'�S�x2�����*˓^�y
�f���a�����9�F��D����:9m�)\���D�~B�o H��@
���gBCy����W��p�4�|��'2&'��lyESG��M[�_��I�	�M��gK�=�j>PF�{�mI;�^����~("�y���_>+ֳ;;�]iU�Z�� ���
��uE2�<�4e�m��lz�0;�3����{9�\���
W��P�H�Ej;ScW�r�bsu�;2�j�*���$�bh���Ͳ5���RoY��\I�%
�����&���)�r�'xݗu�ä������>2칮n�$[.�o˲�x/O9��H��p��JuY�"�
}�D���r��D4���Z��_�������:XT�~�1YG�N#��ɓ��]�Z��i]q���`S�Re�k#�д58�-Q]���6��dcT>��_�����C��No��A�~�E����9�/0��ũ�&x/͒<���	�-���s&.KZ��eq ��נ�_��]My�E�A�t�V,���ѣ�����rַ	�T0���W�<�p_�S������_ĸ�\(A?��Cty
�؇n.8�����y�x
�m=)H$w7/��Hr�pjZc���w� ~>����4�����:�@�a�9��z�(�yU����	� ���c�yW�����TM �'z��O�#�۞��av�C�f� ��?w�b�2����Cj2guHC�\��x�25S�g!�8�u�������׸h���šro��)S�K�����׊Z�fJmg���b�	r�{?���'&��7p���+��{m� oD8.�� KW �^8U�B�f�Ē��?3�`�}4U�7\�S~xz2��:x��6��b��Ql7{7��\h��'w�U{H[��By#1OwL�XH��O�d�Cy�pu��\
2,/�m���a���wޡE���̄k�/Ԡ��@��<Z��������M&�{��ΝT킞R��?���K���F��`�j(}ǒ��*�����ֱ'pjk-7��3<;���1�	��T��p��1K��^�F_C��.��D���6pL��J)��R� ��,�zH:+��4e1o�+�-C����M�{&K|�+A��,D~�0ms�����ƽ��R�v)�:�����I���gZ�e�L��)��(�I�-�b{�Ŝg;w�;���o�w����1N'F���V���枅��i�@�hV�����Y���s�;��=e%Q��Z��'`o�rK,� ^j1�
\&���L�&���
s�t$�O��Ⱦ�ADI3Z�1�����2|���z=�����ϦD���c�:�)}e΂i�|�D=T�n�`��%��}wV��a����C�)��X�L��Rۉ����;]K�먯�N%�v0 ���� <����dڕ4�mX����:�K��i��^��՞m/��,�KZ��[�ބi�!Ե���o��f��Q�o����?� �����ۇ26o z-|E�L9M�SͰ)&?��>�n�vcCJ�<�L@Gy��"��J���r��A��h��ȹ�b>��8���H�v��{QX#��|LZ;�O�*�]�!L@�z���� ��v��1Hfe�h�x���nPH�D�$��ژ�� cF��m�B&��"��h�̪���F�W�Э�Q��+G�A-�a�T��_�`�AE���Ծ[��`�&��`:W������ep�zd󺈬o���i �)+���m�����S�Z�͔]�pX����)�{7�N&d�3g�1[ʏ/VҼ޾J?�Dh������=[����S�:g�o����	���/)�������RG`��0�l�Q\��d���5 �f�'29nP��P�����+�9�%�Z��><�J.D���=��>���r-�����<^�l�N㒨�yz r��Wz2~���7Cb�����q��j\&�1�
䌌��!c ?�^�@��<���
��o��>9�TQFi}z���b�I5cM��C5��~��05�0��c�o�MZ��ܝS�Ko�C��~h�f���dÀiuR�!�E�~�D`��t�j65�	�A%�,�Ġ%�81׽�b�=]>����}U�>tad����L�Q���V�Eh�c�����C|���b��w��l˽��Փ�i}_�ޮ��n&l�1��5og��=��@��u@B}ga��\�(���׼Q�6NE4B@V�:^P�G���d� ��l�AK%ᦂӥ��=}Qi��B��zpfJ��tR�Èj^�<�78�ɯ "T-,��l�<�'�� ejOZ�;�c���*�]C����e��TQ3�xyrE#kj"O���� ��Hv0��|��41����D�d���һF%F �'Z8er�q��% ���<��I�1F�J; �M]H�Ӌ�Oc��F̱6#n��oNۑ��{�"�??H�O��"�!����C U=��&�!����u|�3��-��L
q�%{Δ6toE�>0~�oW�2t�P♷R:�Z2���`����K�O;�L�IL��M6a���`�k����̾F�g�4�۹	�yN�k���n�#BL^��\�:����O�0��F��Q��Ղ�g�A���!+�����UB�<#4�
�pt����읗���g%:ux����nR���P4ȧ����� zV`��f�+͛ӿeNF�BsBB=��2��2�w4��5�f������Z�`z&��R�(B�#�;������Z0�	�<����=Xݖ���5�N��Ap�� �O����85�&�<�fLx��3�ts�3�4��^��_�vϪ9�u�D� �e� Y����ȡcZB�?+�b�?�O�܅���"���I���?rp����Q�!B3�n��\�\+0�}��	�/Ƿ�^_>c�� �t��k��Hp#1���'�>��t�+�^�`M��Z� ��E�֒7�9mu1�n�4�&��վL10.2�[�s<�䋴�H{�?(J�B��CA���_}#*z'�s��k���-��J�֝h�r�0�T��o�V3>MV���M0c�6������E]�ot+�4?���B�ݫ{H�1>�Y����g]F�B�9E��W��C>�T�'}�,`�Ӡ����R�k��RwGp�fh����tm`qdd�b�݃t�#Q�2���L�7>LϏ�as���@�K��䖔j�=<����Ix&N����9����(�3@$���:�0�^ �h����m鹜��L�4�K��!����/w�%�wr��c�^�\�����b�'��!��χW3��c�����m�&M�<�j�孖^���FOM�n;Ȏ=��r��f^)�^(y����d���A uc"(�:���إ����f�8�I��~�4�R�1핗At��+�[�ݵ������ڭ����R)��ҾA� F�7y��MS?ׇ(��#A���y�|�;6@��;�2`���zq�w��j�U�[�]L;��0|���m�.��h�{X	U��j�.@U)���R֏r{b���7@h�0��
��	�H�C��MP��]�M��aae�,v~�<�B�n����/s��>���-j�l�kg`ݵ~g�]�� !�I��r8��2�grs�m����$��ԫ!��p_*e���V�l��o�2��-=�#���cپ�֌���8�̲V���5���Nʴ��S�M�֥@!����?87ek�l����L���*$�{����dvINؐ�&@|Z\�;[�J��8�����)���Mۧ)�10/�e���gi��o/�ݐ���(��_���4�0��N!=�/H��_>f��,�Z����E��u���Ҍ���jK�P(pȗ2���j�%_��Փ����X�y���K�~��Ngq�cd�Mo��Z>��K��Cu1� l��M�ܣ;�2�/��)�"/�ݩ���d_�A`|���is�e�靋�@v�a`%t��ދ�ڕ_Q��I��R<����?p.>�լ�|�;�H��M�lSKl������/��=�@:�ԤR���}�JBN�~󼰣{;���Y�Rx��ʉ�\ Ο+�����`	���J�55dI��[#@'S�8`�a�W��@�L�n�,M���wW�LД7A��^E�O�/}�c`�;����%g�p�̈́D�_[3�6��N�=�ˉr�p�Z��W(x8<\�W_|Y��.���6�⥫���|b�!���D�&?U�]�������6JT`��8�;x�=����o7>Vw�֦����Pa�Y���_4#�	�DgRw![�=ڂ����m����B�H����gN�M��'g9���(.�x>�a�����^���J�P;ZN�H7�ZUL�� �F��_�G�V5$����!:�:�6ⳛ(dH�k(���3K[9]���[J�u����*ֻ�;zX���b��䊍^YE��f@swV��g�t-���7o/�P��h��[xA�'Qǲޱ1I'��}
|��3fR���"{i_���vմ�.�۵��W=�À0![O5,�. z���� [��3A��9��;�zT�6F]l�;|���҆��bO��݄�LB��O
�X�����AC6-yZ~!�2{�\�w��[�ߤ�'������/ψ�B.a��0�;��i�Pl�,s��	�>�o�L�%w|iٚ�ed�����m��T�B�l̜��!%(��h�����W�Ǵ|����,���3���,A1o���/b��*����Kc"����2h k����.���_�ڣ��ӯ�w\d�v�M����2���oC��oQ��t�Q��{����;�y��8����bn
�֓�ߗ�2ո�eᩉ�եg�F3�1�7������l��_�X �ff{q��)t�ّ�Rw�G�-\\/2M�v���C�B]-�5D	*�G�T�Q�	��J.(�R[H-�(����8�Øx��K�o$�����ȧ(���T�4� %t�g`ۇ���t��W_�s����X���Ě�J��9a`�J��<I{����KC���5�I�u'���Fm����V7''�Kg�j�z�|�-� ^�&��уc/��d�i�$�?��ڽ��V���)G���K�k��..�Шd�9IOۆz�g�>{�~^������
��^�)���3�x�"��6��x�^����#Ad(�O��D��?}!P9n:��� �z�s-�J�^y�a�b��BN��=�����^v90��r���o1���{���b�O�-��A�S��QB�4}W2sr&������ht�[(��tw��,d7�� �\<g�~��ˤ��(�<PLt�Z:"I�����Z�L2�-�kA:�]��:�OS�,ZD(�G|Q�a�D�N��wUŶ���c$�,�����h���+?-��r�J`� � ?��'1��w��>�G�3�]eXh���Rwb�ŏk�c?����O�E |���B�����S�lYf9`gk�.��ڿ^���~'��'xU��c��U�唩O���Ď�q�'g��v�~�}�ϵ��6-���r5���J��(�����~����#l�CE"Q��}�4UX���k���uO�J��C�+�h6eVy�槩��=�.�p�ۍ�-)�8��O:MeG�HOk��}�S�]7���(�c�&�Ʉ �75C�ܽ���C=`GT
�s /*ʊ����B�''L6|7�w�Y�3����ޅw�����SM";-vn����j����'�L�]HќK+o�2v�h��\$  �O���Y.�$)��� ��3,�Pz�
�#��魑|�vP9r�'��l*ze��@d���(	�_�p�=k�9����y��3;/���`�2q�%���_Y�ﬤ��>:�%
��ެ���Kf�3����3�C�CZA=�@U_�)�6Ju��,����
i$�U)�P$ů��f[���� �ש�)�aEc����8o�`P�aK��4~EV�����a2��)Ձ梅s�Z&�'l_p�+ߌ|�;��m�͈ߨ��Že��fsٛCJU�i�z�8��Nw\L�������C���&J�.����JƗ����j��E��P�Ta���P�����SM˃�K��s��ʌsC�>/�,��Ǔ�� :nX����E$����rU�D\o�0isI<�yȺ����}�X��p���24�+��S���J�*�AJq��{�L:k���U�S(���~+�0��j�\1A�eM2��G	�B�r��=�1L[���j�{��B��Į�>�y��;4�Q3-+���a�q��r��j�����X=�E�P�	��������搈w��_�s��8d�F{L�=�����I:�^��f)�#��g�<0c(��S��h��v)d_T�1 ��&NW��R5�A+���7�s+���G�E�,Dں߸�mC:c9x��=��W�� ���¿�QWc��l�e�%��dV��4���9��x�������l>�B�Æ5�ι���F�hoJ�&f�lJ�9����C����o�w��,gx�YR?`_.ۭҙ�vl�pHYt���>��hZ&�Tx�5���Ű�盱��[vGϏ־K|�ի���������aƣ�M\�F.ryz$�=׿�<���j��n�����k�a�����������`���aT�*b܈���pS��^ZK�M��ŕ�0d�]��OIϔ��r�i��	�re�]hH��P���S�7�U	@I9u�����m1 �T���1����9uŝ��)?jrl�Uk?�f.'W�^������hp:���_�,g糢�Nf�w��T�uX2j�x�FAͦ��}��w��ce���p�����J�;��Z����:�dnD��P��!�^M�[B2�9��@�!��݁�x�/V����+N)	�0a�r�����-`ɫ^��ױ�"���B��G��K�ì��m��������kIb�܂�|.Z;2c׍���� ��y65Iz�R"q��w'�duD�6:�32�O�D��܀��Ŷ���/�!�G˖�-q>!���%r�M��%B�+����t�`�:�W*4tA[�:�X,t%;g��'j�������͖�?�ٙ��[�%��c����ҬaPL-쐻��D$\11���$�>c����*�hO+ִ �|;�#��'�6��uO|Զ��)W���\���%��٘])�Fvn��1e@��{�"aV�c�/�)����8/w��9�H��?�u�0���ץM~P͊?��Q�e0�&+r`eA�]��Ƭy�v	��)���A��J|�lX�$v��d����q,��B��Jn�u��H���s��ib�f/�A}��b̚3�g��+|[A�!�+�@��kl(��С�?���[���œy�j<�D��8�@s,�M�Qa�N	���1‴Q<FU[�c)6�^��>p�� ��ޡ@ri=��� �*����萉R�����t3پkHGYI�=/Q���<mr,�$n�M���%QXj���+�K��/�yN ���_S�X��)����vCd����)��Ap�V����Ol�f�v���*췁P��(�W�z�p��q��ߊ�q3Va��Ë�XG�/������-��t�!8�� �W5�_����z��(�.�v��ꏪaA+	3[o!��hHn�#e��W�Q
P��&����Ѷ�W*�<*Ŋ�1�2��te	���Y��eu<^T�л:0���M"�#��0������d]���l�Ǆf��z�J����V�w;~=ΰ��`����veԄ��E������k���w��4�F���.���9�7�3|��l�����Q?x�.���r<.C�Q��5%ݮD/����1���ɮ�E�@�*�f�����OpH3}��[�pm�&����v�D�@��2�������@��LXS�S~�������O7��+k����+}��"�d傈}!z˺&H#��ݝ�|�ԩ%�͈/������{�z��b����Ƴ#��w�Tý�5m��U�;��+�N��q*�.5�کA<�@UbY;*2i�.��ƚ8���J(���KВ���ͭ��k�qP�h���o�������	���z�����`dN��P_2[J!H����շF�q���k�sRtr7�1�js����:�n@W�2٨@��	��[�z
���?�y����O��ٽ2��!~L�/�����7xx7�&W����%i�kNڽ�QH͵h_�$"Vf@�ڂ0�2^2��wI(�����g4k�qcZ1Zp����!�u���wݞ�O2EL��>o5��R* �_���Iӿ�7m�$7��s��p�ơ�K���=�>��H2��,ʳ����}�a4����"M!ê�Λ�J�yZ�n���k�c��ϙ��qj��E�J��k�s�%�h�	��W5�+����G��1�ټ�~< ("C�����+�Y&� 7��>��	�|�Z*L4P��ZE�UY��>n��1��r�A�
��S`rn���� ��Ԥkl|g����sjð��Ѵ[��i�5���Q����ޛ��H �HX*aT��]s|'�޾~m��+l�I ��e�� .�_�H2X�{�'�O5u�M�f�B��_������g%�s�ϵ`�2	u���'Y����0}6ZE��X� �����A��y����-�S�o&�M��u/�[Y|��A�&fg�dQ
��+�%�F��`O^���~��y�2���:Q��՝���
���c

�]m��mB������i��Jm��"pT�q��6�%��p���OB�t �[�'��5�����I������Q�:o# H����;��_eg���D{����aϿ���������v�ɒх.��,Wd��(ҤJ�p����Օ�5���J���@��:+�����&��,���u ����, t|���1�,�������aN�*6I���tá��ʔ��+3|��W�A�F1r�����m/�i�v�iB&�>$�n�z��^��.G�X�o��Vڨ������0���lP��f_�Ѿ�-������'ǌ+y��;m�'J���O�toŧ����%8Q?����Lc�|S���#��v�L>'U�hi!�J~*��!��s@qݢ��XO�<��l8G{Wc��CC��jQ���cg"���W-�0�U��^l������g�hF��e��|��W�C��AYV@�����^Ρ�����W@͌���^AGߝ�P%o��0�&]�#�y���~.�"a-��m�)ċ6����[�#�
�o*�#��ȅCx�&@.M#��2սz3Xc���Џ3��{�$$�dX��l�7G'~�H�>�0�(� R�V�s��
@Ӟ�@�:c�4����⹫����A���x�-���e�\k�g9�z����3��m��IU�[Ԁ��M��K��� [G)٥�Gn���FV�I �ix�B#=��1'��GR#ǩQ��՘�G&��&y��n�Y�xKo���E���Ļu�)MC;%��+�_���Q,l���	�~��|�õ�UR֯��ց���>���/a_3�zQ�m��_̑d��2��Þ��YӵT�VM�:"�[(�:`��G�{ Ց��Ny��}���ٞ��J�֌��_�3)���p�?$��\BcXԚ�Shޖ�>l͇/����Q�T'��BYӾI=���-����C��b=t�����Kt�܈}�����͉rş�R�0�meʏ"�Ї�ȝ�Gɿ��1�ю��'�\m����nb�<��х��K�\�0?=j��.�����<v��P&*ǖ����1�K���9�S��7PF!�g�_sO�����|�j6�1�Ƚp�Rڕ�������i��N���K�㲗 �J��$VH(����n��>�~;�F.m��g6�O��*���B�:��qɎ�b,��͓ bf���(T�{<��.�$�����3T�caR4�� a� ��wS_e�p���!�G�:J�zQ$"ם,au�き?�h'�]�x�7q|WY?���2-Nt�)�Dujֳ��3���K�����]n|�:��%����>a� O@yUE��ԟ���e�d���I�;#-G�F���/�UM1)=fS�0%�W)c%I�_<�Vh: �`������8�Gcč~�kf��;mW��J�J��5��|Ĕ�q��>0d�(��7s"���暋�͢��h��ќ'и⁀������|'��1��n��c�:�꩙�Ya�h���8CL �މ+9v*��3��[*U��<@�P|��z�<�Z�(�>�����)�k��n;v�R���Br�R�&3�Z������ �v�1{�O�"b|O.���`��Ӌ��G�e�h�nY��T,v
,-��>��%��j4�Z�;����?m[��|�ܔ�rϚZԛ�w�� ��B!��6��1�$@�Ђ���'�����7�I���!�3%{A�����eb1jÕ%ɦ��}�@#���&�	c�@��7�^=�cҥEmH��VJ/>�Q�ɠ�5��c܅w�͟|<�U��8��5�V����i,�K���৏8��U5�؅\M/\�ʢ��Q�P� Л�)T��)�����W��<��Ӷ��@������~�t��
����l�V�	�}�(��1������>�� �NqQ=0TLϻ�G����UR`8�r�
N�8>堖���Wo\ı�-C��ӎ���r{y$iB�;2M;w�'d�eR��o�s��wv�;C!�M��I^ˠ8�J���Kc���<�$���=l�$,!S�?%gR�E}Z�(�@���q�
�B�2RJ�Ţږ�y��� �/�hOQ�@�=���,s��(�zڕ�:2�V�,��i���D�%�x���wYi�y.�]0d{f.	y��I���|�Q�]|̕jH](˄���̲rL���h�if��P���9�&��R2�)cYM��T�L�+k����bd(#d����L,ѫV����zLO���P=��yR��@�ۧ��D��'�]�����| �65��I��+ ��Zl����5��f:o4y���d���-���� �tK�6S@�]/���_V^��j��j�#�>ρ�D���V?+�D�>7_qN �>I��qd��rfb����/(�|)�7���O瀛�%�H���Ez��#{N�1��nA�ٵ���>��������d4���C��	�\Oջ(�����(�4XD%��} 6�-\�C�<K��/����
��3�����Q͌=b�@�P��&�*B���*-������dR0�Vu`j���?:PT�/Z���N$�)��-E�"۶����,�COJ��ƪ�v�*C�' ҷ�ڴ]W;�'�g��XY���.ڱ�5���;�X�xRt�4��U���a.��OhH+1��bb_X����M/x�[�刏lafТ؁���׭\�c�^y�C��B�AMe��?l�v��#�@=&_xpcͱ&n5��{f���V�ǐ8��e�'!P�杆�e�/"�9�jX�=n���C��C,Y�������o/0�����7��Շ��01<eb���Y��yEAy)����'G�b��S_���}��uvR������� lQ�������&'6�@q-?yQ5�v5 �a)�<'#7Rak�N~�DU��K_����ʍ��5e�c�ֆw�����#�3��2(����i=�0��yjƵp�i[�����V%�2��UП�w��%��Y�u��"p����U���o�_��m�< IQ�&��|{d%���g⎥ b�ʯ��Z�r���H4��{ڭ�j�nBp�|z�^8I����:"K���՘aKM��=�Jl��k�N���s��2�/~�k-;L��>4B��\��� �S�7$�e+A8q�i��o�8tVǞyh��YqXni�@/݁0ha���Ժ�fv2�ͻ�������R��l��U��u���:��;�����L�"�V�!hl��Æ�b�!Z@p� ��^V'�Π�>0�d���~Q��Z%�Jj��[�l��&f"�K���~�����P��;Wiӥ�,���e�s��~.�����Ot
G@&
8�E!II�}��9�SC-����r۾�	,�_�=0�t���
Fj�����2 ?Ra*GދԠZ���d�'5�P&��Y��U�%��Q��OVf�Y�f�
u�����cX���׸���zH:�k-�L9����e���.�Dx@�ҏ[�>T�� �5q}#a����J���)�}�b�`��dC�n�Z+	��f�E�~�����^���d�^Z�di�Rj\�մ����Ӆ�'�ĭu�J^Z�4���qߔ���ak�/je��p�'�/p����}��zh�Th��4�y���~�w�&d�_��>ق5��yEC��Pae��WN��bs���^.���V�ĭ���нF�:&�X=��n�vSq���6�]j�~Jj��ȚB�&�מ�|��}��xIؑ�q�m=�?w�xI�&R������YҶH
��UE��o�<��y�����$���i:���H�0Wp��[��Î�ҁLB���t�	�8����cɒ���?	[/���*�=]X[��mm�ꕎ�}���qo>(x0V��<;�"�%�3��^3�o[)�$"��+/�{�Kri��LuV�K���ߒu/�|������|�{<��1RT��<�F��@]��� [�E�j�ߦS��Njq�Z&�G��d�J{�TQ���ӛp?�,�'���E�J�(+WbY?����
�^iK1�4|�˜>jR�d� :Ld���F����L������m&��&VA��ۧU���/<�¶�h�nQ9}ţo�l>�3D�3V���N�j' ��������U�G��WM\<�sJ����ǙS��'���h5�Xr �1e6:��Q�N.
�Q�<X�U���r����A;����WL{^��5���
���u`dq�N�-S[l�{�_���b7yc�嶿-F�����؞�*C�4_%aX08���eL�8!/��~H'
;��P�����8e��T������=�`�)d�ht�*�^�L�CؐȎb�3��G7��8��l=� D���!��@i���O��������F�����u��{�鞯��ċi�<�6�QL�K�|��M>?����1����s�*�g5P�7;��Q�<��9Z��r�/�"`��A�͛28	�\�9 m���1����U�SB-��A�ySS��/����D��p>5 w]���`�u�	��5�6$�1��E�Q���,S���e�X#�nD.ئ�b��MS�G`�}���(�ì1>2Y�T��3���4��� ��;����:�-�8-����)��j !���(�����bh�%J�=(�!-pf��=Q�
лl}64��[�1�V_P4j�%�K�=M�m��
C�������4�s����.[�Oo�}ǈ�Ԁ�|<K�bsel��X��\#�:��>*G�������\SOh��أ�ǵ��q�+�#�|�<&n��>������$�A�)��n����wh���_h}��N�M��׶s$� o�(w�����ϴ�2�ǻ��T��D�U��2��
����.����õ���[��^a���b3�DE� �F���q�U�7���!�5�N�د�(�y���q��3q����Q�)��+��?R��j�[j4�18��aK����s(��#����z�Ut)r�á3��rSvD��d_&����<w`�����s��9"�}�KQ��.bB�vA�Y�m5���l�B��l�	��6Y^�Hl��z"kĳ��F����1+|uBER�C2�5�ǰ�X�8��ƍ�Z�w[��<[E1��� � z�,�$mN�����'��MR?3q}ƹǩ%`��Lߐ��zc�|�#)[L��W�o�����oA����N���J�5^z>/'�X���� m����j�i�'5�	��aW�a�6�C��k�ٛ�:vh�Ec���Lח�[X)�׺ӲĿ����Ӧ�jᖽ:Z	�2I��5�ia�R)*���!qD��lε�r�*��8&EX�P��g�_���ߥ@8��Mu&+EfI"�2�W����sжW�N������<lR]fJD ��p/c�-+٩�,[Qy��ǃ��B����;xa�ۜe�f���S��Z��6L��7К�Z}��G㐭7�{x�x�� Y��Szlkl
4��s�usU��xQ!��/	���:O$Bv�C	�i�oj��J���p`O}�I���~�7,b ����2~��F��;H�O!ѯ�OJ��@��Ao����L�=Xn��ek}F< (���g��C��PĳG�P��5�MӴ���u��c� �� �a�V��x��' �g.J-�㌬��V�-�`�:ц� �r�e�ӭ�P�b�TU���	���m�����m������f:x�� � �Mq�����޽C�G������r:(��I�mqƄq���*X�X��(C�~6nA�3H1|c�f5��F4� !3��q�fȎ��9��
[e^,��Kz��wH�0�a���4b���g�v�d�,���Җ��t���N$N9�ySm�sWs֣��En���a͸ ���FK��l;G�Ű7���o�ˉ�'P4N�ܩn<���������aGv�&l����!�>�7r�F?�	�����x���U�9�bZfC�yQ���y��?o��D�U���Ȕ�ď 7��$RF�?��=��"`�TAj�s�>g�2�t|�o-���6�� �k���Kj%��1��S��RD�bC�_D_�죕·���ڡ��[31`��_��.g(��*�d�rRwȧ(m�}��`S�7�C��u�$j�x����q&��U��(�ql&��Z�ەF��֫��^��˙��qŎ^F�86����ky�iM�<��/�{5��1y�t��I0�JB�7T3�/#I�RP�W�5:��S��V�H���f;������@�U��r`fFc"y)����VN(���};̯�Dji�W]��iH�-�E���!�%�}����t���2���dbQH0�<���]^�}O����^��VO��ݺ�%��S�dZ�hF��5�=� .��]�"ed�=�{)Xs�/=���sO
�Vo����:��f��3��*�]�eh�7k3gS�ΚX�o8����2k�T�����H �]#r��i�a(�t"4��k���ŚXƃ���~Y�8� � ����ձƊ��A�A�
{J�U~ԥ�a�k�&^��c�; mv�|�YbL����%��%� �6���Y�FQt��\��[��Tzg&���Wt��!�I^S��z��]�=!��^ܿ��<`Z���j��v}��5ʞ���U�	�����{;�� �T����	xK �T��w"��ˊS^(���I4�`��av�=Z��	�#�7�0������d.����kL�*���X��E�h�=��Z�*.��=�aQ����?����@''vɢ;j��gv�蚡�����cS�ޝ����,+�o�B�`a��h��V{���e��;��^w��m���?pӜ��]*g�JE_x�>���Jhp9�.��1u���@�h�'�9@!51tu=��q�$r ��]ye�en����=VLh)?Bx��[��5w_YJ0H-GJ�%db���@�`� ��?���)��w�c'�$����V�A�H�T�����7ϖ'v�{�+E�_��?>)��x��x�ROX>�?�ם.w� ~d����"o�;o�^��V:2t+�|��Ɨ��zk@�|ž�z���M������j��{�,����WUn�	 {*���&^!aig�l��C���&��|�/�<�n��r)�Gۓ8�����i��m�^Iqim$�N�<�m�Q��R�ʶ�`i+c_�0�@�W{�Ϭ�	��_M;����f��eN^�eߜ+z0&��DFNM�%��$����.7Lo������"���k3^-���H#f�����E�j�T�j9>Y������d��F(�eSP9���<,[N��v�v�{��k
U!�e��ջ]^w8 �l�7���-]e���i�n2�;%)�&?S$~��ȟ���4��t�z/&�C�IkL��Z4]��hd�4y��U���!N��t���O�<W������ߡ�)�= |)K5����([ϣOevq1�ɞ�����I����=5N�9ĉ���G����� l����v���ߑ׹�'d���9�3��)��cq�qܟha�YD4Ӆ����2دy�g��(��c��+s�G�X�U�(C�ꂣ�R�� ���|�3�Y���tt2��+�����Dn���m�ű�����A}}9��S�Ak�k�?<I��9���tه�<�t�>.A�չx^�-+� x�e9��K�@ܞ��N�q�OW��bI�cs�B����O�Z��Ͼx�Y��G=����ɺ
4f��x-�f����=�#4ōJU��� r�oM�rso����^{�9�D4�Ր�%ٲ^��~b<��3H�;�:}��"rFIEb��[�i�5��l)���(z;�R�δ��өS�=_��|30�7��T�{�2�an�?�]������6��N�|���.D:�{u��]L��)V�U�{�;���D�C9�^V{$�'S$�d(�@�4���)�,�Z�(�w�"�<�-Qm�h(b��2>��6ex2G ��D�J#T%43ŋ���P�8{ G�T>�Ca�>"W��|e,f�j!� ?_)�II��Պ��Z��pM>�?I�w�PQ�N�.DӞ@�%�e�˝��r����7@������P����_x��L홱���Ɲ&죍���|�	��M��r&r�m7*?��>"2C�s�s��͋0�雾)��W�b����	Z�#N՘�Q��Y]ŷi~h9?�X7��1G�$?�^����n;��f�������y�W.~ŋU�S���n��['Q���-�:Iˡ7�?�j���&`�vn�'�k(k�Z��6��g_7��'�S��Z�
�f`R�ͦ�!�`������F|�h��om0-?=�R�r��0�$�&��Dr.E�q����ȥ(,��SLa?d{g��.voq-ؚ�z�6��Bq)c��F����	)`(�v@�����/��N�����w(�8�jq���c��h��"ⳇ�DȊ�f��.E��҈�������]����7�Tq�:��^R�G�\Y|����uN��~�q���M$�V4:�n��"2H�<�A�谢�� L�Y���C@�Ƃ�K�i�Tp��*���3�ԟ^�]�"������~ ��sr���H�*ޘ�RN�6�,�3����]r����s'n?
y��@(�¿�? E����.P*u�H�d�w���Z���_Z>�U8��V�� �Е�y ��~yOL^��ž������䃙���>�z�;�������k��g};K#��垉�7@�{�g�X	<D;����<��h:3��h�d=��¼4�;w�v�Q�c�a��w��"�A��t8�.ʒ#Yh
�v�*J9� o��$��8��֜��b[���2�c��[d�nOK��8���cj�v��O�֡GS��������I2@�ߟ��i��i�!�c!��.Uc/��L�@b.��v$O�;����o�KLq+�e&D��4D<(�j�և��t�>�oϠ�X[ȱ��SsM�e�ʽ�-���镥��StXtqȿ_�=���S;S��oѢ��6�Z1$�n�UY���,BT~�J���{�S�v@��p�f�hֱa��=RԨJg�t���m�o����H�۽�٪���>�2kP�ئ�i�4.�{*���+V�To�L��TM]73�c;N�X�ь�yhH</�^s_[x[Չz��2��~�aō�J������lʣք�
�v�'��c�M�xK9WXP�g��=Z7�M�@��..��9�w6z�`NL�z{B�Krye���$�$����]��TT�XD�,���3�@tY�����(��r��h�VoƁ����Iߴ|�-*Z�B׾7��HwsB���������)�4�e�L��#�j��8�o���+���=���<r~�l*�_Q�]�ݒ�[f�m�����{���|=����ldPe]��F��6��y���Z�C|�g#C�QpǍ!Y�e4�e�,��=<��Ž���nh���4
�p����6�Qb{R�=Ph���J���r��܈�uh�����P���c"\��k��Rȱ<uU۳�)����;����6�H
�>7m:jq>`��4\��}�����W1(��*��׽ �ޟtB�i�wЇ���!��0O��1Ÿ���������8�l�ŴqGE�w�=� E��-w�M��"��d��:˦�]_{`ٛYrq�eaΛ,15�kf����N�.���;��c�f��`2�,���uڢ� ��v�*���9^cP�6f�i���Hc��x��;c��.��D`'<0yJo�KM��y��]���N�YU�o܌!n�z�nw�\n	<�e�|9�z�{F�=:�����%��NXA���Z��� 8φ�^Zl�B�>���/��H )�̒O��0���뢜%y���?c�P�o?�:5��̙B ��w<�0�
PSP��_:�ˆ��[Ƹ]TK?e4�3�F�Ak}y}]�
Zo\Qx�<�/�rŕD�ۈ�4�e���e1w�����hq�	'��˽�;�h�x�R�����h�)������7Z��&�%�m��ь,� ���Tb��:���_b	��>�� ɮ
p��5$����Z��z�O�q�Q�z����K�k��ڕ�5�O�a�#"6�ȉ��[���׬� �>H��X4-��x�o�م;��Cи� 43=o��
֛�dY��E��񜇐 ��1_�_�����Y_Fj���q�p4�N�w]�:�>�P��`�P�uԐ�՚���,��_��+ �5 ��;�G,�i�Y[$��a�I���4ngKj�A5��d��(bK�i�hv	���׀=�ڥ�y���e��/>H���̿}��hd�::n�a�茶���њ��Y&/'���py�z�@Q=���iP�؝��T~��f�n[��a%�B���%=����	�\��uc�����G�dA�Qΰ�[e��,����y^VVd�yD2M�
ã\%C<�M�����B��+��q����m�ͽ��Ϥ�v�6��J6%a:���!�,v�������a,��Y�����Y��a�9������lĠ(��� t��BP}(c^DLg{(�75�7U�����Ж���vw2���, 7���?\4�q��[��u�{�8w	,N��J��o��~9�{ipu4�=�(q@�2]\�����m��v�l�)̟�����#�L�������VY�bU�5��US���f�<�NɺH�ꊥ���D�����#�	�t�n<�BS�Q!㎤���k����/ruc����0�6	��YG��c&,I@�K�6VCo/K��M�`��x�΂��R��K������^/_1:�Oҙ5Ԩ�8�;^x1\G�a�/׀�S\]����z���)�IL�8�Mj!r�Z7d����6��t��M;)oP�EuAN0(�d	��J�v�|>�{{���f!M0�S�N�)-��P�%���6��7o��`C	�x�؊dn�,pvE��c\���� ��V�eT".,Ȅ���i��V����|�����2au�W_LQ�h��EJ��Vi1��?�tiM{lczӠu��A8�1�tЅq��8���z��@��V0vrX����"ы�N.�K���-�?��j&l($��רl���cNJi_'0�0i��w�{#T�l���Ż��r�~oͰ��-���O���k��&�i7N�}��Fݴ�m⥵Z�n��h�LW��?�Yk	�8�C��_P��Eы���Z)ֻ�h��f�E�Z���	L�)>=�w0�-H�=8�]���ut����ր`HY(sQ����iNMڳ�T�h����0��C�j?�/����*�tr�Uۆe�;#ХC���5nS?�+���.д%���N����x���F2F��Zi�kҨnb��h���&���15������]�ro�c�FA˒�-��V���uچ"�M)��?�fP*�m�z��B��8ڊ�;˩t;	���xpn��G	�A^�n?~��.}[v�p/7����7�S�Βڽ��nJh���q��
(OK��=�[���p�Q�/	�veS�v��6��U��*H*�q�������.�@� ��`�Z9��D]���oO`ccBZp?�ѻ~A�JF���y�z�����TϜؘ���9N�A�=A^�(�7�R3�'7-sdn�y���Ac�:ۿ
����/Z��o_�ۘ�dB��5M��ޞm��&Ĝ������ï��\�I��S��1��Ε����8='P�Ez�4!s��zc���b��X��)�'.�+�Ok���c#|b�U[����#�f�C����Ss �r�:�A��J%���r���}5)��D
��zx�ǒ-�~��]��mYuKQ�,'���o�b<9���Ә9i]a$����:蓏E�W~�&�)�< ���cz�]_�i�ˢ/R= L�o��[�|RZ�T1�@�h�	
2F�C������$�E�L���M��f����:�7�­�xJ���㚦�9�kɈ�nGRh;AK����A�5���A��K�C٫2�"ĵKUb^o�+�&��>�K�Z���/��YH�zDd�᯲���������]k��d/��K�0�,��?o�^'@'�o�^	~ʌb{X��ʄ�/Tqm}Q��3#�c�T-�� eX�R��$�H�l;�/���SmT�&h�~�4T��L�a������k΋'��s}Lx#;���*E��[M\u��Nw$��`��o吚����e�'����=sM���3�Z ��@ɵտb��m4A��wQ��%{���!zu�����x�9U��!���:��O�S�Ӛ���@H�4��m���z5H!xp�C +}�/�zڌk��˻���H| �Xz�d��!hV]�2��
eC�{�� ��b�F�$�5)J�����s��
�� �r��#��j�񑞰�0-�Uh���δ��U� i`iC~!�v����]�_��2Ww["�>#^�)�ih�|@RH.�0�'GC��El��2�l@̷D-.�4,�d�*�)i>��7ˎ=�@ÅG�.���qt��"x��c]����5OU(��W?�%	N�-њ׈q�FH�q���T��ߢ
�
Yo�ƍ�r�:���>���k�O>x�3:���]�<N�Kc�����/���mh�#�	@ॹ��׋Nߚ���I��4zC}�X
�:�?ngN���eNr,	��Y�H��1�a[;]�DTO�F$���w��{��{��ϼ���_�Y����&����f�@����M��QF8N��jǦB�F��;�T��A�χ�7$���ۋ��/x�h\ڋ	�F5FJ�4Qj�?��b=I����"�4��<)���n�74�oGZ�F���b��L�(|��3x��J�v�\��Bba��3�E��k�v��H���-��e�_�I��lIt_Ęp��x$��
F\a\�~�A6=�v%ed[���g��j�8��||M),E��ip�]}�}.�+�(����t���l�n�:����n�Z��ڞ��,�p�l��	�d6^�xA�����*"8D���gp�#�����`���o�:��)X��2(zO�+Chr�W6i{�2�3_uo�H��ɏGU�[�S1�[����L��<��c��+��gߧ �7�zJK2�o���$e�#��p!Oď���d�R&��M�X���᠆�
=
T����cZ�7�;���.3���H\C�p=�cy�A�~l���xô̨Wޜ��p]>/%}�G4�*q������ �kA����� EU�묞3Vܠ�Hғ�%��s�	&K������}��Y����f&��w�>���h,-)�0�r�Ρ�[�,ʹ���N���h����u���G���p/��4��~�ۊG�T{H�I!V�*|q}�@2��:����e�%�@��Ǹ(�%�[�+N��Y�+���Z>�PW���T}�ux�2�f��	�ϡ�S�WL��?�]�X"�Ǹ�*��)��<��<�5�π��PDв������'���!?ۆe���8	k�FDq�p<5�!aU��D��GQ��o��!V{�l|��8���$���Ǿ~�tk�	n������#�Hx�>zМ>���$�!lI='Ȋ��g8#����2	�#Q6o�+�B�_�D}B��;�{��T�_���QMN�\��FY�@�:�;�h2/ڑB�!m�u��[vlh*m�r��N�&;��b�����Ա�׹<M �������eO4'��{����v N�,A�|���=ƺ㸑(�r)��O���*W�>B8�N̨�������2(�Ǟ��kd#	�)%�I!k~.�*{U�D	�Z���ְX 4��4qP�,��Ś�Nmޞ���v��`E@�*�I��³�K>%�u�� 3��K_��tf�m��'�A���2M�&Y
�ĢL�Z�{��Bm��6��e���8��;����|[��� ���a�eD\���L�#��a�5��k+��35�9VJ�S3��89��1�rvP����oL^LBa���9o�j�}�㾛'�$ppZΓNv�Be	���N�=�2H*�����EY�C���(7��3@!haM�Ek�����jZ�y^�����q�s0̤ʈ�08Yj&Q��O���G�5�)fm��]�T3���)+�6�i=̗��oO��LH>�/�A��ʺ�'�4ϰ�1��=tj���A���Y;��p�s�y�ݍ��F15�o���/��#�࢜c�xn>���l�4w t	����P����A�>g��ڐ��hi0��;����{��ZV����ڂ�>,����� 3{5al���'ml�> �e@�L�ʳ����c�c%�n뒹��<��70}�x5n�s���H�<�hb��Brr��,�_3�@x%��x��o���%H�I4��C����47��U�n�/����i��M�������̩�shܯ���<�X��W�<������^�0����� ��a�k�,�V��|o�4�Lr�s���}�G��ƇqW�(�S�\&
�吀���/��~�v�T���a�t��9N^?r*2l9�i�=�:�O,\��\,�o
8���jU'�3�$���Mg�Tnb�/%�3�&R��'�9�����/�C���Mí�!��^��%\ Ұ���.\)��"j+|_qı��J�P3��N��8��Y�ҁ�f�e���t�ЩUiL�f��"��U"h3�w�vM�#�ͽ�C}/��������OET�_�a��}%v��f�q�t�M��cЕ F�Ȅ�K�?��6���ވ����ɿ����%�(^cK�Ov�=��ua�x�1l@Z���CDk�Q��0U}#�w�	��E���Y��p�7
�L�Q��Iw��h�NM�+����G�����]TM�ؑ1#�V�| js6�7?��U���!����V�x2�>|<<�C^=��������b��9�b���J�"	ש��}�xm�~rpI뻘
��)4-Y�������f�>�xQE�zx�b��v�P]��	Ӓ&�=�`��g��x��y�S��3�gXJ����>ʣe����STBE�����(0]hv��н���񴿰����孎`�8֌\����<>������z5D׺P��~�e�����qZ�淿ZD��P�Q�V�B�&8��Rob�Q��;<��͆�����%r ��.�������6
� ����@��N��x s�t�GHtċ�Q
�n9#�*� �k�l�$ai���M~����C-���b����P����В�r������1ғ5��ަ�[F�R��=g ����彔�ܣR��DO���y�+��=^�A�o��T��Z����#n�����[���JT
�!9n���s������wJ֞+��5�f���5P�C:���Phf�Y��;zճ9P�y8�9z�$1�z�q���&qKK"��� �]{B��1�+��1�t�?����Ƈ��P������p�>iJ���0س��u�Xɰ��>W-%V�.�B݋un����{Z~�̴^�k<�G�o#����w��T����$R�WmYs��R3�7b c��B��g�)XR&z^?�&q9!9){��ލ�̤"r�ы�BR��E�޾�O!&��sUq�V�U,�-A��i0�RB�H����z]g�Z�t)^ܦ����~̦�|�h��]@��<�l�S&2��U{R��0���e�R(��M,4W�3&Ifo�`�I��Vu�a��X��m�UjԷX0�����pX��:@F{}\6h�ZbBVX5������ϩpIa=SVs3$�ʃl4�8����V�5�,:0���6�+Ug
5��7)��g��gJJ]:}���qWv��Ю)b����ڊ�	%����S�<W�����=�������i�K�hHur�w�,���#pR�$^�`�.�k��&���;�)��~r!�d��c�ڦ
]3�8"��V���,8[ߠ���+z��Y�;^��L�ث_OS�v����k�x(P�:�A��
�2�&7���rk�8j	8�RUˠ���<5�x���A2-��@m�|d�ߜ"t�s�N\�p�br:<�����+d�������ȥ`�ҧ���=�j�acz��tG������5`�i�x�H.6��_q-ig_�,*�PL��|�i�����#?���n��dH���I'�M�1A�B91"��X_)������#�ѬW�o�S!Q �kR�=L��X~@��{�{6����;�x�0��k2e�0|)<S0@|G����L�#Ivs�>�qz���>�,��������~�,Y��{��3��fP(�\����o��B�h.\�KԠ�X���~���@HB`����4¶[9M��'��L;����t����{����~v�`�uHc��a�"�3�����H~x����dƐ~}���}�Ԟ(���3�t' }aFG���dcAi�Ų���E����� ��ٱ����6��#����dzO�ְ)���*��u8o�JЎŎԔ�2��J*���;�������N����j.. �0��CB��R!���'i��+�U>r���K�
b�K��Wn��¬u]��`?u�~=<�yo���&)���\ 0�ژӿ0r�	�w���'�
Ĵ,�(3�Ҕ_H��)+O+�J�J�X��؀SHnw����8��	X�;צ��X�4�5a����~�{Cϓ-(�-�m�,nO��e�՝ �70pbLfa��(!��9	�铓����rb�E~nM&p��֢��/&��q�7��r2X�1��p���*ؽ���u��P{��ϓ�П���0C�����Q��!K�XȟGS�~Q?s��_�ǖRڴ烁�P"�'�n?�0�*�������2-:������ߓ d'̛�l�BM�%v��b�O�H���ZСг����I>��6Y�e!��[c��Ak�������=��[Q�-/����y%�C9���|[�QF�)�3�tL�&��4��8s��H ��3�KM6�̥\ �m���_m~�KҟЕ7'%��0����N�s`�i�P�Y�"��ۅ�ogi7e)��ET���6��;�H���b��)\^9b�TVf�\*���P�	����y@��X"��*6���I�A����(c[R6R�����q)LڬPJ�v�=�Y������Q�t�Ѥgɰ���m#�O����2
��z����Ypi��{GF�,Lpm��B�ny�<�G���9���9W�z�����Θ��}pe�X:jyTW���a��Nٙ��������f����D���b͵v��Q���{�`Y���Ad�;2O|�N�7�����''u��K��7��	�Ҥ�hs�j�q�e@m=�/�C�9$��ٱjK����i7e���]��n乶��*_g0���,@�9�fۮǙ������X�͎F�R+������6	�Q$gz��� ��R$��|�Iy 5����ӠǦׂ�U���WS�t�����r������h�*1���B��Ʋ}���s����O�N:��/ ��rP�?��>����m`k�1�S���K�O}�wU.	J��H�8P�ZQf�vNí՜��d��v�U�b}����L�c��.��D<�P/没q�d*�����^����i��rO�qO�/��EI���9Ta��{�JM�RH���q��\xe(�jR,�F�,G\��?5U��%��U����b���?��{e�P#�&'$��8��Ly��1�<i���ZN����e��E/��ހ�[Pd�!��j���,-����ƽr J~����廇6��#���J���}1I���`�5����[���+�թ�kHmBYD!yB!2����+ui8���6ʹL<���yύR5K`a���Q���!��@�6����`�"b �#��#��O����(:�������Ե�m���b'5HA^�ӻm�����1i|hH;s�@q�.��39���XCy�L���d2ׂS��&����޹2C�[�ea��vUFgb��ߢ@8��:�!���V�!�Ό���|b���L23����YD�k0����y��������W(�����.����֕;'�n��sw{�����x2$[Sī������Y��J�G���2�ǎ�n,t
��ko{�T���=K��)׻{|�`�j�[7[sM:sA����w��3�[�ՏV�R>��#2L��+6p��YW�O�ap��$��
����~ZШ�@TƖ�Fy�&ِ���iJ'a?i�M�5k��B#�w��t~�v=�I9���8�:��
�׸���q�H���8k^��Pz���Oo�'dk	KeOȦu��D���Y	ET�E�@(�;��P�8J��p�1A�Ӕ0I3�Jis ,�k�	���3q�4�r:K�ʜ9�:�1T�bq��4�p�-��\8��8�O_��M�e+�$�5�W�>gd���k{�:k�.J�`Vp�22���b�K���;8��u���R�i3T���@�aiDi��>��QH t담��o�����q����3+���o!ݐvL�h|���+�?̑1�3����d���h��i����d쎼#b�"����[Sܹ�����8�"b�������u�5��ұ��,����!Ƅ<����m醳��e�������d�g��Ґz�R��P X�L�V�e_J9�5�ȳջ��Y<�-~�EL��*�א�|sϥ5NL�E��,�i�%�"'���|KG��X�5+Tćk̲-phu��'��/g;�o�48o�ޙ��~�� �)jМ�m��}���XU�ds1H�O`�Ψ8��l�Uº$���F�$//�
9W.&z��W���y�sO�
��?��[,���H���'
WF8Ơen�'�'�� ���U
�����+�lr���?�j���ޢ�F�v��;v�.���M��i'�}��"� ,��e��R��Lz����}����'x��b�]ģ�)�]�d�4 ���lC.ø�R�x~ jmY����=b�� ե��|�!�.�"ʙ���?�,s@�x�NE��Li�����nވ&�vG
�K{yK�n�XР_��o��ҹ��� C�����kg��q�Ew�`��T͔�����>�m0�m��(č�RWx�C�yG��`J("W�Qu�m*��M�Þ��^�:j�XM��J(����y���[C�Z��{��N,�8�� x#g�V4�� 6�M���DH�
��T�L�t��f�A�/�)8�E���o�� �7%2����m���x�x]�8MZf�V,e+B�w�����}��� %�R�<�����i�]E�0�c�φ�c�[���`I/N�%� .V��^)-�ʸkw��H����9����r�%�\]YH��"�s������\�ӗ�+s����� }B������p@�<{��'�!$e͙����;�NY�]���4���W�CV����%P�B��\oB�~�1���	2�y��0(��k|��Q��t�Ah�D�jY���.�ҟMn�������G5�j��d�y�`�����8���['��7|���8�ۓ��bӚ���Tp�hy}m����l��~��Ñ����N*o��Z5r"�ȼIYb#-,Omb���+��O����YO\�b �z9w!;	.�RL���!-F��,^\�j�Ͳ��ͥ�.���0�;��Rpr\(��!X[�V\� k�v����*��	i���煁0��2v��=��H{���J�A2Q��ు�S��_�r�<�Zj�~�C!���U����s�tP!�g�[n����a�]�6�
U�C@�2�;��'+����V� �׊���"�7V=V�Z;D��Hv��Y;�;����D���f9/��y/��Qlb��%�1����M�:jV3�&��9�&'��	���j�tT�=���n���L��M��p����Z'Vf��/���?���?��a��A�]_>0&��٨_ }���*�פ�_�Du��X
ޞ�� ���[���R<&�6��/9����@�� :���鑫�!��c)2a��6鳛x���م�{�EN�� P���>�]��#���x^�#9����+9ZPk���q��>_�������;�xı�Ƚ�����2�Fb{=��مW�����Gl[�&#�v��<0qZi��svc���#5~���X�y�3p�Y������#��X�M��2���l՗����lz7Ì)�E޾�FUHKp��=8�6�_����OxM�}�<�eљ��v^�˨��-�����t68�Fm63�ఛ�灓Ǘ��։��������x\��)���N��6�~<&����/cL��(`@��A����6��Tz-�}�^�8#ð:��f�i�:�h�[oj�r���Z��U-�kst�,�W�4���үc/�	f_5�.�gNʿ�9�
ױ��
���10N�w��ey7Ԏ�S�q�X�F�d������ټE6�U�?K�����C80����!"ZB�ԕgl/~9�a�;x���X���M5%��m�4̱t��<]������*���0�C�= �6�����g��o��p3"������\����V����Z�]�n_�֊�P�#&`s8	iqk��p����2t��׬$���N�bO�?K��(�SЎ,^��j��?��G<Hv��(?�#��z����հ��N@�Q���V/*�j���=;�v*ŬR���Xy�y/���G$xO�eœ4g��tR��D`1'M�o�����q:;j�V{;2�*�_I�����I�,�}h��J����z���4��=��zo�w�[�~Y�j��#�.W��B���5^
�Q�E�E�b���K���?T.yn��+m-��-+8%�S��bٕ�0|��7��jl�=h��W<��~��#LPs�_�3���_�	_��ͷK��~qĵ���% ����e�<�)�ꡌa k������Y�ն�]�s^�A��%����#���"�.���(2/�t
ْ6�o��1���Ҝ����~ͳ�}<:�J�F�ԐCٴ�[�^->fl��EB&��a�p��Ο	�E�<���3>>*��K�DUs� k7�o5����Z���,e�,IN�����̱���=|�����H-��ʓ�ʾ �Q��� 6	L��k�c	�A,k	�$�'��Z$�.䦺D�8u��$���C�ľ��y�D�� ����3�l!�?�n�Zh	~�f0+���0�j.8�='Id��ɱ�Qŵ��.���왕������zzb���Y���F��v6�" .�&��,oC��h�߄+э��˼�5'0���<v`�I�sC��%�"�#~��d�P?`��֎'��w|���i� hj�)�>��������\7#�o.0���cu$�é��q=f��j�+�t��� �p�.�?&�j�zx��.m[ �ߴ�ͦ;���5]��2ʬ�B˧�s>�,a�Q�}"��:"�P,|���4z:��.�f�x2?��.��ݱh�+��}�ĥq��d���XM��� U]�CWT^@Z�su	<Y쓬�lԀ���u!ը��H�[��s�`5,$\���-�R؂��s��3ϒĺH�e�����&�[\UY;���epz~�^���&6�*��{��|7:![�w��萵=t��w�	�q�Y�qeϘ�C%���fgo7��if�6�	��ۇ��l"����?S�[OB�Gk" T�c���� b��'�6�Gh��d�sT��%���S��<}(-�8�s�%* �H?��w8�N �Tr29q�_<{��5�b�Zy��E �q(�����n��Ѝ��Bft@dr�w͑�������)���$��� �W%�	�����'ם�;ZP{`�w�fκ�	�u͙Yn�Ӭ;��	��XC��/[���}��hgz�BkNm��Q��J~��'������Xq�PHɲ�30K(� �r�|8����W�&p�F��W�N���<c��q��7o6j�Y�$���w�Ƭ�n� Jy�\���|��40�i�R@R��[�,�jH@!�?����	��l#���9�D�Ĺ�mX�h�b��	��ߜ^l�r*��"�*a��V�"���Y݅�]���j_�ke�z�L�1į��5���*�N�&4r��b|6p�7l��3��L��Q��8n�M�B'RЀ7�c�JP#��VbJ�0{��?vԳ���!
8zv�-%��������Y\D�Lf�W�rӄ��7������tzr\��dB�f�诔C�s�x�j�C�a(�g�JŵYiÞ��7�T��C,���la��]q%nr�_�3�Ǆ,ܬ�c�v��2��V}�}�����`^awل����~b�V+G]Wm�Ä��*��<�|0JQ�%�r<�<��!鄪hN�)���'�q�v,�|U~#�{�G$5@e�M�cHn����]Y�zί �/!7@z�u:dt�����Z����O�G`3e��+�T��,{�^��h������
; �p�{+n���M��=�+����u�$IN�`qUM�Z:���S�RGJ�ۇf!�#C[��(�}��9-v�"P���F	��)���y(ֆ :Bg�J����>r�'%�(�Qݭ���[�5�?v�;g����,d�(��߹�F]ீ7�X�z��9E2Yʲ�M*8
<��ڳz��
5HMxK+�㬫l�dtN��xv�@��Η6Y�^���*۴"A��0���s �8�n8rB�
!�lR��~pS�(�|��K�E�R�ў�x F��i�q3%�1jZ��>���:��9v���s���S�j��j�J��	A�κiW���#�Z�WO��sx ��Щ�i�yыfݞ�'�Y�צ�o6GK��Z�e~�b� uܺ��]�F5�ei36�#Ae�^��%>��9��C�w5�N�{Q�Y��[q�=�Jh�K��Iu�i��S��n�n@z�p_OSE�f�S5��|翶oJ��$��p
��!�P:��3�TcMkN��@Aᅞ������(��K�wG��*���lE�����̯�s�&Ok�1�W?)B��p��A�&}�؋��=��;"�&Lr7u�5� >�v�źҘ���7��EA/%vl���N�Ԅ�%�Ƹ��k�	̻��9�of:���Js�/��$tE�x
㬏1N�Ǹ ��������]�D�tԢ�,�k\��8�?��P�����Wg۱�˵��i>G��(}��`�=��03[��n����9�����u�(�t1-P��+(R�Y���e	 ����Z������D+�?�q�[�9���7D���#��GLd���WZ�_�@6�d���9T���;�8H'�V���&�MU����!���@��W��.S�}y�7�$�r[�D�E��Ai�d��O�T�c�#l�-% �U�V��ɉ��J�c��';
�J�a����wD�s����3���8ewb��T���
��H����'MS�7+�qXv�^zO���~ԧ�����K��+Z^���H��Z�fB4�i��,�\�����\��Zۉ��}'���*��X�Ja_i�$S���FF���-���h�"�|V,�r�调�~���e�ߩ���FW�D���rX����g��6���6�q5�����ȍ���X���.S�@��ĥd0�"g�&��f��&�����:k�Q���</)ɼ��	��1"���V���;�Y�D�R%-f̣�w�Җ.ОKXu`��K�i������5�w�Z/$��7�����cA��f¨�֗�p�s=��r3�����duu/q��`�� '���'��N�=U:���0�\@��i���Pͮ�sAW��������8oMb�f\�<ΓL!�y�O��r=]E�Wq��d\����F�_�(�]��66Z숐}S���o3���l��Qh�N���賕Q�y���=�S�q������s	�2ݝw$�V�q����
)��e�Cl2��} ��Ĥ��WuX}���TȘ�,UֺY@��ԟI��O���m�r����6_�0�j �L�P��I�5mQ��J2mg��\K�F'9���ߓ��_�yu�z��[���Z�&��Wy��a=�zemMm�:��s�~f/�{�A���1}=k$-�֥{coO�T�{��P���&5�q!\��醱�%uZ��'\���ϛ��~�,�O��~؇&A�U�Ӑ���N�*<�'2
�>�=���;��7\�8d�Y��hj�E+���Ù^0���|��z���8񥫻��v��ٴ:e-<{����(�"��� �%�{[��E��,����2�6���S�m��M=g:^Y-�?��`��N\�V���qݵ��?�����z��8t�[y�b��@9������<�nɏ��Ϻu(=e����?���VK j�Dj�6���9�I��GI��/ ��� ��òn\�=�1��a���"K��1�s,�j�\�>8R�W�u�0c8i?�2{����|����W&������N�P�o�.�L�7�c�kZ�)��q��CoD�!�2E�s ;�>5��P#�¦Yr���{�q�au�O�2���=^�����	>p�	k�)i�q�Ul�sݯ�j.��n!�����]�+��r��!��Bu�wQO7�-Zn�e���������}�>G����d/P�G�
��C�������mUs��{U�";9�N䌿{��������jL3��Ȱ�G2X���pr�y&�������^+�<3;�$�����D��t�t�xӯMU+"Ǝ99���j�m�{o�/%��-E��>�����gWߋ̃hu��ϙ�#�v=�m"|<��Ɯ�DR�;�[��E1~}��&���{�N�+��A� 
	D�=�5Ic�k���5۹t@��!-�W�Z^0K��P~�^����C��I��l�i���Jz��*�p��µZ,j��W�2��G���vՀ�e?�5���B�U��T�hA��Z����daL�V�O���Ќ��W2�F��j0#�~�,�d{��>� ���n�� ��Ȳx3��@���Wb9^��0�T�	za��V�J4��-���/�԰3b�D^n���])�X�� ˮT��2�M���C�Yl��k���+y�^kw�/`�k�vU��`�����,�i��̹��ڞQ�iAX��}�s�
�_Jal��XQW�`+F��>������/Q|:
�\,��C�"��B�.��2"��G�������0�u�b%���`Bf�7�m����.\S�e�n	�o=����96�d�5+�zFl?���O���:L�ʁ}�Z�k���S����Q A�����q;S/\C��@�j�[2���¿SG�x�=g�����Y'���$�ҷ��6�{O��4�1��V?�N��I�5� ����/��?| \�r��4)�}� ����7"�mfP��(G�����+یI�v*��C0Yʘ.#ɽ"yg��#��r�;z"*����+*���v��~k��{v��R���eH������s��:\��d�LW{��l{Lur����nUړX�l�\�� 3OŒ;@$����>��3
��Wv/N»���۵���(u�e!��h�лޖ�d3���Q�H:�Ǻ��8\����`���c��
2��c��hl�̃7ZQ�!^�EH��(�K�T^ζ������_GЫv�6�^�p���n��TJ�a��׊[M)t0!ռ�m$�ݧ �<`�_��hq��1�	8��T��;�H���tv��Ȭ���&�#�pF(pf�4����pG��1�?7�n�or2F����1͎��$�%��X���~r ����ܫV$�/�.:�����b��6i/�h&��2Eފ@���9�����P	�;�Ņ�^@C�^tl/�`�N�/�)�ES?O5�=��[=��N��7�k�Dw�>!Ցӎtt���dp� ּ�ϙ=~DI���:��x�����G�
9@;��a���L��U���Te���V3[x�ӹHR|H �Ï-��J�3�Y�o�	R�\�&}k��K�+qD}�U���D'중ߊU^!�����6 �lP�Ɔ��V���[�n#���Z��J.ZA�^����G���^J�k�>��/ �i��P��da�!����b[�8a�&3풠ш~������*�\�H0ۅX:#���wy�GD �]�6v����T"�j�̑VN-q�?>���ɋ8�k�:�G�*i>Ѱ�`�_�1o���㴸���f�X��8g���ͭ���j��[F�����fW����J�����^T[�k�h���RM�����ׁ����j�C0��p@�
sw'�Yڿ��8��A�X�5��������&��P��J� R�Q�f��~�� � �M��C�>VJ" _؎��d0eq�)�rm�.sчwLt�(���m?�h�&�'���ֈ����ѣ��muu���2�{.b��dO]��;7�`(����7d?��u�g������]��;M��a���J3���dgٓ�ަ3"�[�\�/��E��cL�� �	���e�)c!�P�� MY���B�l�7�뀯���1��H�����'@j�Q�D;����/�Rl.���Y*&O�>�&m�}�Uius�eT8�ʗ����<J��U�e�u�NGh��/��O�t]@Q��@!q~Ǽ[\��I��T��[�R�4+F�F%��]0I�'��Bu!dP���i;!1��+*-yR��[8�`��"$o��CP�{����Y�����R�f���*yCݷ�ΦZ�f�C�����;��L����~|� :�,'F�қ���J��5�a\�i�D�2�
�X�
c�O~p�w�<3�mQ�)�r�i��B�V���bt4��`*a��DR�h[S,vs�M�]����n�'x���_$��:�E�P([���f��C ,O_L�'5KV�� �h�W���u�VG��x)y�m�L�|����12�4x�2:����#N����h����+W�4<�������1�X���0�F�������|�	�Z9�[����a�{�z_������a����e��y	K��&��}>+����v�Ο�[C٢em���g��H�'�z'����R�b���?�X�PY3/d�A<�P���TV^��?SϹ�0B\�:v[���0��艄�f�L:1�w��g͞ȳ�����%�a�������f�M��>�Ov�k�_D�}���jrRg���^X�Ŏ�;�s�$������Zvgq�|����ʿ���ߩ� �AdB�t�p���f8V�p:[Zc���X���  l�J��rD�K2p#oY��͛��ڟ�h�?q^���h�빸�l<i�+m���	��|zz�R5;/��=4�3�r\M��F�KG��RG
z�Bj�f��5{�y��|Xr���cCaҫ����Ȃ���
tp�AlL�%���{�`�^W��%����>�	�o>h��t��C�g��H<��/4�X2pO�������=>P�x���&���2�eB�R�<6(̆���Ǩ�T�r��S��D�b�xй��)z�[߀��'��xq�v�f�x���-��s��-Ya��i�;���!�?Z�N�Ѳ�Q:��o�F��D��`���y��8�{�Գ��l?!�9���i�<�����\\�����!�%�p)S$��C��n�m�[��d�|�M��q,íh]�ek�� CmI�d �NȊ�y�x^�y�J�#wG��굾-aat�L)B�:�CZ��"�Ue�=��#�2\�:�o�|����ګ-���zkY�$�s^�����:�h�aV�_�a�P��pÓ����C/��<�w�M~d+�p�<菓�i�f?Gpvb�ۜL��Ӹ��+�KH\ɸ[?-��Pr�@�I��f�Tc�.��8�9`x:������A,��S�ܾ�%¢^i���Su?#DI�o �
f�a�e���#���F�J2 �U�V4��>�Zz�Ϋ��oGl@�n;6� 77!�i��E�.�4{;�䁫���᱔
�y��ʨ�\	3,J7i��� Џ�f��b�v	�뉎�������A��P�s����k��Bhc������<z��9ݷ����3S���^�EB~g�'��25�G��7#�����N��]���h���V�^�:��{E�o�n��W��g��6�jCΒ��IA�⤣�0�R�S/�N~���9���%�/Z�6b5Z̊nv�̳���&�#�Ҥ�������"׺MAq���/��kM��z]�&U�+_�#��h�'����I�&��d2\��[M�o�EeX;	�Ȩ$k�r��)�U3մ�������|[�����=Ew���gNG�-��ES���o I��8={W�N��{w�SQQ@_]%l�ѽ��,�ە�A/bGR�lA������p���q���;�S�	V�0ͅcB�w���R/l�.����Ձ䡍�)����N����Љ&�@��i1�D$�Y���y�h��!
(��d��)��(DP�n�+?x)��HC���7�d0�5�#�SD���q?��c�Y*�va��.w�T�,~�^��+�ߝ�Tu��x��'5�E[�j�s�0x�����=Հ�|۹>Iт����]aEsz�U���j��ɐtg$*��I���V���Y��^-X�<����Ų�1�Pȕ2���2��:*r��S����`,d�`�$���At��|چ^eH1)�~q@.@8~9Aq��MI����<�	Dbc��=@k]��\H��Tf�IXuI��q8����ȅ�fR&�����I�pj�Q�_r���J9V� �<�J��0M�J�|��)[G���9
��u!�v�-肬�U�Ox��G?�X 2nǕ�T1$~�>�8f�s�B>��=3����6^��W�I���k�s�5���FlFU���Y�#�Q`Od�n�+>���y&�_���K8g`v��̤tl�&�D0�Ƭ�3A�K�w�H�o���P�-�O�H�b��S��/x���|��ֽC�v�R1�	 ��@�E���J�z�]$r	w�A�n��H�:��׹�� �/2n���RO�A�2X^�ȓ��� �ӋǷT�ͤ��q��NsZ��hUrh	��R&�_uh1��F��Hm�!����s��ś�2�9_��4g���u��B��A�Z�N�1�ܰ�A��.��F9�*�r�r(�Y~k��fj��l��>���z��D���
!��և&ˢ_[|� ���4u%�:Ń�ċI?�磫}� ����@�����<��,��K����^����w�؜��
��a��4 ��
u��+3݁�����=�LV���2�3��y�Jnrl��y��Ɉ2��8f*��%��w����@N�,OÈa�� ������J)8�<f�FL(�r��;��%��#{����}|s�3��\���r%� �N���n���'}2����_�3�ʚZ"��OZX��m����5��M��p��{�N�k5�m��[�� �@J���ʮ& ��&��,-~h;f�a�O�W0=��U�Y��GIf����dQ����0d�q�$��^���-Q��A�T�J�h��j��%_ah���q��S_��C@7Y�ߏ]L"y���J�zWd˔�b�?�p`ۉ^��%F�񘚽T�KŠ��釪J=��&�/���hź�R<��+>�
⢨&���*q2K��XU�44?ƴծ���ZC4
cq����L���f�*��� 5��k�t]��n�Y>�ԩ���88�x��|l�rX�tQ��w�`x�C/q��5��`fG9�c4��U[̝��r���4�e4vQ�e���0������.䢰vl_y�;W�����s�o���h:G���Ӥޒ;[���,�`<	�C���a˔&v�!�6=4���ԝT�J q# 2�jC�6�A$���W�$@�tAT�u�=�:n��ד~v�>K�r�֖lJ�x�.��ֺ��A���r��!��4vZxw�^�C�NS�	����'���i)�%� aO{|���?;|%��� kG)��
���;5|"Q����ʻQ85X*��.�{�=�c���қ�ᩈ���O����i��N��
��C}��h�����O;��xp��;��3�;��H��A��a���Eּ�c�\����*l��:}��G��@�:Y���CEp�O"���\��h�4�ϗ���J��̩T�!ЭZ��+ҥ	�vS��:,0y�*4.aѐU�:�
~�{U����Ba���ɰ�wO��d��+�i�x�A|8�bi��=�|�:{�'m�-��D@l9���/�͇��o�(rH���. ;�"#x�.VO�T��4Ԕ�i��J��R";��}/�"y�ʏ�z��`p'_�{2َbh[W�U	ԫB�[���\�U{��_��\M��Lں�8�s�O&��z�}���Mw��:�?X�Ǖ�7�8�U|	Tȕ沈���6���	�6�+����x���X�S�����,z��N�O���Q��^�x�
Y�Z1�j0��⺑".�+�r��M4�_"����i���m�9��=���z#|"Y߇��>	�9�7�S�:{�m�b���%��&��j����Wpq�e]�ǛY�	l�wC���i��0_���r�?�������ڼ��C�������mg׫y�=jZ��o�B�m�%{�!�����3i��F�?�Ժ�+�c��M+�O#y���>'&�<��)�H�n��&�9��_	������@VL�aw�����y��f ��r4;	��4�,Ё��`������U��R}r{33�Y:��Vf�F,]��GɱϪ^Hy�6���a�k؇�j�E_��_3�?u�G�M;-�c��o�R��SW�)[C��^lEH�9�Y?� ]Z �)e`%aoʔH�vʟ���e�A5��O�^SS�c�裭
.q�����υ\�e��s/$�~�vV���a&����CQ)*�͆���}��D��F�Ğ<P-�I��a��zQw�,;���E:@������z����Z�g3��r�7ĭ��#0n�I�語���u�s�b�%^�JM� c\zp>�X
Y�����6$��l�x���~֩�X��	$�2�#=�e:�<��E����5�-͘6D�V���j�C{�G��%D*c=h�ܽJ�
�'7ի�kb0�X���;Þ,���[d�,y����o(�`���:@��&�凒]��Ia��1�{�Lb�-ޞ�t)�ey�u�W�cRl�*m���38T~�J�q���B�RbHb7���,��\�_����tb������ڐ1i��P�J�#�y����X;Q�Nk�����hY��c��������	�E������c}a�3���|���(98�\%�:����g��\><Jk�����x
4�vN��J+ ��1d.i*k��8oQes��=ϗ�Ǌ�X��h�YI���6��45?-��g22�N?���G[�%�й��؄��W��y�^�G�����0oP��n�]�����H�-��hä�g���Y?�J�g�=2)�4��d��fTr�k�
����o��d��#!��I����:2�ܹyS����Os�xjc+����H��|��u�Gf�E�1���"���2�S���e��6ߗ���g��U.�O`ش�&+��@j26-����n|����ʳ!� �>�� #�+B'V�Ǆ�,qP�O(�- ǅ{<	�+fTqZʶ���7��kA*5�7�.��d�ݾ�H�żڜ�wpsHE,h��O*�k�"���<���s����nQrG���W4x��.D3�O_{��vLr��Ƽ��]q����KЄ���I�3�-�Jun) B�vd��N�eS~s���fۘ�Q�����gITR�)�r���@���"J0Hƞ�r��afV��C����ҏ ȷM{���T�3j�dD��({薁�#-��v�-��3��\%��P̍�R�d���&�\E{�&��;�	F�+�[��,�П�L�U��Z/� �+�%w{���@/��	K�)�[�ӑ�E/��Z�H!�s�;�)DT]������(�mI֌��}y̓��_6[ Y+.�"xj^�y����K���N9�E�3f�>Q�h���UG�p���h�m,��d� v�u�B]�V�����;9�=_�Է\�o�к�����.^��l��0�V��i�r�o̕�B|W�Wov���t\:����F0}AF��1{*��2j��I��ek̲�?)��K�Q��H1׺:�D��y�D��Q������v�|'�q�c"TC��d�
i��3�k�2&���2�'�+i8�r�,S@�$��%��)��]���<�g�r*�V��${��qB_�h��%��@�u�KO�ȃ�V�Hû�U��F��4hE�[[�g��m~k�;��&�\���pk_T�0�W��p"%Cf?x�3X�֎z�b�.���fȤv�ʸ]�ڔ�&Qf�2͌�Sw�9��5
���zXV�b��	CV��<��Vځƥ��e�v8~b����*F֓I� �'뼡��|�9$� ��]q�Υ��5� ܧ����K�!`=������O(>�j[���$
�6r@��ī!��+�^:���\_%B[��>�m�c{�'�}_��c��n����4z��������3_D������kh�Ԫt�$�D�֔��UU�EXG�����WQU�ű_�xj�>�{l���[��s�Q=W5���@��롭"���TǨ�y���7�5iq��7߮>M-��)n����<�FRդ�ƾ�w��^v��E�/A��fRhhѽ�(��rk2��V��^��5d��DZ���4�8�F�X��w���3p��@=#<R�3N�lY�s��y��W��9�t"��ñ{b�ױ�����8T��i���Z�D�nGj�C;����t}�;s�:�tM�ڞ��+��I��^���w�8Q�����B ��H��]9�{��3a�I-�u��V��4x�,n�3/?I�x����TN�0���d LCPG����u.�Wo�������_1�}��J�Z9c���C
���(硪���ý��h+[��_U�G�bk�1)jG�W�^{�D���pLs� �ߊ��О��HؼĹA��ķ�!��.�`��e�F��8a����D�<$��E�6F�X�(�r)R�<G�sɾ�GN�%oD���AF��۰�T�k���p!�k/�-� ۰0Jc|����1!�.Kr!��.�{�}�W~�fm�Ye9�=f���ι�ԙϕ}I���D���%�t�u(RSQ�a2g�.�d�"]y����RS��W�'z���ְ�ʂ�K�C�>�%+QSR����ܺOրS��¹�����!ږL	�m�6S���٧�~]tq�q���� �j�<-�wﭒ�B��_�[����1�fҐQ��L����N�j:{��qj�-w�ʸ�րz~,�����f(6�"�H�J�����XQ��?4�.R�RR+;�e*3j�����<�v7}l��>�H����J�le=ȯ��������b!�;�5�b�Ё�#�;�@NцhU(�Q�Ԧ�ε+`[��3�4��C9��Y,���^��-��.���ҋB/0�H���j[�W*jL��8�)��u�+�f��
Qy)�T��g�ѵQ��	\"�L+W�z���y���Kf-���*�]�v���感��B�CL#�H1���geaN�����2��Nf	���Hh���4��
L����*��;t���]
�'�����k�'iG���Dx��-f��0�2g�W��_3N^�bD�]�e�+���4�c1�?��20l?c�b���������P3��Z)H�i��TUw��L��aV��0�yJD��3��S�V�y�:�*y� >��4�Q���g�ߍ�Px�`l�<��%��&�'�}��[���&�@�èJq9Bf�Z+��_�?$��~H(�=+��E��ץי�L���	9�;��r�>����7�i�KG�.|���6ކa�mߢ��o[J>��ݹ�>����ڡ;)��T�t���B�0N�4��jR�v�4��(��Au>��)c�3$���<�S��T��уZ�R��3�#��&c��/�g��sa�3�˅����`��ʈ�x��0�\Y��/�d�!X���ua����<��[8��$$A��h׆�t���E���_'8�?�<�Ī������}��p:3:\�>��iҔg~�/m�U��<Ǧ%�@!�]ã�*��$`PN_� �_侩&�ol�>�\)v�t����6�Qmh]+��
.-hVUHB�,��4Ș2>.�������;��#w�_	L��)7��я��i>���g�Ao�t0!:�]��kS��3T�&���J�^�Ā}q��F��K��0�6��)e�����˼�+bbF�y�8�!��3Z���\��Fj�$>" pg��H�FS�/t"b�9A>F<�D�x����{�ɤP�lv2�B�_�z���c�%�	�l��ܭ|ۋӊ]���AF�f�#�ra!?�͈�)cY�	u��-w"XW��4���쉤q������o�T:�+8��JZ���|ꐏzKvM�����_�!�0y����eAZ��	�.V��Ftd7?�W����n]�vkF�Tj�rQ����.t[�~��g�?0��?��tx��$g��T�ՕC�)��`�Q����!��ʾYw�9(�r�\3�w䀜��GɅT �*�Ax�/��W�`����N@��վ}�<!����_A������ϝ�zA͗�󀬲��K.�6xԋ��?�׬��9�@�"#s���'"e��o2�M������/����oj����*a8�����Aus�8( ��y�����,�l^�~�6���ېE���F��k� �g��D�^a���-s�O~/�Ȼ��^�z;�:��j`���X_�D|���u�{�h����mu+�������$Ve���y�(Q����O:��_z"�����)Y�s�J5^�>R��?�e�m>-S�ݍ�)�%�Ӫ�R�V��N��n�[ދ=�.Xz����sG`�x���U���COӦ� Pm��,(s|�;Q�5�D�����t���m��K����Ϡ\ŌX�&��̳PŽPL�k��Ƈ5���=X�2�c �K8��D� 9C"�'��2jz����=����4�1����R���&�ĺ��qÊ�L�Pe�4G��i��s9:�~f��gi�Ԑj�V�hjp�����*Ѯ���b$���,�_ܫ��t�C��Uj�ScYM�U���-V͘��v!�� N�����cL��5�M�<��0���r	�_0YL(Ka�R�:��P'e��ѭ�(@##��D�ul��B��x|��kt\��ʋ���`��d��?c�>�D�"�؃(vD�;X�������K�����DkO-g��������=yP`ˢ�*x�b�udJd���pɞP�P�K_�]o�x! ��(ߡ��Fd� ���W��ߜrQ������5Pn����C�	����_6�Y����K�0���M����s7�}�NA���	�n0,-u98�n{�#���29����\�'a����il���t�	�x�4C�W�~'��a'~�7�Gi|�rN��f*4]G����dx�ِ��C
8���j�|$ҙB	Ma���R������'�)��4_2�I�Fu�ພ�F��ek�'yR�YB˜L9�-��B���9�p�2���V�K��l�&�f_BM�Q�q���c�7c��A���� �J�
G��:Wf�`�f�=O�z)Z��b�>(y2���1��]Y=_�-�hu�]��*��Qٔb5]��,I
X5D��G�_��D|,�5ƸP���:+�}�)�RW̾��1���{��G�	�^HA�aVމ�7�j�;J��#ao5×E�M�ci b�Ư�B�?������UD6� F��L��R+eua'��2/���O^� C�*
�.nF&�b喦���h�U߭A���M�Ý�Kc2���ȩȮ�.��'�ܕ����MEc'
�y���p�b�5v�;%��̻sb��Έխ2]��w#�}Cg�����C>����j�8`M-�f��u$�>4q�
!\�œחLȫ@.�9�Heꏙ��)_��O"D{�C�*r�? �cw~�'��6(�do
q2F�x�y�#x���� �k�4F��xr`1I�Aˀ5+@�����WQ9;k ����ĩ��1�u+pῊ�7:���^�!�:k^թ�NCH�!̸7^��v�^���T�6���=C�>���l���O�(���h��V �@�����q����ة��v�mc>�S��f0;8K��v\K��@t$�4��%���!9�W��d�s�llL����oqԔ�b3�6�ݍug��P�;@�Kv���7J�s�^�Ϝ/�آq�'��T4~k�"���e���	��4�����O0�m$A���P��e���^�go�+!R ���Ob���  �kp2V�D�^���|F���CR�Y+)]����^���d�b��(�+Y�0�� %}6��~#e��[ЧF�;ؤ75��&�&��^����8���� D���z9*x� s�̹h(T��ƚmUz���CB�R"�I�]�7 �|�ҰbE�߾�n��ɐ#�� �[x�:�$0��k��(���z��L���1�ȑ�P�Y-S�������p�}O�$a>��t���!7�2G/L,Ƭe�6���-5\�>�߀���R��d�N� ���_�m��5{�2�r�I��4� Ph=�W��K�3��m��P)�O��q��_�E���xP���0N���^��t�x�'�@�-�d{慂�K�Q�I���B��S�d��Tx�ԫ"/P�'��s����.��n	e�+�ˏ{y�.7�qRS���Aʳ�Ae6b)Φ"�hv� #�����<,����2�5�>z��^v}L�aFyX w'd��N�7�K�Tbi&����k;+'��3���A�d�.p,�1oֵES�a��O�']�'&��U�$��{~�0�����m��ҝ�8�r�n�T�p�)(%[�[ ��ǻL��0���]��
��㉃���]�̀��r��������\�B�[�h$]����d!$�E ]�x�g�;E��0y��k���]�6�Tۛ�	[�A�A���� Q2K]C6^��;��vOg�t�^�s ���gz��
W���yY�p%m7��ZZ�S������������?�����=&o؋n���~{�����Ύ��jyq��ʗxa��^_���+GQ+�>���殆��<�>a�� �:"}�)���ҍ�[S� S�7�+�������U�9��F$��G���/�| ��S���>M�*ݘ#�z�e�O�y��n�O������0{e��b�hO�!{@��Q?��=��$v�A��'�<d�����\���u��@���+!9���UC	�)�!�
�_ƔI���5_����V5[���#7Ok�ޏ����&����`�]H��c�ZWl��(�@��I!�Ԣt����H�FJ�'�ˢ�,A� �Hz��&/��L���!�\N@^�1niW�h�ӕ$v"�sD��޲�Q�tY0�/s}�2c4_*Yg�~e����� �zK�6��q4@}_6�{�l4�sDm� �;1��m�6���_���coY�9l7+?^Т�,�a��=�{�G��Ow搅��/A���w�J��-��P{ё��~1l ���&��J�Mȥ<��B`7;_���0�+�	��I�~�ܫ�N� ��8T呁��6OPqǈ!r�%��l+U����9�ҥ@!OGa��	�ׅs{�RSw;#Q���ٛiV{ەh��1 ,�}I�.1�@��@N�;�]��z�<эn`������B�@m��v5تF\_���A�q1��{�mM?�}�Pm+��@cO�sD�)�ӄ�U���,D�v!��k�M��*;�eMnW�K�=@���ϳ�"�x�L�r�ܷFHj#���_����숲ᇖ)*����"D�|sF���"?�\��]��eR�|��]�5�-�,qn)+Ԕz�.�A��@K-�h#*]��6j%���f�/��!�ؼ���z�
fJ��8ރ�G�'p3�]�)�t-�7,^֘�m��b)���������h�$�L�A|;W�c)�p]��9�7�&���MʗQ1�8Jz����ٳ�	��#X�$n��/j�xJ�Z���c�#7��$Ȭ����J�O�� �30�zSZ�m�d	|���}!����T)����K�	�k�i�sU=m���l�w�ǩo@;��2��ج
!Xm}�$�W]�4rQљ$�po��!L0��v02�����wg$7��a\i�}�A�~*��	�k�E�v{���P��p!k̥w�a,\=���&"����uCLڲ-�ALi���:��������͗:lLP_����#z�o��jyT�]li.|4L���`3He���lC|��|�}$%����c�53x_^�p'�Ѩ�P���.I��kz�P
Q8��B0	����J&M���N�Hd�(���£��L��h�Z�]�ñe_J:M;N? ��e�͐K�Ee�T�v
D�
i?�HF[.��6��ʮ���7X�n��U/��	b�:���K���C;��M)����T�s�6�O{}�c�= ����xv��pP�$�~T��f@.��������'�?�K��������|�Fti�K�E
��W��e]k��eݖ(`�ʣm���S+��|�tp��fG2x�!E1�W���
$ ��
���:�|�a�I�d�Gv�
	VH���o�̺R,rUI�j����rOȃ�<ө�5X�q�7� ��,JH����7�M���[�.��:�������t/�:l������o>=�K��Y�@�YS������Y�G�tE�7�z2nK\7t���2Q��ȇ>T�t��Ǩ�6Ϧb-�,�{EY#�2���T����$�2r�^G/�.n�+��ں{b�N�X�[�~��%3
o��qB&�.{b#pX��6]پ�?���۩I_*�i��Ȃ��6� ,wɞ�Bݽ��Q]���
���z�{��~�*Uc��@�,4ѱ��n*ngn�n	#F��O�]�B��������!L�O�K��{�JP�i�e�H���R|���o��8yN�ߖ�)|�e)򦅇��\V蠱�\q�(�7S}�-W.���r��r<� E2�ǫe8����hh��
:,%��Q����$;QV�q�9택�}�����D\l�"0y�~��rɉ*�rWM�P�&�|G(T���$�(X�6�v���1�H�ɘ�����9Zzw�j���a�+��iͭ�rO�����ӱ�5hh��Mg��C�묯�����i�08n�%;>.W�x,Gi�٤�J��W�g=f�v�n��u�X\�@]{Ӟ�:*���s������*���C�+�ݽ�h4�S�ʐӑ �@�."��}w����>�A ��J/�^��_mB�Bb�u�]�or�DT���*]�Br�<�>��Sf>�ϡ�o"��_r����YL��{�t�=��'�E�oL��vS��<V�5����d%d�f]�f{��o�f��Y;(�_��'-B�}���xR��4�?��6��z��8�)�"��6x��_��Z�I�&�������ѽ� �  ��a�|u���HSYܽP^�#��z����,��Q�t$4d�LD�T�V�o7��kdߒ���!��fM�@КY���,j s�O��Ɲܢ���z�m(�Bs7MW�Lw0ɶ�t�=�d�����ᏻӁ(Z������M�(��ϒ�+�����^uc@�A`�u�\��;��x�4�l�>V}�<cW'�j7�?��]��f��!�:F��U��	�.�cuY��T�գ@�_�G��е`Y�$ߌ�����T������u��]Fv�D9P)x�r�ڔwg�)��hmz�r��e�(�Q;�J��	�a}�w�P�!� 96
�PO�dV��C���_3����؈��&����H8����e ���L����qr9s5�)�:-�����uv9�+��Ч���L�y�l��0h�X��:��<��1�L���P���)���m�n���ȋ#:�����4$���P9|�oC��Kո��P�B�I�z^J	9@��(�E* ��|��иq(��������&8��6,\�ét��8���Ot^�gk��	~J���W��������ޡ-ڰ��y�S��l�)���-�l3͉a��������̬%l:�ӵԇ���ށ����yӧ�#�U��AU�i��9_l-��cA�v��ް�m�$�U��-[���� �la������:������"×jg�
`>*�����NU�C�f^(�[�k.���ѰF"G~ \�|*�};�퇇�6��Ǔ3�e��P��}/��"Q���]�!�8rW�?E�
D>�����4�!����ƻ��:��{@X	��,�α���ߌ���>9���c�8�I��0��v�g V�5D;��m��t3o��NÄd�]����R�"wuIED��J��}��	�?l��l�I�����ot(�[}���P[�ˏ��F5�][��4Fz�2B�Ln��"�"t���B�w D�Ʈ���� ���6��"�oz)����Q�!0�2��}�*L�ɧ�d;~�����5z.�ԋ�+�䶖U�Z���W6us^�6��x�FS�jwzW���(A�JԲE�[�4x�B��]!�)C[���. �;N����a���֪���$�]�_�N�Z���4�)���B������]ly�/�dWs���e\�cgQ�PVٱ���q����i�A��U(��h�280��������I����,t�m"=A���)F)Tj]��`���u���ٖ�I(��$�I��Z5���E*�3�0���w23�ap�r�༜��Tkρ,L�G����+nH�s9�4<ni�׶����|g�~Q��0z��J�ZU�K1!�ӑRQ��?i��^��e�6����Q���GEWR�5�dpN��s@DZ~_g^����Ÿ�ae���!W8MHF�(��LT�Ε8y�Yw�<S҄�'!W��4��('�����O���3C�/���c6%=���6�Ix��i�a9_5�N)b���u�Y�4}O�>>�����d4��ćY����51�*	��5|��=s3�3~9"謎�Ջ�܂�����Y�����y!�����RX�p�+�䪫�i&�����1�H�m<@�_��[���_T{�*�ދ�̡>��/�J3�&w�Lr���GJd��p�5�DMu$�7&����)��9ʑA+���!�%ʍ��k�a�s���u E��A���y���[W\�-u�Զ��^���Os����{(Pg�������F�͉]�ȋ��2�7žl����髳�؀�S2	�,L��}ZʵU�ƣۤy�����1{:��Ajr�nm�X$Q��3,���ٸm�_��70��d����x� ����j	�Ht�1����n�xDrXFpB0�9�v�PD׹]Kc�zM�	��o�����,V���--Z h4%��L4�o#�Ĳ���+�MdCD��D`Z��%
W&��)�3B��(�,p|�8���c��ZA��;��R�{0	�@���,��|S��[�|_h5����WE���ľ�e���**�����>pX��,��Z)�����sp�Z����"J߮`����:3$;�1M��?��%n��6�"��w�-��DQ���Q�.���c��U�����ڛR|��U��fj�De�&���P�U�`J�ں䆨xi	���Pk�J
��w�Y7���� �w��b�Q\��RQI�UEh����<[+������iMrK����	���aZ70Y�H�bt~Mm&�u���m��������k��3=1��x�f8�X�������?���A-��%ȣ���e�T'�_\Y��.�Y$-�C�+��7EC�/�M*X#�7ᆩ�t2
J���B�X��#&���J�������1ǅÇ�sg���N��|���SS��&͈�L�{��8K|T��Db�Z��#\����6g����D��y���uT��!��K°�~�܂I�N�	���Q�6�E����팭Ɔ��V�elѵ���Ԁky`��(�J�:Hsp�d}$�q��H>���j�8O��O��hA3%�W��>��E���G��m��E�Ώ��;�1��1}�#θ�y� ��a�'1`�@����J�8H%���k�X%?�HM�ץ]l����ߪ|�ְ��S]|ϖ��A�R�h.��$�V��cZ��W���U���j����CE�c�ڑ�E�Z�3p)���t),o��dQ@b�)�"D� �%�lB����u���8~�[��2j4�]H���1tkG ���JX�w핆ҽ�Z��j�����ϓ��a�>�H�yW�����<u�a �xa������=`�]�2-��7�:�S0W��N����B0�*e{��ș����\i[�;ufiQ�
�۔��%��.�غ�v|������'}�*�ы8e֌�~�z����-5ﰯBɴz�f	�@!f��9��}:@1�lf>�T�+�{� ���Y��Fs^�=������^Ć�2�G/�1;�q��>�=�W H�8�'gee;��D�C�� @�P.�.բbf�g�z!�*��:O�8���f���R������������<;�Y�;�0ž�A�R��(���#�����}��	QRo6��]#�h��S6��Of�! ��ę}�U�i0�����	*��Uz`;ur����<���c�K�k�kR��l�x�F���a!�@�3�{pe���,fV��oA0�v�GP��*G�[���ƺ���_�a�������g�1w��N�Z��$���pl(������<���*"	b�snP��D+�J�s�Z���/>M�.+%@���<X�r���֩#�+�یH���";�T�m��_��Ǫ3zMD�o�UjLD�n��P&X)�Μ���ػ�v�ֶH�BW�G�B��*���&�t%���|OY�<||NN�I�:�X@���OXo(>��n�~��1���;��,ְCGW^DX�b=H(��¯ U��lt�l���(�F��
d1t#՛�-'���l��ա�-齹RSZ.I�hx8�P �NI:���'��}"�I,_���]T)U�Ab8�҆C@�\�i�K��;�a:�:�@'�H,ʡ_"5�����aP���,�!Iڠ}]�O�h�^�ȸ<"vwSy�^���t���7��G\spg���YS"�"lFa�� (d�8sX�yŦ��e*)m80���)OdP�Q���և�,o{��_���(²��g�o�n"Z��*ci�&���[�V� ��ƍ��R�K�s/���2������l-�6�;�澴[+%�Tk��4�L��w��3|&!C���-8S���̾ڴ5�`��u���
�R(�wݔ�P:��'m�+>w*����@���A�m�I%�J��o������8`=��U�ۺ+��!�W���8�-�,,omZ'2Ԗ�)���f�7��{�D(�/'�)οf�?6������F� ��#
h^9�� ��X:��p�v":%�E��
�0h@K}lm2�N��x���^���U�s�����0S�?���YUy��b�8��Z4E�t���P9K���������}���!�s2TQ��	��t��`�(0t��S�C��X���qh��2��������,#G���Dz8�X���o�u:������g�-a�׻f���O-	B�2(c��@.��x�ΐ�y��n��x��u��3ў�L���u+�6��`Y�I~qtBT�ɗ(�]-w�%ojL��n����������G	EG���VK�La�W�a�Y��3�����{����Hū0���Xv�!�Ϟ� �iF<q���z��B��?8]�ɸ����׍��oa�,<�?
��X��3o�k�ݱh,Nv�~�]�5 O�Y�5;f��:�4����c�# a�q�{^�!M~�ש#)u�� )ݭl�(u��-�H�n��jc�Uf~y��G�����:ef�	+��Էh�*��`�д�j�g�ģ|��X@��5���(��c���?�w죊�)^Bڄ> ���"ƃ�TX�/��`�6�B�$�ﶣ�&��@�ӂ�!~��X"i���LohJy� SVL��
�f��~���͵V�Ą�I�W��E�ڽ��hw.��q�#���S�:�k/0u�LKz!�6�� J�v�7O��CΎn�H���#5�:��(���/.��B�k��Q�u�k�x�FQ���}9���
��ni��b��Z��Ц���)&�"\�m`j0N8��[i-�����碞�����ԃ�Я�d0�%V������f�v�+�R:��[]/��?���K�;���6h"����jqt���'2����73�4�O�����(A;����X ^��b@y�|�:�����o>5gR�I9�(۫H*�k��/dh�v{��5��x�EC�"�С�D�;_��+n.3�}6>ʁK�as�����U͍u��ӕ/ 9���%��G��%��ǀ�y����oB2�l=(�1B:~�jH�*�JmxR�<.#� ��;�h��?�v�^Iz��x��ϥ	�bY�K[
��d�<ݮk%��oBr$����FH�y�����GVbhx����	|��H�\�J{C�%4m�~�l�&�`}b;4vla�r(�U�k1��p�T��FJ��zE�B��9�/I�����/�W����P�P<���w>v�I@L@_� ]�j�/�����e�m7��O�\X��Lތ���f]l��\~�d�*��qԑ���_A��D�!�w�g2��B�]�@F��~�C���%�N��T5e�X~V�Ж�Dc8��4�؟֖�Kl��IZ��z��}�3H�t%˿���Q�I�P�_Y�	&��K6zH���
����΋9~E�'PN��wcr�ݩ�����q����~z�`��P*�B��_��X�M	�� `�Ć4�V��Z�S�%����le�bQK�!E��J�ū�̣��/���n^h�1��*��;%�2Z-�خ�����	��G���w�맖vp�E�_��s����mXb�}��RUHF�Z��J���T�����o��D��7�C��VI���_����v�`�Ϸ�o�#��7[��|�����GWG�^P��gy�" ��\�Nv�+��Ǡt��h��eM�\�;��	��o��G��	u�E��q|���K�X,\�7�T!�[w��x��-�+>ֵ$A.C13f!.����J���}��%�d�
绸+���}܂)z�@z�q�hU��:�����$��FNm�c.�����_`�vG2�����)o�t���l�B��oZ,�(H�K>���
+
D�_�(&�7��JJ��seCO��Q�ZNs��+�y����x���,���h�yp��U=��>�b�jN(��@�
Q�g��L��{C�����H��cb��^���(F�;I�������X��
-�fe�9���=T�مpc�'7���F�����n���`��~|7@y�����הK��\tw�Lu����5:����?��މ�NZ�-������C�B�Ru�4<dR�#�z�M:��x����:�<��=��J���u�6�4�c�A�o��e�[��z�\��j>	��I�Gy)LaG�s�ѩ{ X�IheU�#H�ϒ��2�G��l|�1�Ȣ|t�՛N �}O̙�V��D���=* f����C�ӛ�«�sB8k�z����g��,k �9O���8�UJ�v$����'�){�rn\
�Yջ��ɒ��U֟����Ac،Jۛ,�]/:-�lՆ�ch���\����<���o��V�~�#��S겭J�1�3H4�eu��"6��ҫ��>c����jT��f�5�Ǫ��`�2��36�Z�7�YD�bc�Ů>��7������X�s�br}]�<���ۏ�����a7	1�}S˖n��ԅ����n���1q�`�PH�m���f+oz�NT��-IA ��*b����af�J=�[����ؓ	�I�eZ��r�""���i��g�<�Rr|3���2�sCX >Q���5���d�t���ىeL��ڕ ���j8�m�:���T�4�K"Y��&!,��{��U��#�e��� �P�9��_��ز�Œ,F�BD��Q��H'��;�eV��k~���z2�5��X�� !���������i�Pz��Z�y�;�ч��]�%�XV{������*kp��:����b�s[�L�f���A7�!��B�?���^�C;һi0"�;z�?��6��b3����[�U^����[z��W����a�!~���Tt��G�o���H��A�a>*J�)m��*��5�VS[�=*	��c,��ǁ��I�N�����-?�����c m�j�:�Zxr3�~����5���"J��Re��� �4f�ǼWB�}�c��&���='W��R-���Հ?)��*b�C�φ_�l��
�T���J���y�K|��O`n6�u��7�9,9�R\��mLH 5�[64F�G����X;� =��ZRw[��I�Z�]Ns��'���e֬�9A�8I�mk�ر�7d8�L~�VHs���f|	�T=J����p^��W��o熇-o�ͰxeR�!��s���A�0]��]��06:!;��FE� 7��]�e$�H��U�\\H�^XŪ �i�ln�U��Ȉ(��M�NQ�C&nK�J*��� "[�gV��-���%��h+kU�'��C��(�R�ڷTyI���J�B�L[�Vw@�7��O�&D��G.	��7��~y~�/��x��W�W�\�_��W�a��VMŜrr���^�3<^8/#�K���k��U�͛�R���ʁ�&|��#��@;����*k�\J���Nh�B�a���1Ɋ	�RzX��2P�$b��7E���������p�+�����(����:O6{�g��o��B �Nd��]�|�S������29V_���#�XѬ�	�D�����'*�n��
�J��H-MK�_�\�1C%��4;�e=/A�"���) �3"���D *��h��A)T\�xsuiZ�#,����oR�J.�{�+ǘx�]q(�)�bM0��g�V5-��08�Ωpɮ�&���Q�Ao���}FL��O�vM
�
�sL=d�d�Kx捶�z���:�g1wԩ�v9R��9��ԟZb�#����3�PVez��E3�]p�V�7����{�`���a�QL����lc�����P�Ȫ�׬�u+�A/���/S0K�Qߡ���h�k�âG�SؔB"_�x?c|�կ�x- 6���#����mph6B~'�}[l��Xˁ�Z�#4��O��n�j��.�┅�zX�d
򎹧�H��4T|�s����vͭ�e$��x���@"�H/]��U%��"�gs7�D��W�����u�.M��qj��V޵�P7	�x�M�bhl�=�PO��Ż��}��QnFi��_YI�DKS��~Q�T�~q�>�������_��P+�4�Sp�4�Ԏ��`VP����k臬_^��H�����η�[B��{'���hq8Y�3���q;�Mz�	uV��O�f])/!�d������9�(ǣQ	h�'	�++2p��nظ�[��:1��B�lPCS�ޗ�E6�#,褄�EX���ص�@Ez|�Q�H��j4���[qC1c� *f��a�:��=:�H�G�^�������b	�( 	ɦs��?�6{΍P��S�6R��C���Q�hS��� �(+chn�x��	�nm����Yں�Hgo�N
�:Mk:\Arey�݇B�e?0�*2�PyIH����|K�l��S�X�[)�xhe�0���^��<3o	Q�7yez����s}��Ax�*b �dA�q����j�Bž\0��a�36:�0�!���~�ճ�6�U� T0fD1���Q�X��y�!�@�XR��#�v�B�-3�i�;�q�ZS�����?��5+���M]v	vTk�Ƚ1r�=bLȼ�a�2H`�<�����>�����>����Z�n�z��wx@�֔��e�8Jv��bFB^��'%�]��C�/+�@���;S8+��pׂ]���0 �&r#Dޠ6My�b9�~Ђ>�{x1J�]W��ц�|��my�w���b�7�4�� �M��l��0�M��4�W.e$��P*>��y��ˈ4�0«���}Q�}^x�l3�_I��S�^�����p���&�ʃ�9����a�ĒI7�B��rۡ����]$�0���n�x���I=��Ed��(�Ȑ��xN�N�����t�ה�&�m��gi����n��9���)��9sw��B��y*C�x�7��.�7�����Bt�xV��[�M�z6Jt�=P��m�φ���c��2�(����t���l;����+�J��u���{3o�$DO�n�q�w�b��!!|�b�텻����7�d�?���i�ʕ����\�OD/��\�v9-���&�H���d!=��a���>Ǔ(�T�n���WK�0X�(R��'%�z��ĩUc҂�=����p��U���������fBY/߅�i�\C��Ƙ#p}9�!�}${%m�&�ֽ���W^�dHn����*�͕�y��P0o���P	����/�\�߫�9D��Te�UQG�d��^Z�5���ώ9�R��:d�l?�F�p2�[e��K�� ���?O"��uo��2�)�5N�u�ı��v��>��j�,'�|���F�߷ƼI��3U0}4�AI�����mJp�VW}s>�fǲ3�:@�X14\ϰ!�)u�Zq��^��Ij���t��vFp��8%Vy��aپ� B�elV�l��	�6X�bXJ�2#I)�e!�T
�j{��?�n�m!�jq��p����>�p2���_]��@�_t��G؇4��v��!3=h�^GWO�{�S�[��O���4�}����9x\+�?S%ш>��!G)���}X��Ȏacm^����+ԡ�i����D_��"��t��Py�����,���'�����a&�^�� I����U�Yɔ�_s~�l��e��8@��B��M5Q��{0Ǩ�:%ݒ��@f�?ϒc	��ưR������O����� Ӎ�+��=x�!W��o�(3���"�uP�4�%�x�Ӛ�v�����ɪQ8��;`[���)����_��f��h�{h������`j���n6?�.�;�O&��$��' )��b�u 8� ���è`@+B�w�U�tq�.�]�(@�D骝�>�(ʞ8��,�ȇ�#��$@��"q�d�55/��v����"o���H��,�����% 8Q�K��5���_�����o܆0�l�ޖ���(3�����F�������Ks�����Wu֗�YW��e,�NN�0�%����0�y=9�Ƚ�S�nRb]{��)��P�j@h��9M��$Dz-�J��*��6'm?]��	q�лu.�jx�B�������R�·�CFEp��;�C\��v+D' � �9M����pr��h�!S��d�x�sq����Q�;rF4L�x^U�Q<W�%c�3Vr��!�TӀ$��[߯��ݦ�98P�i:�]��:�E��9���v˵i#�93Π�r���$v�;`",F��
��#�#����C��,]dYP��4\C�$
��!�qO��Lz��?���#S@�9)>.��c�h��C�|���CA��a\?��e�6j�'�V��:��>z��"�K�8���I�}]@��Z-\j�A���Pz7�>�p⨚���,�c�k6���������V@l��z�u�hϮW�2�L�!�2��� p��m5@3U�i�í\h�"��|&]sl�t���Fp���&��*=�
��[��-7�MZ��2	)aϸ�^�w��PA3(���b��b(��F-P.�@�O=:�p��9I��Lys췃]���*L���A�O��9iJ��A����*ޙ��զh�_�j�H�l%5�+�(��Nf�k\�y!T.�˿��$�	M�׬c�2e�i��56��p^#s�>�J���C�]h�?�<�,��y>���v��� �>���f��5r3&v���@<X��Cм����N�Qq�r���5��#�׎c}�]ő<?�c�D��2�|��/:8��w�.�͌3���Y��\:A��\�e�)b< �^�v��C���>x�( 1�.�W���g'g8\���
4��c��n����w��k������Q�&�k���21�W@u�;8}N�e�Y�Y��c����T������Qvс�gH�E�����i!�ꉌ������Ԋ������A����������i_�ã����������^7A���ȅ��"k���u�. ��	ߴ�����ךn���=�6E���-�.����L�3�{F퐬�FJ>�q̌y�K/B����!_�9=�>�J�Ƞ���Tf?��sɂ	��<�m�����^K�m��-m0�=r\�C��?�9�6��n#��h��	�U��N���Q]7���ذA���^�μ��1��bR�JC}鯅�=y����jfT�x��ER�6,��л���p�������F�X�M�ҦWsr}]��y�C.��7�b��c�l=�>��:�~r����Sq��Æ?hk!,�1��Lx��nX/w�V<�~����LY��C�l�{�GA�F& �A�J��>ĺ�`���,A7����v�����}��MR� pA��J���-��Aa���\v�a�͚ K��M	��.�@��lMR�6�Ґa�$�o��#�X,R	�31�!̖�zа�Z�$�`3mA���L0�o!Ml_ZeZOn�._�*��:���ʒ����〴)J7�Օ�uI�b#�?�)�����2̋���EM���Ay0�GS�`=��|���=>�+�<�����ˍ��t�L�s�Lv&^KN����K�f�3��vἻ
����W�.[���`����Q��Qf7��h��+�4��z���\���MH�9}<º�����Bu��w��"#�,W�$[#��RۨG;@ �s���y��G*M�|z7���|V���ՁU[���y9M���]�n^�ps�{�w��N虥׺��Y�;j������^�-��W2*>0���+�m8.�:��}�E޶=�+r�pjP�V9o�}��aV���vw�@�N�S<B_��MH�V�9Q	+�w�uC����&j6��5d��R�v *� KcL=��A�o[��G9�b ɧ��t�hz�P�����i{B��O�\�.����f�6�)�`f[�k�^��Hi���.��/�5�u���|��"��J�|-D�m�,ԞǼ��ǎ�oC�<�3T��B�dL��g@�8+\wď��s�j妥(֬bQ�P���Ο�J��	*�C�?��3^҆-��8� ���g�����?��w����82�X���H����J�Ѥ��vYB���Dt/�1M|WA�q�+[qh���?�-�>��A²� dK����@�Nz��{� �%� ���a�xR�)�q%�.�!k�ʳ����:��#�6>	R��%+BW�<�̎Ue��+�DN�z��:be�������#�)����GŤı뼙S���u�_?p ަ͂r��"�6OѲ8��Nx����:3�C+�������)����R�~ù�]?څ|X������y+�a�E�4F��l��i��?|����]���e���B)�ayκ�6.��\uF<0D���qo�?)�r?�Ng�J=) �X��UT��8A;�"~���a>ڢ�ĲjH}����Ο��ͻ���\��"���{ͻd�c�����64/T`ӹ��*C�����y�}WKH�:��dBf�N��[)��$#[��� ��/a^j�a�"r��	��:^�=:��l�Dŧv=���U�p<zGe���3Ib'^�OIf^Z����0����Z=����a@x�]ʪ�D��-�(�{�1"Gu%ި�6=��$�/[�ߋ�H�6�Έ���$�l���'k�ق�v����C��lp:�_��V�U��%I����?{Ыu�g`���Xz��k�JR"|B���8��1�/b"� ��1@�����Y��\��)&hˬ�96����N	^�8i��=��~�t�uN�_-��nMd�G�с2������.��nD�b�b)1a`hj0!´2�^Cj3����A��gwp+�k���|(���1��J��	�<L$@i�C~@������߿�E�$l��'~�"�,l|�¦�FI�
KYR��{6�^I����B��7�A}�V �y����?�|Ă&}����w0��J�_� ����Y2알7��)>#���p����D���)y��^bW�{��fϘdO�1��>���ݑ���z�����C�e��F���@!8�����rc��A��y��e&�Ȧ����g��W��- ,�9��u��O&"��-{3���b���!C��L���V-.7 ~���b������	�]��w��:U>��7:���JX��ݏ'�N����Z]�y-�x=������پR�L��Rˇ�.q�"ŧ�%i>
<��~��q�`d�A�>�p�t���ߔ��Tw*�-�&5�,�������#fӘ~���L�,�r������7@=^��%�w.����z��i闸���a�t2��?6V���L9��.~���8� �o6��j�F���i���ɶ��S��9u%�+��3Q0�ܧn'�>Ֆ�z��2�k������%yʱ����\�)�!ޖ�~����o�҈U~�o�̥����!T}E25��w~����{�
\�/�Y�qs��7@����4�<І�K&�M��ݪ=&�o��W�A�Y:*��X�bИ���CX8j%��@��v��T��e^�KNn:����FHsؠ�gyxܘ$Z�����7Ǫ�_ٞ9��1��^��gurK>�p$~���3�y�Z�o�������Yj1�nY
�\?f�$I
���S��K����l��J!�d�3��>Rb.�]����B�b�J5p���zD���um0�)t��G(�C���C,�bu����(k1ۻ�gab=��򒶏������_���xo�DM�� VZ���"Obl��4�g����M�r�g�c�R�u�F�2�Tc|{b2�ԙg΂oٟ9Kg���r�[�ư�Ǚ{��(�Dg�K�<�8R��8�2|�F+�T4�'� �atٓ9�F�-~F ��a,)^4�������L��U��L)#��x��@���3 ^ר�H��6�8���v�S�6�������E|�!�py��3��o1s�~�E�U�6�f��?P'��]�^k�rh"��n_z��>�g�''Ľ���^���,�����B?���Ɵ5|4B�@ۑHC����*����`�� �@fˋzC�m4>wIʻX���d�bP'�(bgU�X�ώ[����amE��I����_����N�Rʢ5�����2/���y�Z%N��s�q��Xx����j�}��� x���?L��򑪝�á(.�¹9� ��zG��
�\1Ǯ�g���s�)�dc{!^ٹ������a�`��=�������I` N�0!$��u�݄@�[S�"ւ�K(��G������G��Gw��~�L�����{�ܻ�j���ވ�?���o���I��_&T�N;C!��
5�(O�A���nN�aocW����F�2�����N��K�h�nu�b�u��gT�r G�[�ĕ�2O��N���K�t��mv�-����0��\W���-��+�`��g#:��$��/�k��Z�8�].%r��ո�t�T�u�@J�>�� �zޛ���Zĵ$�]`Д���#,xK�j��:
=��u8������Ƴ�=���u�"�XUݮ�q��nw����,S�� �;�J��W�p8���q�����垑�&3 �����݂�Hk·���A��|���V����aQ��\�*|8<�&Z.�D�v9�֋�	��J��L��VQ�?�_��V�1k\�$1�XA���>$2��u+��q.Od�Q�;��6����x��	�UC�������Y�� ���3�p���\H[3� �#�i4R]���I�+b\�Έ����
���"�#�{䌰\E�G����fp)�Q*GڭNr�W�W�z���y lchg����T�:[�"��2<Xt%�{:�5��{:�r��:/.1��I�����<��<9�a�K��q�����
�0��夭"��)���ȴ�(��� �Q���D��>�@��x�^y�����w��R�d�Q,NF�&��8FܐV2S�H|�J��lR_"L� Y]�N�K7\��q����+����C��R�o���ЭST:q�h����G����#S���km�0�k�ь��_t�=��$���a�Mct��s�I������Rܳأ{v��G�)6(�:Z���7f��41����8a�
�6{����r̴�/�$+��5��OrF?�u6c�K��q���7O.��>W�-;���<,�0P4Q�D��^K������810x^�*��x�+�OT�o� �G�z��Y�^��zU`�3��y�I��ӯ����?�/ΌO�t#w�=m(��QJzI�"��Oܱ��5����9ȶw��迳d������������Ʀ����V_k97k�'�\�+}����M涠�r�`�I�`��f�ӥd��Pzkf�����#����S�g+[Ue�|P݅�}����9Q_�w���l�fI�in\�����?m���-p�Ic�H��&[7g�n�T�O
��P��^9M�Y.E�,�k��O@n��%��/�;�|˺8�:������ι�l'����6<�oE(�G,�(�2�f_g���~�}T^G{��:�wo^" ��=���%տ����hT�%�i� � �qĊ=�1�.@q���=~s�!H�k��Jä�����>��&���E�"���h���o[�D�7'�f�7�k3(<�+�OO�m����˼�gd8�t���K
��o��x&AYɝ��P�J�	�*�����E&B��j�o��b^\I/.���B�"I��Y�u.S���p������,W�۹Q�_[��L��
x��\1^����E}��,��|b��D���`pIH�q<Oe{���k�l$=!}�`�q4�!Vv�;m6�u��g���e�B�ݲP�!9�������, k�*�b�z���
��-�6��<�u��Y[�3���,KǕm���w���\��;�m����1�A��u5}m��|����F��b��x^�"����� 5c��� ��?}A,�CAp����S�,�(H+T�ze�6�ڌ�
�֗|MU?Y���^�"�����h�p -�61��~������_`</<���B\LnuW�w�V��X`�&{_Peix4F�R�IM�(W%D�g��D��dJ,�ܦ�&ߘ���#e��%���Ι&����8��S����� T�h�)�ePϔ�a��H@²�D?�>���q�go��	�g�W��<Խ}X��0�������`@�-�/���8��V#kj��j�����!�<�o¶��"���{�'a)�BB�9� s]������,2SV�3�0"~�= Ԇ�������+ci����u�=�^�,�*n����"=Np,&J鍘7&fQ{��,�m�B^>�}�̧�-��_�|�U*~�4f���6��Yބ%�_+m����,.��a��`�Iz�¾%��C^Dn��(���	=�4�1�� ��P����aV���Pb8c\��Aʥ��5��dL/�Dj=9e��77/���Na���-��� �ϳ0DB�%�*�����c+���պ0o1�L���q�"bٙ�A^n�I���i��mXX�lц�/�$�������F߬��@��ʌr!�E�H*k�Bk�%��	��{9���£r�.	4�����*�ƫ��I�X�r�d�d�MӆiR1��z�����N� ���T��1"I���h�s�c�j�D��(��a��E0&�l��ğ�|	�8�����|C��6UN�b[Ǿ	�L�ۈ,Z�"m2R��zh��G�WX��@[� ޗH����ր%c����dJ��:�6�D�(�B���(�9���y��m`������Up�|`-���]b��ݎK��9��ǆ�/����Y�_��v7+��#�;o�bPQ�f���t�f�u�h��Vb��7�������k��+
�k�M��ږ@1�TZ؈9g_��]�"}9@�v&�`�h} �K��6���kG!^V����ۚ��F�G�Ҭ�A�N�K�㽔I��*G6��h�-h�`��M�W�=+s�S�BL��	�LFL�]z�k��!2�$�3e���7��+��@�����#�y'�G��Ё#�$7]� �C�"<E�+�u:�x�>o{p'eԀ<d��3Pqd���E���8�:�W����\L�B��"��s�M�t�J�c������D�+Ṛ|���pA˄u�K(2\���X��b+�Ң�g�m��]�z��cU��_k�t9Ř��G�8�qG��}?ɝ���܌>��9��4 ejO���S��1r�m9D��(�P��[�8�6+��}Wȃ�3�(��CR��x���@P&���u��yo�"t�%���
VN��8ƌ�afؔ;��S��� [�襱.�G(:��̅��" e_��o,B����Em|U<ݓk"�qs���:��*Ԍ�I�m�ʡ�����o1~�"L����$�1�9*�E9�|�g)^�RF��W/ے����[��sWT�������]��/᭎��D@/�q�݆X`ܿ��t3*�'�ܚ//�����f��i\�������]�8L��i6��aކxK˿�qb��,��1�p���.3����!��DU��œs{2T��BŦ���(�P�~jڡ~���79��s�n� �d���T�˪�(7�{�o�N/#�e@��������!�g�0����
CDa�S�L5�@�-; �p�HF<�r* 6����Q���L�S{�ו��CÀ�cW*����C����A�q�p�-͍���@���2�QIB(�J3Aы���g!��\��&SG��8�c���v�q��S���ՠ��h��JX 7�E��4�t[�P����	�
��[���PAP�=�4�S�ϣ�|�|�Da\��ip��wE:_��Y?�����~K��s���*x��&�Aŵ�T����cN�JT�y����,de�o>�^`��<��ݝ|�pؠ�`�q�u!(�M!�Ɍ�ɀ�o��)P����g饰8�sOa��.17ݚx�d>�^j����R���FK�׼�Fa���3��y��>4vLXX��E9�B�b ����Z���Qy�{������ �4?溞!�{L&Ql�O��3w,XZ�hv�!%S l���k"����Ńţ�]޾p���$&�['ͬ�f̧A0c��(�� fRfJ��deLr�����=� ��(����<�l�����ao.Ũ:e{X(3�5r=O�*u�\(?�0���c�l��������;�5}V��U��[i}�
D;[�����ʷAݗ?8v)?�o	� o��W�ȵ^�ؖ��-@.B�����^Q�\I�W+āG������A����_�۪/��?wrݚ�}'��=���@*������k=]�mD/��*�i�~�ܒ���U8c���xg��-z���+}���+������K�A����M8�Iޞ��mg��<D�Bl a�Ȩ�_a)�5����9��Q&����a���SbՀ��pF�������a���S��˹%��3oy����c�S�����-�z�����}|V�L2BP�	�%V �ҏ�w�_uC����,a���l�ps�"�D+Z�I=Am���簟�~j��N���ZH����%�ρ!���`>\�w��s��@�D/ ���< �f%qR�W�L�C;t~����.��������"Y�+ߤL�yw̫hh0��V:C]���}���o��B�S!�z��eFs2��1�#���q>�^"?a������]�)*�/����Kb(��PV ����UST
�wq����t�%���p��=���!��b@�����?=]�~�3��m��J ���"Z��ե�=�?���MP7�H�9*=�ޜf��;�<��_�����f/Y�u�ς<[*9®�gE��L�K���,�)naK��^��Pf-�w�g���"ӧ�QblA�Ӭ5F[�|m:��Ys������"fq�bJ�c�5t ��U�)�4HO�OxB��.Z~ J^���P�52�)�U0���Ic������Dk����<:����:T\���+mUxig��h98RHO�o�}"1_���s�?��F�(��P���Z���
�H�.Ulī�og�	��!��>��#�Y���b��iYȳ���z�˚��%泭Ԃ照�:�/�m���Ƶ�|0��Ȗ�U	 �;/�}~���G^��� ��x�?�Ӧ��*���V���VzY����m��6�!� [� 3M���'#���t\�Ȼ�R�tC�b=cՀN">*��s�����Q�a��<��М��i�Cĝ�ɂ���Ƭe_�F�ݸOiK9�]"٭�o�_W뼢�첛7mb�tZ�����֧r��:����`d�JS�%k
�� �J{ꝩ�/|��:.6�7���.lˊ�C�E�A���?�U�f�9�����t��j��Le�H��vS%'[�	�W����az=}��^ݒ�j�R��l����J�ҊiF�3�h���8I��Y�,����^ԬD�5��L���j_	3
�N? �%D�a�TqL� �r���8� <���]�3s>$���z`��8�������e�[I�H&�eK�sPRj{!�$�Ê����1{����À�Zښ���%��Av>?��5�>(fq#<���O�S6���7�N�]:,���{�_����!��b����\�g����{��r���k_�ɳ=td��W�m�� �i{��rg�5l�n�~C|�,�tV_`��*����W��G���e��/�`�p\�t𪵺�i�@Y�]bWFA��s>�(�P�ָH�Zۃ���	�\�f��P���`T� ��w�~�g��|���h]�d>5T�����;���;R��1Ecߵ͆�"�Kٮ��*o�ϫH�s<���7�e8��TV&3�+��=8�c�z��-#��%S��߶�$ֳ5��ir���1m�J&���*��`2N��Cjf=����F�r���>X����vFj �hE#CLL�&���R|���L&�WZ����ᩬP)Da�}��)$��팝׸���Њݐ+͆D���v�f��:"p�A��5���,��ps��S;ƼT,sSXK�E�Fh���B�K�l1����A��r��HN;�p=�lZ�0BE���@�$dp��Z �I�V����SN�4�Ľ�x���P�#(�>�>���6@liC�{V�TQ���;*Z�øb��~�,��ƛ��jrx���\r�V���}8�s���L^�X���$�y�d/ ��տjEu;"B9��C���9�nZ�sM��ݕ�c�̫M�� ���.1�i��"�#)^(?zAa �J�	�QuzFz~�r�G���.	zȟΞ�&'��L���Q���}��ƽ6ف>f^f�%��6k��;G�������Z�x�KN��Ǌ�� �*O:Zg��c���J�X����ID�Z���O���E鶁�jeK$T�T�"mc}TM��[��hՄu6�')7�nX�65�|h=W�?�,���a����fX+,f�:���I|��x�,A��,y��'�n�8ƣ�?��Ctm�����,A��:iIӱm����D�)w5�n��t��Ձ��,!�%��]����x�έ�}6�-3�q�~�9;'[�A��g�Gt�� ������3a(uW!AU�z��|�P�r@z�b���N��;oO	�ϊ��ؓ/����e�C��R�ӗkRY���#`n��.�k�{����ƦM^��k��c�~��~��L��o�C�G��e7yL��H��5/q.Ra�󸠦�9��tp*�u�0�i��@c���.07+�ot�Q��<ցXIՂ�1�"��@�9va�o�����A�)��<xwx�$�^�,��8� e��L���{���b�ʣe�`�4G�v��o{���,��Ӫ�2�����L���̇@��q�(��7���複����uf3���N`����m�z��e����%�M �)�&�"�����0�Ռ����!1|�+��t6u ��! ���"�f��MZ��	�﨡�oZ3R���*��9��'d�jD�W�'��	$�3WىД-B`�f:����bz�Go~q�Q�_�h,m%Ho$�z��i�M[%�T������`_���3�F𧏼��'�����u����z���d�rnR�?2�CFӋ�c�%+"�?�U�*<��<�l�#A�����E}Ѕ�p���L�'��4aJ���I������ű�
�>^��^�Х�7����������)�B 8�
Cw8�U����v�s������osS~�A|�+�u�l��������g��P�O0Q�6X�K��$(�c�iRW�0e[�9'$�b?��A�6������q�z<�&,�K�h�V�p�oS�]�x�b7���W�.63���9��Z�rO4&6�B0���OC��p�x���y��3���@2�ܪ��<�q��j��%f�$I��u���|�=� ��ZzUf������='!�>���ii"^z���k!�c�g@�K���V>X[���Gc�<P��=�N��p֠�^s�vE�E�N���iݢҵ�0t�b020�׋W�l�o��`�.���m\�N]�y��J������{L���#��I0�ؙt�zP铤D�>w�\�}��Al��l�}1����8�4B]N��J�~�}��A�����p��@�/���6�<�=�zx�O�Wi��I_��Y������x�mu�hFz���E���TVջ�����V+�܀ ��ɩբ����R��^��$ƪ0J�Q��N�5?q-����^�);�v
������2�+e��-����ci�#���=p)yuX�����Q�U�}���9i�i˶&j��d�w�b���p�Gz'��a*\vt�B�7�����^ߵ˪��rw7bPM%����X�ŝA��J�`�or�(a���Rn���2��2iSNv�������G#f��$�*7�]���M��bR�S�Z�ǰq<��#u;o࠵SR�����Z��z ��]��>��V�F՜q}�^l�}ʋ�u�Y	��uU��1�������ʶK�])EE u��]��/�;=6�'V(�j!�*	�/�v*Nŝ�U:;̟E��Ĭ��VP>i/U���0<Z�}0�z`�����R�/��@s:�h��Х�F7(�?�%D���<U�����?�g���PFF��|h��q�Sև�8�a���tϭ�X*������dh���\�<Ź7������9btA���]��Α5�c�b����G'�T\���~HX���T��>So��B5�Z ��
�'��W�$ڻM%�Q�A\�y�S��cF0��+��`��f�u�o�ڝ�Z]B?F�rV0@�6�p��#@?0:Q94P��Z���LԈ1m�x�_%�zGUk�����}��|���e?�/��p�gQ��ཬIn��͖K����x�{�@m󲎺Ϝ�B �3\�_����� ��b[5�T�4��XJ���w�����32(�L+��<����/T�R~��ކQ�A<2�K���DزB	\ �Ϫ	�BK"B[ ����D��`��VM0��e�ͣ���fE�Ϳv�/3�>�gF�ACLy�wǞ4���@9���L�%�_�&>4�e�ԥ;F�ݬ80^ЉG��ܗ�M��j]�^�����3������aP���Vz�+��.���Q܎?2g}��j��])��j>ZqKoD�NRV��;�W���yA�g��kKM,��Y�*��G�u轙���I.�~�.�m?��V	� ���v�U�;�Cb���+�tI�aq�}2rYB\X�z��9�@-x�ty�c���a��e�`�4۠�<�'m�q!�FoBv�VIz��Z�X���>�%ez�ik��.^y�F���}w
�0<����Kgas)��F��O��PNۺA�������x`�l�U�)!�A����YcjR�lS����zݺvG`f������g�o�2j���,s���ki�����i5g��O����9c�D�}��%w����>����?���m̿c8a>�nB��o����u�]�����K}�ҫr������S|Ne�ӱ�Q�?]9:�m��Y(�)�~%�S��/���fB�!p_��`�݄io�$|���u|"��TM�"��3x�q�tby �
IP�In+A��%����,+R������72��-Ʃ��~�#�.(����O�Z�t�C�ү�ԭ��1��)�ۧpqyrs`����*���szT�к|������6�֩KՋv?3y�GT�LX�v�0���j�Y;\�v/q�E6�?������ߍ���5��/0mc��O&���52#�{j�#�v᪵�WGF<�.���,X����:ku��+Z������j�,0D0�R:X�s��3�Z��6�1�L��&_@�#���xYDz�:|��!c�m�0K��a^�G�щK +֙#iL�;{%�,� ��eJ����e2`��� '��gt�t�Y5��M�r��B�p��e+��<O-���S`|-AE�$5 � �H�K�;����T��5@H��T8Ee�Tkё?��!��y���0�����q���ˋ��U�RyT�	�%hh;t�8�dP���j���S��A� k�8p�i��^KϷ*�YT�\οnX�|D*��p�7�ӂ��r�5�*N�zЉ��*���2��e��1T@�%��Zi^���t<��M����f��{�τ���V SM%�)��p�����ڵ�6
i��`�L����m\b�!g��������6:^��D*3�:��s��^����ɣ�q���µ�����
Bp��`t��DK��wƃM"?�����)Z������<��k�;��+�\y�	~` �����c�XI��E���kN�vF��w��� �����*9!<�H���{��{���-��I�&���'�a���XG.�JO��?�,`{�YT_�dM2����oM�ꑠpo���{
^��L��}��^c�ZՆU~��B�E�Ii^��m�F��Mk�ef�+C�T��M,�;����)�FG���W3j�B����T{�T�T����\u[���7��{�N���o$�֓��q�S�8��Fo�!�����`P�u��[C�*��Ch��K�k��ˣ2D�����4U�iu�/v�%��=�r�%;]U4�"4Z��b��� ���ltk�1�%�s<���)��D�6���gC]Se H^ U��W�7����zKރ���N�E���'�T_�D��h�4k����(��{N�C#��9�|��ה�[���B'
r��b�c��I�����+l�,�˛�:��J����+�6��RM;-:�;l������Q)���[.85�Z��_D��D�{��Q)<2�re�g��� "���d�����t���Sܪ_tM˟��B��0�Q��O����|���;��M]D�r�U�-��eΣ�nƓ�΂�f��>N��y�Ί����,N��#ѳ-
�ZHPR�N���E�~���?fڂu�z9Ui"��u�x*�7�����XY��ۀ�(�ȏ��F뀴Q
�TH6���o�B�e�Z	�
_�6�GU���1R�Z�k+@v�і^�A����L�ؙ�V�d6~�=[[D�d��(W�6=�ف�rpo�0Db�ht���q�_�k�=w�楆��s|s����%�o� ZK⣻oi�a�3p��t�wh��S��>��y� �"�s���wo��$ڠ�����E��X�6�'�ÈE]��`=�K�QYR��8oR���~J�a����4Y%�,�g>uH\KX�a�9�����^�έ�p��^K�pEζ<���T�eܴ��c���^^�@�p�Ʋ��A���Yt�[>e�����91��}!��Sty&����a-]f~u�*%+�%Ԕ���n�p/ٮ�|v�Q� ^g�) �U�y:�j�>Ag���Du���\��v��<s�c���7�'�fƂwn�1����D��$��̈��7Ԁ����l>�DHnQ>�^�5�1.I�jS�k������Ʃ��E���̋V�i��	'������p<u-��h�`��U�r�YRG��0�<H�G4���ڛ�|���(
��m�bx�C���$1`�=�'�]%} ���R�#�#	Hd��y���t>�I����v�_���fy���S�zj�_����J����^9x��X:I��Ylf�[)�[�ΞJr� 3����Ļ��ql����Ju�ʖ��B�1�0��;��#�X�UE1$�E������%%φ�2N�P>=�[%[�|�R���~X�Z�p�����U��/1hd+���((�-�/�����jQ�@��:��g����6��in�;ͩ�v��9�
5a�@mD�*C�7 �kv�r������s�qYGJ�*�l=�REK �Q��8��;ۙ�Z�B��,>��P�#�8�8;b�"�}�CL/��O������A��G�<p�f�����{d3y�\��&4��{;B�Iwz��P����H�g=uu@%E�+� M0��}-+]�C�-l���*����� {A�Em��D�����zOC_46 ���V,P���&�9��AӀi�I���Զ�����ߧ�ZW��Тb�����؊
���eQt`��]&W?N5>�Q������J�o��	t���b�<s)���f+��0Q��(�I8�vG���݆4�q�W;Uf�n4���[�� X�
5�i�R"m�>�68�L�6o�D��9H�e3���R�N�^�D�\�	�m�p���" �NA�wC4�[�4��
�r�׵QX.��om�/ə檃������;T�����T?j�yEN˔��?җK*y������ܖ�����b5")
�lL�	 "��.բA��A���9b���?^#�3H"����SkN��~=�]M^���c��үL�Y]E���xh��qm���t��<~2v� :����A�͟&kS��R��V�W>T����k�JX���CQ�jE>L���6�8��2XH7��u�� ��06�ι�H�%�����R�^Z�Nq 혺bO�ỹ^�������ܜ f���j=�����.�<H�O�3�KA.�U����}��l�D1't�߁�X���}>J�s��
7cN� �C�(Ӟ׈AO��j7�,2gO^�`�5w$�:@�Uֳ$F�2Jc��?S�w'Y������UC��9���ي��/ݣ�!��aP����v�ٔ�gfH�[��ւ���``9�o�/�/+��H^�����o�anQ�6����t
��d�uD1��9�Z���@�&f�Ix��������i�ZB�V1�;����c�>1|г�.�Ӎ�J8VD�ŝ� �6 @=NYXa���ynd`�j��'����Y���ǽ/\��n�!<2��L�r�i;���|��h}�@�����f�AS�k�Rls��������]ǔ
v����,V/s�W�0��BB/{�l���'^?MX�ذ�~QfE�����6����x�d�1�툉�,����������8�K�g��G��+6�N@C0�jܓա5�"��B����0'�>g��ȟ������c�ͺv{Ru@ݸw?�˻l��*��~�֛製��lM�@��1�I�Z�~u
��<�|���'����d.l�h����f'�T��;��4 �d���4щy
�w����E�=��LY\j
�R�7H�W�>~�WPm<���/f��M�T>��t�4��	����r�m��M���D
¶޴E����x�I@7���t&�b8T<�e7'�W��%�?�w�!�ޗ�9DH�:�6,l�Uo����j�Ro��!��P*�YI{"�v�c2�l"̻㚔����V��J	����A���#���_t��J��\��ӱi�D�jR��w=��jk�P�P�	(�,=�u�[�"U���QѾ���v���t�_M���e��_pU,�;���T�m`61sb���[U� N�3O][�?�_g	T�x�E���|[��Y	�騹B,�*��� yߟ-5��qd9|m����!�����8	�T"�탬B@�� �	�����ǘ��(��u	����8t���pRcj<F�4:�y�����z�Tt�i?����	
"H������Q���ʌ������\���L�rN����W���]Pe~E�8<�d���z����?ۼ6 ��_��9���=[�h.�-h���=�v)�Ǵ��)�D?�N}������O^�ؤ���M��g�0��᩵u9�-;cT;O)%l������ǩ�� �Z�M7#ް�}��41s�1���*�Y��,.V������<���A��w �$�U?�-&T#xJ*�21�&r�݉�J�y�R���)���X~r-`;X���6�_��R�!�̫�$�H���,t�1t�a�4zч��x5�t_Q�f���_C��>����@�!�:]#�'�;~�Z�[գ�4��x+��۾����.
4�~��G�6s)�!�4�aJ��(��g8o�M��l/�I&�U<��ؿr�b�<B��M��׎RT\ ��F�9S�
����w�Q�Acé9V����j�{O��٧b�(���:�⪁1���h�>��5��b3���U���8�vvѫ| �� �Y����5���7��k(���������.��f@�?��d�8Lq��<ZYxP�H�Ʌ���=E�e`��Z��Vv�w1d!���y��wX���y��|C��b�Z[b؆���h�6��Rb{i y@�4ĉ��8X_X*��歁�����N�ag뛚�%��}����F�O�n��\*�E� 
��5{F>,(Ge������Q��SF�Dϋ.�j<j,���=f����$��Vv'�!
]=ڭY k ���I�Nixy?sCF��lm�Y�YZ�p�r�E��]��{��L���J�J&g�\�0��7f#l�'<�4������g�һ��=�|F�SI��-@Hx��J)�ɓ�e�)c8T��m�?��ⱌ���囩ݓl���W˰qyhgb7.ң���#2@*D
ׅC)�� 3P�>ѣ٩Eȧ���J���c�C`s9̲
���o[\�9b��@1����s��&^ ��C�Y�,��4����-�q�v\̧T�����͋�.8݋Il�O�.X�����}'@Y���!��O�r�	��[�����ΡN ct�����'���[�i�;��b�r��'���ė,>�!6OH�&��N�t���� f8�"�R;�r㳹������$���)����0fؾR���Z��8ra�bN
���4=��2N����s��w�㭓�*�Ę+���\����!��>�Q�'kkV��2!@�cs��z_�I�ν[��ޯ��u��1��ܹ�an8�����"`6��
�<��Pf�se��K�F�/_��yVxj�z��#Hv�}��B� n�M7%f�����r|V3Tj� �M�>����_b�+�"���t<�M}Q�Ϝ�0L(�W�b�*L�_�6�X����ЎB���.�� -�T�nxH�ρ��M���y	����ј�(6�mE�Ϫr1��9�ۼ2���Ghx�\���,�G�q�<PǱ�Qp�i�鎟�:F�ښ��1-kǧ��?��m9�0��e8�N��!�����	4�͙�*��������|Ëb�-@�N~u��I�-Zk�³���k<;�vc��i�gY��,z����P�L���W�����&o����50�:����(��'���Y)�`�<��Ci��_��8 Jh���xζ).�Se�}���+�^���?\!h8��r������$j�����h�h<$K>�����㟌�RC~��^���VW���r��S�t.X�
/�18�\���,�3�N��2A)�QL&�f�&�b����P�
#R������Y{n�����D1����>�����2��C�#�����!<R��@bBܔ<�Ԕ;W2�1�O��RY{۴�����Oq�r2K�̉t��� �0`�8�*,�M�Zɨ0�%{ '�q��&|/8�Q����;'0f��[d�ER�g���^f9��t_N@��Fs��#��i66i_��ºvLND��u*�Ɯ����0��b2�K�vKy6�U�y����6ӮD��Я|���h�� `�5�/�ΐ���[3G�;%��eQVK���DF�#�RC�0�V�b#s��� ~�����C�z�i�%�8!�dܗ�č�'ف*��o/^V�c1�CRj���0�ǵ�2�X�V���b�"�,�&�j�+�"��y�
 GpZ���agnt���˩���@��$��������-��x��V���Г;S��Ac�8_�9�`�2�cyҫ�l��w9Y���%����o}��\�#.��3��?D�!�oV��ڭ�����=���=	�P�\���I�i�x�ўu���/֘v����ֿdDm�0�a~���x����J��H�������+9s�`���YGO�����t� �������X����by�b��Ma�u��P�;z�Z'B�KQ>U��%pHXe���W�~7�Ďtv�{O��6WǸ�R��n@��}���$Gd�8"��t�'hÓ��߅�dQ;����s���4g"��!1ܶ	 �b1��P�'��h�"�Ea��?߰�e��s�E��x�5�I�x�B`��'��m��w�����5�;�O�3ܙ֔�!:,Z(����e>'6X`��������[�j=1�P㪘͆� �d�0ʉ;H�(|3=���b��k3���_&�VN�X������8�T���8����\e������g�BY����ţ��N�C��"NX��?XǕU�[F"qɥ��i�A�|�L�}F`.�����n����l8�T��ޯ�6�1�[UH��,�J�߼��.�J/K��?w��f��,�[Hs�"p��aR��!"$�����.�]�^�F��k*[L�c��(�A�+�[-��H�������o�C�-B	�(Sf�g8�v+�F�}]�W?�v��i1����ڠm۲���c���y͌���1�2��ɐ�S����9����=�z{좳Q�Gb;�u;�����.٪��}�&���L����y�:�2㛞#y�k��ř7�� �5���dQt~?ŋ��!Y|g�R�Bi
g�d4j�ٔh�R��Ū��A�i/��o�����|�J��C%�ݎi����=7z�F�Ĥ=���P�V|��%�c���Vh�ѲwOg'|�0Z�7٭?^���5�üfF��O�6���ȣ|S8��2"$t���AF���&2S+��<��0��'�U�(�] I���W�'�1��{��l�f�=�#-�r��R��IdG&]sN�
 
A���4�P�����cv%��ы���>���)����/��	2��B-h�OÉ
�q�O�^e���B;5}h�v��c+����Sj��*PCX%��xIK�k�
j?:?7�5��3��TP��K��ȡ���9�+�n a[W4���Κ\z[�"�i�NY�S��΂��G킭�+�H�;U31�':)?m�=ԗ��ơ�L��iOz
l�=��1�
�Qg���"+��7�XEa�R���9	�D~Mk*̒�����x�9��t1� ���,KqG�]�E~?z�*}���{q��/����V�Kǖ���8#��$����N�<�*]�����[�*g˘�^1&�O(��3g�[1�l��G��xk�2�~�Q
��)]C��(Kk��{�X��$�ߊ�~��*��Ұ����f����b��䂱��Y6�Ly���=?��Ma��I�<��EeKՋ:�g/�+dy���]���~{[�����n��;P&�j$u��I��;�1��
�w=O�����.�ft�{�^�f���g�)�Bs����"�7�j��,�= }�SWoGM2�#h��S%���A�2>T_����}]�� 5\��Y�D_�N������NE�N ܦ��o� �����3�Mߙ<m׻�x����K �dai�p�|D�f���g+��˭:�P�|.^[v�q�o�:��ᶔbA-��M�D�YQѽ��DgY'X�>V�y�%�-�3;C�	��E���/�W��6�1%�~��WQw�LA7k�x�� ��x!ۀʹ��m8*&��yH�34�i�*�����	q�1A�V�,oQW���B��l�^��ǹ�����O���'lM���O�ͱy�ת�0_M�/�_�����=1[Q�Ԭm��d��T�F����wZ[N������n���L�̐&���c�B���b/Z=T�Ո�]L��@�����Η��
��!�?��d�5�П.YttA�(�gF,��=,�jȠnƓ֪ty۲�Z���+p$�_M]�0�ԁ�r=N�T���:�Q4�/���k�K��I(�����r�w�Qs�yL�f)�8l�i�H)G�ۚ�{�	�&�ݙ��V��]&�;����	L�m�q��>��lX��KBe�1>;vi�����l����5Tm<C؉�����B�7B`X���aq�N��wZh�,�,�'f:O�/v�]l�H��J�%վ��:Τ�~�=�#�-�E%�⽦�� �T�HXV
�{�>���zí+�2 Gd�t���7߬��*G�썼v�M���ؤ_a	�/�6Wa+]_^��n뤇��rZ.�����I�#��HG�n�y�	4@āo���ָ+˔A/�W�[�*7�L9H����1� �明�0IBʭ>8���_�㵕�#9_�m�ڳ��N�L�K�ET]?����e?�-�9�Y���|5s�='��������o/M�0����d4�K�L�(�@�t��!:~�O5��]LD������_]����qp���IֵoC<gj��O���o��M��a�U���f͗X ����y���\��"�G��s������a������;��C�m�˘h\���8v��C��a�u��`�+٪�T �^���x_�cB�%�.�Vn���9v�%�ᎃL=w�� .*���]�v�2j+nR$�b���ɖ����"�H��� #����\��|��xrH����7ڹE��_�,r�ƾ����}	�������v�;����<���8a�(����'7����'(���%��j��uk4���5���K֐�� PT���ĤJ$�.�U��m.X�$�g�g�]�;Sw�)�}�dy�25v�U�P�:M�#��#5�Bpٵu&UY�P1�	�U+�o+���5���Ӗ����=�J��X��j� �N>ٖe�p�,^K>Y>��
�ܜ~�D	�SL������X��H���=��!��o�f��P� 	�,5m-��C�%KB�ǔ߻q�{�s����x��b'G�Q��|�p�+a'�x��59��&��F|�H'_Ƀ*n�������{]Qj�://r\�����
\,iό��<:�)�zAdQ��5 ��o��i�������!ПS`�fw'�q0�wBO�5����_N'�/
j����c�'�s�m�)>��ג|L�Jm�D��S�M{�1\������Hv�v���>���d�U[tZ��N?�
�� �}c�	>%@�h�1.�Ak��n���'�"�4�)�~s�o�vU�A#I�i>"m"��dО���@c*��_I�N6���G�deyC�ˬ���B��Q7ALyr���mN�aΣ�]7����L���6I�VG(���I��]D�bv�~�g�������+�#�t�1H� 
���tC^[�BD�=���u���*���?Ф=��͂e�^f�{IΦCA���M���ÓB0ۯ�9ֻ���[�$�{μ� �,���2���h���v�I�&�D����Т,�7R�����_0�Ȏ#|��)��/4��ay�Ǵ��Z��c�i�ࣣ�\�{�b�io��7�^��`�����tև��O���z���>I��(��I.ƭ}�SS�ꑶ��8+#2�*qr~��D�����]"�>�ۮ���E����3aS�~�.z�I�e]��jn�;�Gtx/��RG5�����N�h��#�-OQZ?��
ծ���!7��?dFr. �_���.Xߑ��I��p�Q��-���ӷ�C���̒�s�/.�w�h������u	�dO�%e��Kiԡq@�!���!�%J�'�l=\Du�=��ۘ�rA&��c��y���K�N���z!�s�s�Z᭒�LOs�Q�&I�$�T��zop��f�+=��H�%f��bo(��X��a��n^�1��Ȗ�|�Z�tZ^����En:Pjo#���	�$ɍi�ĤV�ک4ɿ	�}�eb���k�L�* Ql��?΁ʹ���+�^�W�Ťv.A��\H����*���֏F��o��U�XX��C��yt�$��	�2+T��R�I�ar=�+�ʴ�  t��^_^c��� �,P(�����UL,X�S�4t�CV���Z%�_فB�S?�Ծ�7���mb��>���M�VY�*y���v�,�,�s/O�
�D��k��_GC6��ު�p������1ҧ�Uv��I�葅�R���\iU���S���,���"�����0m�O�J��G�7�������T�bTg��8�$���|�o�y�Ww2%�a�'��a#��6��n�Qp��K^H�y�� ����	����r�����.}͇w�+��r'�]X=E_��<W��\��:/$[U��_��@@����b�<���o�Mi�/��>Q���_F����6������*�D=�����<���̘��U:��I��^���c7�ʹs�ߟ�K��?.��- ��e��1�PU �D^�Tx���0C�b�5s�B�>S�9�u�}�0P��ז�D!t��w������d����^n�^>jKD\���t�S�y��W?��P�_j��P�v׼��(^)�0s���lN�B��x��m_��V��Fʆ�e�؀���ZΔ���3��#�_��W�\q���i��}~"�c�������eH�8������$1�Pn�}4�DB�c�X��-��ˬ���)�� {V��XQ��=����p���*" �`�/6;b�ͱh��Qť'	��jM�O�Ǔ�aV�\���3�u[v��f83P��h��9�]�zC(2���XkU�P��&8���vr)
-�<�q�>����|'��}h�an�7��)�M�(����ȓď�Ә�r�6�N��A(\��wB�����鬓5?��V�@���]e�^f���w�5E�9�e��/>�2�1d��|N1� ����AÛK��D���=�8I�J��zD/g��1�%;p��!����ǹ%K�^�^�:��F���8�x�F;�D�0�D�m�v�=V�4K����=�;|��T%���ڈyD�������J�+W=�z�~�3��v���U�>@v��	BT�N�O]0��RM\xͅԎ�z&I$�O*������\$������k&\��`��aH����	��뾪�	�H��`V��q~.�
a@6b�&Taf��A�{�����f��C�w���������j���%P1٫	j����e���8���b���T�(��Me�<N�M���	e�(ꎍ�~9�q'r�4��O1�v���Hm.�/����:O	L���Hp�|h�/C�b��r����H���Ens�k�9Qs�>�A��ږ:����Ї0���t�{x�:�ј�.�0����WN����6�cF䚑 ��"):�S��X�m���ÅV*���}��I�	0���t�R����R)�̶;Wޝq��T�B�#���J4-���?�W����%�{!��_�����>Iy�����pR���Y욧7WDn3�~�CB�RB�XYLܾ`�9Y�/���w~i�m61^jl#�u=g�zZ7ɩ����4����R���Ia?�I��#�'����$��92�G�<��'��G�~-��ڧ�=eNnC����N?����<�Ε�H�Iܩ��^C����������{$伌���ZG�d���[�� ���SFc�	�������0��+����#$��a�ʠ����/]D�?�/}ko��OTT�2Ř��<��i�/W�Mo���"�_�5�M�w�/'�M�?�5����oUF�y����P��7�P,���B�y����J�`��Z��kCH�3!���h�z�_�P\� 8�jj��tD�/���ALS�ڴ/6 ȁ˗d��bC���c�z9������͓ �'PL$Y�L	vHf�;w���q�Y�2ZjI,$�d��[��鮿2��Lm���H!�0�"	���(Lе-S�[;kW�K�(���Yi�9�Ѱ`t���kU���ʩ����V�s2��L�&\k��	3�y"s��.�h!�Zs≟>��{H��O�{9��6��b�D�y���$�!T�(0B
��&���Gd�e�mw�8YD��~%��q��\��䱧"��S�` 9���w��0`K�変��=�� `���ty����F7��t=����#-z�ew͆�X� Bŉ�Oѷ�`�r�|�(�����u��%����EA����h�qü���5śҸ���q�$�
�ʿm�~ojI��R�e��*�C��*�[H��YRB>�����6)�!�K]8���:����C
�\�SuX�h���+�Si���
�rd�|�L�h���T���˧�,��*��.6�Z �*y�I��s�Xb���|c�|Аh��w���u�Fl�H� b�,�@�y�����p��{c.�	Qeu��[[�9��:Ml]z�_%)+%���n�tb��l}4���dŜ�����]�J��Ƭ^�s��u�+XPn\���5��d<:h���0���d-8'9�vU�ެ���#"V�P��
��=Gg�M9�z}��8�,�'7&`Ui���(�K�Q��e� �K�x�����+��缲8�j�F0 �2�(����Fi!�`�r(l��h�&2�P�2���Κ�c����5�<�w�	/D@7Ix�����Ԛ�F�Va*�����t���3���)��UR�����&4���s���k��I[i����cou��~Ј�?�����M�S@���n3d�y��A7Q�G���)t��}	��B�O�MٌD�d����࿸N��L( ��*P�6���g���g���ܾ���C9��D�'�{}���w(YL�O.;0���{���56�ҁ;��%xb��b?��Q��w��Ьѭ�f�+��yd�>�B�>��lf�.��!�4OJ�br��*!�x�j�[Hȧ`���B�6`+�MpǅǊ��@�V �evh�Xl�.�؃_b�w#�<���@�@������֥5=X��aݣ=KP1B�MwL�7Y���N�z��p(�K��ٮLߝ��B���R	�����/0^[����!i����R�Ɋcu�#3]���?٬"1	8m*�9��r�Ǹ]�n`��,�	�8%�l8�eaPĬǨ��!g-������s�W�P�|+A{��/���PK����� �Vgꇫ�XhҴ_�$�Dω�h�b	�c$�C��a�Qf.2yg��l4�Ah"���L%y����C����@�U<W���M�~��7�����H^m��P��:�%����4����&�q?f��ş&��͌~�}΂L� +P�$q�<�0 '�&3N��Z�C�4�i�t��| �F�A1J�Oܸ������uؠ�g8B����D=��S���S֓I�9=�ᱻ5k
����$���R���"<����k��u@`]��-���xX-�d�
�:\�\4}���6�G;���l������m!>}u�b�j[�ZvgG�����i�
,��4�J$e�R��ϜNb�^z2�CX���@�م�0W*��ꗻ%���^��,��n�S<�ي��=mGPD�e�"��q�i����-/ѣ ����|gL	�z�K�g}?]��0ӣ��� ʬ��$%��`�-�Me�A�f���(L����5^�d�m������XP��)���C̕�LWqu��AsP�j���8eݍOq�_ޕo�[I�p�L����d��B�>)��/����M�Ϣ����l��<���p���/����(��Xq�dB��l��㦅�)H>�i���u,U�v�����"����ER*]F�5�m@΃&bC�7\���aT3���y�58�{���s�>����Ӽp��=��� -�< �"�>�@^ub�w6��~�4;�s�� EI_�����4!p%��i�r�!=���;�-�V�O1<^�t����=Mi����bBD�j!�}�G2>SRn�� ����E�V<�p�V����XX���z�B�?N|5=m�fu��� �W9�%���$=��Fw�s�
y�.-�S��8��I$�hP���qO� �;�����b�"���n[Ow�8�0���v���������_)������@|]cĥ
+X��"�n�Ц�E�X��:��.0$F�Bx����F?.c!�b�ܟ�'EZ�T��x4'9"���w13���u1{��/�-��c�����tq�,����	��? =�A�,iu�_lY
qk�+:��7>��}01��+�h�:&���B�Nw�c��RC�ש�9h��MiC8�'�|��u�yF�._�F��ۚD��rɶ���`�Gk���#�wb�L�t(~�>_�9;4�`����k`��QE�A�.��:j�u�A�*�[0C�
.�#(�49�q��	o,;6��Vmx1:(~jg�w#{2F�^�!��Z$�$L���|oUv��Ⱦ��#�p��YO��!b�{��#aJ���Rp��ˆ5ɍ�-:IVG�=v�Y5pV�N#|���3� �פLKU����m�rƘ>����u�J��q�.ȅ�ld�#\"#=��W_�⾛oG�J(�R���cqZ�k�ȵ��5�;��( �6�-b�<�,�Ƕ�*0Y�Kd�RR��s����3�7Q����Wr��j����}�r���{C�����&j���P�bg����Fh��	nu��	\'0�+��8��n��n��æ��:蔆X%��U��h�	v������E��X-ɐW����j�!�r��n5.�U��,r
��<;z��%͉�(�l�KaI��W��kB������1��];w�B]�)u����Fm�
�Bd�(]y������5����"�sz���[)Ԏ�$�o"]�|�{Z��rd<�o��X]k�A�Z���Tֿw���Rf���[��Y�_[�2�y����mo͕>��["s�#֘x^�
�aE�I��Q(��VPk}��[{G�?E�p]Ҩ�CZR�!�w�A`@/ܯݞ��)���說�+2�����.��N�y���S%��='�_����Ft�ae�.��j�B?Y;�� �$1���o� �'I R˔Ωe�G���?��C٠���YRBb(k	}	�D��_�W�+���$1R@.�w��(e��fNvX^R����˕��_UW��§��"Eo�M-�[��-Î��,E�Vk�����m;��z���>Eml>�DH^M��b���7��Fw>�s�U���oM<)�3���0Ez�ٺ��$Z��|Nv;�]xO�� O�N�b�4�;�*_ޭ�N����4�䧂H�y^�S�tА������2��h&�߅�!�\B� ��ˢf�?�󥀱��ŚB2�e�w;Q��j�ޏi��i��=˶7�*Ѫd��^�e�r��2�?`=ؾ���-���BG�Sl�(�J���_Q��:�L#)�
�Iw��	���+�x)^�/_l�����gB�ϐʲjM�l_���	�-���q��Z����;-N�_뺎T'�W��F�,�{V.q�ɋ������Z>Z�=�]DqLѥ��q�jnF_B8������%�������{�_%t�|!�TC��
5x_D��I�T���i�b3yd�^x� ��*v�	�@�����Zd�-7c]�}�����,X�M���D'��.�>+Q]%�kSCp�>����N�V�eaM�W�۹}�#�+D�BYf�l[A�Hd�bn�Β���9:n̪����߀qk��e��]Ԇ�:T��
�Y��"z��B%�R0��J�S&r�խ����#c^��F��9K��6�;*l�3�K��I��1��rGS�ڢ�!��}f�Q�BOZ.�����e����~�G��������7��*|9h�"��m��=j=C&�Z�(��(��wmZ��)�,�ɡJ;���o[�*2]���H��(!�~6���}D���}q��m>X
�����R�y!C9`j�|�����˯�t{�E��z�h(���T��ԍ�m1��(�!?�wG#�}�x4n��~������ؔ��&��~�kH9*P-s��&kȷ�rᷘx���i���#U�c�x�j9Ve:]X�c%�p������JJ�
�%�B�#!o��i7�%�>2���U}	����016,L?�*��^`=?{R줞������.52ne�#:���ܕ����J'��I�nNV���n���f�r�3k�uN#Z���V_RL��%�h�.��M&��2~gת$a��� ��������P�fp�w���&n������E96<�y
 dWd���f��)�*U�wNb�f'�j[fړZ;NT���X���%­q����`�����+�7���x�a(p�Ӛ�qw�V�P�kx�������%ќI�01i�kä��q��ߎ��B�HXkL�Rk	��&�vQ����Zk�)�jv�O�A��f���#�muO�(�@��*���K�M$J�T���K(�%kÙa��F�z��h�/.�Tkk31���>����v�^��i7]�3����i�����A����~�?�%-a`I�\!e�w�0�8>�P�U#Z�u�jz&�C�t5u���
)�l���7�$��>�z�:w��>����>���{�

��3Hzi�����^{5�/�؏y+�������<a�cG�g���j�Z<P�YُrwN�\�t�P>?���p�����~�>j��
\��B��"�BѓޒDs	�`�ge�B�r7�CPwN$&DY{
 FV)�dY���?��sr�0���\�c��X!�l�G�^ �ٞ~	�QK�R�^����(�iG�^_ub��ɜ���#�*1�VG��U	3�Re��#F�R>��S��3��u��;���<{]�*�0!��p�岩Op =��S�Y#��g7�m����8\5��B.d1�[ec�jfzaNm�	Rpl�]!OϽ�$�H��%k����+ �Ws�p�;Y�ܰ;Oer-��t�񷭳1Wq�S�(�T�L��{%��)�o8H`�{��%z�̼�g�O��R��@�XS��� �C���p��c���i��*����*�Y��8����5��a3C�w���զð�ы��@b�¤j�{l�.�i�A�@�\�2�$cq�N���������@2��.�J/r��D"�)䜪�����!�!(���d�61$��/�w�j(^�>(��Nr���섷U�社��6_��S�(�.ބ:�ӈJqSm���y��ƚ��5�s�����.37��Ѻi�}��L_�����	�CU��79�Q���`�H�d�|4��ef�h�рJ���9��'[\�V8��~��E-����o!E�q�
�ݧ��ퟋ��6?��t���s1_��>Eт�*uH2|�c�ʘ�cI������?_�
e��Zc��������$���0����V�A텮���|$���Ed�����r^Ri��;��=���"l���_G���q}{�����C��L���GA�0�_z�5�=_7��+��d��w>��P$�+�ýIZˈv�t"��������:,�+��kun��վJŸ�"�=��O\�K'�0�-w�ڦ�f\�2_KA�W�e��D���'���B0eU�x+ĥ�l�D�0��L_ա�������xD�h5�/�^C%�^�6�<A������B�����l�,D���0��!�ٓE�zNg�dǷh�鬚��r�^�m��K.d�'�����U�$��4�2ȿ-���`��R��f:�?X�e_�$u G����~HX��i#� ܃�4E�>	���OtǒwY�V�3��v�8H� //�E롥��ؽ`��2�.���l��L����r���+r|��$�r�:9�l�Qn�H�X5P{���_���A��R���/�$>;-Y��8,6u��}R�-�"ˁ�	h�q=�`v�jҥ��T�n^2@����E0m���5��ԋ8H�x8L�n��n'}���YZ���5��,��ޫ[y&eƖ�܂v���|r|����y�GA԰�,۰��-��Vf-^CI�n��a7��.%�I6f�ҳ&��I��`o�S���~B|���E�߉P�:b�n�U�;N�����.$[����A�T3f!鲏n'�Y9���T��ui��T�J5:�zl�2i*G3tqe����%��M����e��,@��.'@�ș�����{�[������x)N*C�5Vx��`�p�˵�<��4a�_� ��d�;Ѷ3B��W�X����<%��)���Va�6I>%Nt�6L4��D������rXT^;7v�B���e�n`��aIٛ�]�@o�Z�-yS8@�L�AK�m����(�PN���F�!�6^E���ρ�F�n�?��Rǲr�.VaQs1M`����>�����Gχ�>'���_U7L�Bk�;��o2X쯛V������ro/ݬ-�ɦp���n������9��� ؤ����B%?��9���������2�-7�g�#�q^b(BY�9uo����p?!cS�^�����H�l]L�*y#HEW���Q��߻1;
�^�B�ok��ݗ7��	4| �M���N�I�\QAZ�UB�t�l���ӏ=o+!]7$h� |�èI�
�cGX�����5}�t�p��Y:�x!t��Kb�<���}��A[P\V�?�sx'��rz
�tb���̌��jȟ#tX�Ӥ����9���C �����3TJ���^5 �vߌ$�%�MK��U�#�-��<��X����W)A�c��h�l�~����	�W{��a����KQ$� \#�_���h�l�x^lgWC��c�Ԏ�A�sQC�fW�.��W���8��؋��b��mj�^�I&/��70K���7�D��%Ҋ�'���B�q���-�ΐ��z��+~���ܲ*�\s�&����qs1�;�`��lR�t�^�Yއ�v�P7�׸����Nx��?��_9D�Y<Z�Ǹ�~j���n8ٌ���{�����`���'NCg�	���u�� �1Q}���-(��B˰�9�j�}�˳;\���2 �wЗ�;AO�"�&�kF�lۧpaDdB��17�g*�st3J(C3m�� +�7K�'���׹���5�b\Px��<U=��V����9:4���ϫ4��f�쐥d�$+��<`�m0h��Y��X���v��4�Yvb@���h�1�{/^�TM�P�Z̬$$ӌՌ	���R5��?�?Lm N�?ܩl�&_�a|��"}�����ڴr=%A$k�m��(q�:�!U�$�,����(dYC��4��|;.��[t���bzXNn��p�x�V�J�� $=)%���m�l�z��3�����L���[�τ��ѫ��O��xڤ(zHs��_���r�j�o���&@���N�{�l��M�0Zߒˇ�^������E���g���^�d���(���gF4D2��&�k᠘�5��-ϭ��I�~��47F��E49%�>�bK��;�(�E� �r{�	 �_=c��p���S>M�� ���C����`9�)cJ����@�@����~�'UWKW�b�U� �Z:���]��}Ւ��|q���*ͺ�C�e�A#�)y��ȼ���K�|o�B	�(4\���L���+p��*[��@�?�J�]�^���^��b=�5�[���0��йw:gyv2C�����gi�n�w������\~J�0��Q}��d�k���>��6�:lf��P!?l�%N�CY,�k�<	����yZ���x.M��~�<�����L����nF �`9��1M؉��D�:;p%�l��岾�[��g�u�R����tb0�XG\Le��4<&P�߯zʛM���$	y��,��JJ;�%ۯd������6H1�]�u��\��Q{%�*��	��p�&����ܒ�m4��;�^/Q�- ��t�!_P_�E��]����V;������ٗE��糌ec�o	0�d�o\<�k'z�����'(����h(��S���-���FPW�O��4@<Dy�#aq���vu��2B����B���#��_��Ai�J�LS����`Y������|����q(t�ix����[���-�V�&)�t�P�n,}���;-�zo#�'�b����SFz�g����&%���NU� ��Rl���k~IVkE
��YW�HG��	�4�#�"D�ޢ���O��c<jKcaq��>E#��p�v�w=�GNp-�]�E�c�y{������D�G�Q���6��}s��_��%g4>�zʶb3�=��Z�Q:�eO�31}��	��o1G�g�M�E�I�.���x��cl��	�>�D�7�����%C�`��N��f5��L�Vņ���+S�v�_p���r,�{{b�7���ح�!�_�p V� ���UC�j�$���e� tު���Ge���QN������B�2!�*�XqJ#g�п;�Z�TW��5i�I1nv���u3�1B�^�[���b�C}��r�f���}�cNp�ޅ��:Ia�*����F���q<KߨW��Qx��Z� Y��zNa�?9�)��r
�!ν����Q�.����2������3u6�r܁X��Q����W���K�|�J�%s�l׃4q6s>2+��Ą��^����i&G���K�{fͥW)s��?���t@I�9�4����y�㕲|���>��'3E��' ��Z����N�H�v�J P�O�L����LP"�Ult�>��A��B���:ѻ�۴�7��m��0l��ɘK���D~^j��X��D�TE�X�r���UZԺ�W���U,���>��hYȅ^w�-l�=���L(�����9���좋N~�0����*�:��z��JfpyIF�|1-�qF���b��o�|�ģ�خ��ᤲ���x�5lmܜF�M�7\�dBH��;2��4��]��8����_Q��K?��l[S{�'��"�Ğ2��Z)v=��l�p`�O���!*�n7��T�Es�����K�	���a]'+��{*ؕST y�s�6s�P~	#(9��`P�Y�.clĢ[��n�fޠ�R��= 9����� u�݌���s��~f�p
~�S|�i���)B������N"�L�5� [��f�<��痒���Y�`�m	�V�og�������ip��-~cf�(n�^���v�B�O�hO��g6$���D]'�k�S�-���
�W?7%O�{�Br: ���X���:���*ÌkA�Í�ry[2sʽHm�����	�Px��s�~-iv��<��V�E�5���J�=�B����1�	QHL���6}�I �ڍ������Qv�Q�$�t.J�É�KO�W��@졏Q�|�^C�y�`��ߜ�ڐ�Ǔ�01ڝ4����*��6H����U5a���/[�jG�Ȝ�z��������^�pY�~�
�����e~y2�+����J��'�m���y�[S�7S�b&�9�u�����M�2���a�_�`B�g��mwo-���`,�m�~����HPc~ϧ����s`��f�s���GҚڇd�ˀ�|�O/8�eh�
7���n�ʽ2�{>�z��h�F�4'SC����=�"B3L��=(na�<T���w���x�5\���C3��s��aUr�e�{_]�+d�/���֊TX~�c����������Eq��{��O�J$rE>:���A�{c?�<�ނS�P�f,�C��<�2�@�pX�5cյ��.����� ���F�aY@�$�c����/�����=�F~(D砌��Ym��{=�,o���C�h/��o��K�6��������>猋�l����}�9F]�,u?k��ُ�e��c�?�i����Ż�_I���j�m13���6�H�q�{�P'� l�b���U�Ј�.C�6���;�֕!9�b0�2�ӱN�p"/:�翫�/b�+��6���=�
�xW�P�0�\�
%K�������\��5{��^�^��T�Զ�����P�3�|��҃�>4�@����ZЅ����h�$H����I.{G���i,����������$_LӔ�n���k�'m�tfDg>�	{[K�]���	}F"�u�M�8�Cz��u4)�S�� �\EX�m���Io���yt��DtoZ��a���q�kcY����E�~0����ˋ�/��d������؅��~�npv.�<	X�����(���wҶL�7����Y�fslQ�.�tг�k���:��~�x3�@eݸ"$��]K��G��03�0_�;z��sw9�߾6gnL���6c��^�� t+w~��P3�T��#�N�y�ש��YQ�u�P1��4%�by�S�\�l��g�H4�%��Vͫ�I6�7@�Gm1;��l>P Y�ũ����H#>\v���[|N<�܌?�uV�H�mi�l���u9?:R�����Qjn
��hy�YU�L@|T�����(�co6��}7s��mXօ��昐_bE�J��&5$��Ȫ�>}JL	�7���mZ,����F�,�~�"Jw1=+%��q@8TS���O��8��}���7b��c=���O�$ N��ݨl$��v��ٗ��X��
�x���|��H޶R�f貱X�ʇ�,n�3�Ϥ�#�#؜���)�LxƼm��qR�iyj�T<�����S�U4����&�<���KZpq��
��Rr�����< mԥ��^�"��'u����*T�zG��1n��*lj&�
��yv��7-�h"��t����v���]ɨ*�w���j�;�n��?/{��O�#Q%_�Kc��d�QH�	$�^ɟ���-q:��A8��r<u^t�b.��ay�&:�g0��q�<?��y5k�*�Ѕ����l/��b���s+N+Pg���\���8�3���rZ�ɫ�� ����I�B�ۄ:�>
br �
���T�[P��������~P��k��)��Ծ�4�Q�M;���#�JY��Q-ŝ�&�c:�M�YÔ�Zz�b�M�^V׊$�}D�7z��I�U���W��	qԾ�U������j��r�!�1�{'n�<5��#�?���#c��*�.����X`�����&-}ݡyo��r�ɦ��Y�����4���!�Bg!�5�gs���V���KU�&]�$``�p�Y�ő�3���8[�{oAy�!uh��mC�g�n����ۈa8m�G+�j��X�Ź%Z�^4�2�I�厫���;�o[���՗a�5���?��1.�~��H����K�d%4j����XeC����A7��3�<_}G/ȗ^��0Ƽ�b�mH�=�P�H*�Sr��	]��1�� ȥ�� ��x����ŨƦ|)Nz���$	[�漉LoWR�D$Rd�N��VA�w�%���{�@�R�8R�����Qo^x��٘t�x0L��#�Q�C�Y�ml0�Stx1"��|��S�,��ע�kK�����^�cV����Y� rw<���8�&A���F�Z]��uy���N{�M9���sK���E��
���7n|}�	��Lڋ��+c�oF�9l�ȟ�<<y���Б���Ek��
��`�c�1�^���*T�Ҵh��N?��w�6w�⢾��{Q<<�k]�T�;�.6X >��pC��G#d�3�(��|�W��Q��D ܢ�;o�ߗ?�iR|�J*'��׍�k�p�E�����ڜ�uT��T_�lN0���]I���L^�I�wE@���Sn7Ut�j>ET�xJ�vK�8B��<��v*'��E4ǹ^�y��:��E$�&:��J��Mǔ ��N���8`��eO�;��M�o$ZJ&�����D`H��m��7 ����\:�o�vdT��cjי!���Iv�<�W�:OO��p����)F���'`��G@ɥ��8G��K��uw�+��=��^;/�2�տ���l4j�F���$k��rA��ы�tX��Ω���B�"�[d�#�u7cUţ�sW�p��2IK+�;RFg�:�t���Á����6
���l��S�#5�Tl��U�W�$ԩ����D�*#�0��?OzP�F?8��EU�}_�"�,�sh��
�V�'ĳQµ*�r-�?��mZ�l�6j���?����2/Dܱ9ξ\lGA�O�=��b��L�ŧ�nm�h�b�L����V�Sۅ�Q���=[�a�}�Pn���[��~T��u?/�|��M�����#���`����vꓳ����:��i�2�b��m�}#�Ts�Ȯ�)[@ϭ
�VAu�ͺX�z^]n_8b��}�N;����6��3���i�u�y-���I0_�̀����Z�G�/c ����'�z�����ϫ�p�\����~�_A ����b�;zqX�_U�+�!G��-�=7�a`������z�ĕ��v�Q��t8�mX|6��� �G��X{(���~��bcP��� �&	�9M/n�?C.�EТ�?�HT��$-�����؀��������W�L}��
m�0��3+�f�n�����'i�[��#�������7y�T%�q��C95�	�^��L�~�^��,��$
x�� �B_X��(^����̠�����D��we�I2��Rͬ�q��������e	-(��}�8c��;��Aj��I�G��
����C|�P��y5�m'>�x��۾��ʖ��옕k�;\˟���L�~&�m �@��-sqkѩ|�{���i��`>>�'}ͨ�+\ު����q�:����k�]�"��$Y�����2S��0�Y�9�ٶ��]�0��_�-8�ϟ B�� ���3&����x�<�"����J��sf��x�?�^�/�$�B���̿fڵ@���%�h9j�N1�O؅�p�Uo;e��E��*�{��� ��U��$��x#KR�~j��K�m7�j0"����|k.�e|(�~�<�z����'�4S^Ĥ�UL���4�k���4�
N��_XIN�yO���H�
�#���
���I6a��*���b�m�h���R��[i]J`�k�%Ԩ}��ΏP�E݊y|����
��ɴK���tl����o@9�-���h,���]���e��n)�����]�c ɨ���~����8)��X�x +�]_�5Zd�:�K�k�1fg��͞�E��:����7�r3�6U��I!�|��=���N~��x�AωK��-�p!i�.e���a.�7�����0��7�[n߃� ����:B�xҖ�12$�?Ν�`5f�R�T\W}���éÿM]���q�5�+(�y���Rsڛ��yh��bI[�t��%�C+0)�zv�
��Hs��س���������G?�/���cf;����]��� ����B���~q��r�a�3qM�Z�w�<�N6��#���+�I�4�z�)�z�+_������Ғc�]/�������n�1�d����~���9&�A˪����S�*���T�*�p,�[�F�y�0�ͥFm�3_6x�|���â��'Y`���|���2�v���i�~F������GTT�2�w3�#�ެ�k`����$���~?L����*��׀J!�5�a3ƗM��Σ{a�?����\u��$\�]��4r8V���9������<��5t'�#���l;#.��@�@�"C�-	��Nt����jHzxƉ����F%a��, �Q�Z}9�:͑��ѰȠl�sbr�t~��lD�"���:e(��r�X��XP=������gͼ RR^�>��|[�ŕ�-d�~��Z����=��W=�O�.�s����؝�*�י5d��
Q�CX�́l�䗊�pLo3��	.�������{Y�� 
�0Ј\v
h���eW	�O��d�%��^�u��^4�ҥɚR��Z�^�N%m� �e�"� �۷(`��l6��xՎr��U��K�%.�J��˨#�ݔ�&D�\g�U=Q���4��ץ�[�����-9�!��~��F@��+*���z���kȒ�5�Q�*�d��	���R�տ�NGQ=��8��f�ܔZr�_�V̄sS�\�C�`����~M�t%'�� �"sc=���@s먼?�B�D@QW��<57A+ŦUt�x��H����:ZJ���@�/��z��K�7��~b�3u�L��
e�����Ig�H���%L�#��
9�'.9�$�}��Q��^�)�Z�b�*Z����S��'��]&6�/�6'rꗌ=��qY�q��0#ԝ�G"f�NvEҖY��Y��)L�'��r�u,�;�H�*�������E#'��vf���y-��v1���I�"�MU.Cc�I�mP#:��3��qd�@{�e-e� Mٷ�q��R-��O侥������ӥ~�����ܪ+<�x	v�ԥVC��L:t�)Ï�-Z���r6-iȭ����#�2�w<�ӂ9Z�x~�{��fWyϫ���������'���.��g-��Z�q3�<�ZٿgNA`D+(X}�[q��\�`��_�
ૼTJoE�쏎v%A���g�~I��y�7��&�����Vd���(O搎�HNی�����9^�#@������h�_�cZ�Vר�����{{bQ?�F���;�eHA��(pJy�5���fM�xDX]��a�@�R�@�"4�i���Ղ�<����XĬ�qj�k��+��0�I#�޻,�p�7%���T��{ʯ�c?�?MS�>M5��pOs�]�����4]��!��vP�.
��N�pt�V�f&�pEs(�|(��{T�)�E�K3k$o���#(b�V ��n� T����s���&^Ro�ɶh���`x���na	CEC�vҬ����Z;L��|D6I��d��v��p-+-5u�Vw7V+����d 6�lM`A�SSmIZ��G9�n�0� %d�U����ǘ����rKDgg��N-+�K��l��7k�d}k� �_��8�H�R��N�^��j��[��0��"P��8d$-�%"X(%�Y7��]u�T7�k���}�ޭ9�����5�fä�0�e]�C7Gt6fpr�2�Ӎ��Z�{kS��$ܓ��p쬄q)��5~�ܨ!�"�&���'��l?EoC������i���_��.ܽ��0D��1cj��@bVf���j<	���\5�f�oD{f�Qʣ�mD��|�G2���E��U�X�J���A$Eɹj�B�y�V��v�N ,=�?�REA��-a�t�@7P2����\'�{��&/��&�h�mb��?�>h1�Z� ������@rfERb ?�6����"��A}2�<�P���B8�z2vG��v<�Ŏt����+P���X�^����	9�>�k��ӏY�#���G#75���X�5k��"#J=s�G[�aQ�N��$���=���'X>�D�HB����6�^���W��AT	����6+�+޾A$�c�¦��'�V|�������ꀄ���T������YNs�# �zN�K��O��|a��X��H�P�[�S ���(�Kf�!yL�@���78o�q/�Äs�m�R����(>K���v}A���?��<�����UQ�����2#6b7�Z�j:C �ױ`�ꡔZ��AL�(h����[�$��fHp��ܼ��b:w<�ʆ|�8@F�e�b��v��i��v��؂	��^���Lױ"�Ô��~òQ��߷�������(�%���j�1?)���4.g��q�;�b�+E�nToxEz8R�ށ�J#� �lC}�����}��uҞ_q�����*��:�� �Fp��e��QL����Qh);k(���k���aQ�4�CD��Z����Qu΂��ݙ�%�������*��[QkC��W�f��*�$H�ܕ���ǜ�q.��flne+3��~���lΞeDL�`�}�%�{_�ݰ���5I�݈g��H᯷�O�}�K���Ꚗ>�O��K�i5�t^��~�ⰾ��Y����`��bC��-�h;�F�Aѱ������wl�!P�O]%��;�3��l��K/=��A�Uh�bA�½phcn�Y5u*xow'I(���V\V֎��(���D�!�#���_�� 8��etك��	��d�ZPOo	�	��N��qPvc����ym��G�k����AA�>��dR̥�t�O��:9�)8`�{��$:C��Z����:�;�Չ�:�2���>�1̾]#?>��Unj���3u�� t��6����k�H�nC�C���)W����C&�����!�wLQspYV��8��m� �%�<��@��#����|K�1�W�x��GRV6�G��,*e�,_�yi��̲��}y��!���ԩ�5��s��c��(�o���.T}m��T�Z��J��)�qp[��%ߍGC�kf"�)ޝ,�up���YTMT�t5�S���ΐ�hv�_��F�8M%y��s���>�.2(�4�KQ���ߒʑң���"2g�<*��Cf�\f+�����Ĝ+`������ΰ�	C(b����zk��.���ap��ݒ��������àU%W�gh<�A�'��e.�&dW�#nj�̸����<�$��5-X��-�v55����|���`�A�P�#6��]�B������s����H�z�%�\k���k�	D����?�ae�J9��Vo���;��Guh���\M�<�>�$���kٚMVxFo�I�o;�9�5�����(���;�J�,c�7(r�M1b]�/�3��zI��nz<S��ں91ք�q��(g���B�S�u�]��~Z���"Z[����&��pHK�g�j):�Q�Y�3���p� �$N.���L�oZ��J�6�����]+�^��՗d=�yb'c|1������D���1uɪ~l�ڡ)A�HF���y����48������ ~�<:�ȃ��g7����ORVҚ'o�Ԫty�N1I�T��t7 �ۉ�]��2�8e:����v{�|�C���k�=)wS�
NH��E:�5-�3`ԑG7h6�p���k��{�&4����+�]��A�P%:�ިm/���@�4�x�t���JT}��sc�������R¤h��>��R���+C�ZRdU�.�H-�{��,u7����:v�O�[0�� mĿ�\Λ�2���oF���]V���P�E��J�^�#�Z�_��g8B���	k��u�i�Lj��������#R��c����0do(D���63}��O@�&�)���e�Z �[���O|���aE]�~~�'�Z����d���{Ћ7�	'!\�8]�����G�T���/��9�%[u�@�����,����?��5j4׶�-n�L)2�)�K��!�S�?܍Üf ��K�����-�AS��Royc�&��_��8@��K� �0����1ʅ�-SOW�=n�=����r�n9��.���i|`�KR����[��e�6����e/(�1,�l����;?
A��� ��*4��l��Q8f�Y��Cn³+E	�"����M���� ��C��!���� �cX�u<�;ۛ���F	X�)��$���G���l��.ze�i��w"��j�)���2�L�Ine�x9��Db.���&�%����b���M$Y)75i&���l@Va/�����V�P�`��"O��02��Y��r�/��9��Tx�p�<���&m�q����tiآI�I#%���P.O��������R��A�&��sU��L�mN���J���8����=����B�D�c���ɼ��L�|�6���W�E�<S�t�<�`�B�g�|KAa,ղ���!���~\��]
P'�����4�~��%���װ�y���E��<JL�w�)�-B琲������x�;�&
�H��� ��vLQR��/jh(�7��$�k8z��M�w��dկ��)��óxOۮ:O߹���6������[�:�n�[��e�G�޺�b^v��Ϝ�c5��n�g+|Z˛Xqɿ�Xi�]؞/Ȧ��D�p�F��|�D����MC��� FCrӀA �K���,�t೫�1i�rLU
%wu�R����No{偿�9�=G�`C��@�S���Y��QG��f쭓(�Y��#���6p���<h��<8UfbU3Y�oZ�g���Ѷ���HZr��n(�������^��;/χ�������@����?#en(��V
t0�w���kN-����<
�=���7�{���VQz!N�������Õ!2���k/<-RI��=K�����L���Y�.>�F�������b��dS4wa^�����a�h{W]��5� �ݻ��%m���E��X�C���(e��69�6�����ɼ�|$W0�x�6zo͙���#z_���A�����R��@��`��03�4���D�Y.ȼ,���_5p�3�G(�;޿#��;��f�۳\ �����B�0�G����o�p^y��m?¥��Ӆ�&�쁡�<M������v�%z��aϦ]k��L��x�C�$�����U!a��x}��na�6t��qf7H0-͊�$c@Ey��m��!�]$Dc��,ĚJ����S��70��$f��|���*��oƔ	�E刌��LT��7Y�=5��I�H��4�~U!oT8�cC�z��_'��еLf׭�{ɐ4��8%5V1`t�gV�Nsщ2���a=���/�\F�򆌮��ǃ�k?���L�N��)�`�y���#ڻ��������{�l�����f���7��26zy�
��f�]�{��Q��/,'k��1e�H5�����e�/@؋�B��T�_g�����+р�8GR�)fg��O�ኾ�f>��X�ү�����E�w�<�)��4��zs'^��,h˒[o]_fG�J	5%(ߙ�G�]����׎��J�Fw-�:�� tw�MjV�a�E��ޙϏ1��܏O����#)z�ؒr��&���QR�ƭuN�̩t��1HRz��1�X���_��el�o#bZ��A����*�@ӻ�!��� �`|��(մ�H�
�J'pީ�1�k����.ɢN���$L�{N�����h>np���gg�lGW��	���[nc�aMC����v�vv]�*@�w�UUs�I�K+1Q�qj��+{w?�:�?���k]0����G=��b����P�	0}�����?��5X"Ը�K 3�X7�IY��ϓ��܋�J�}�_<\@��oe.�F,�K�nx�e�0za��6�̜s4����9&������H�A;�b�g T8��#jA�q�OU��9|1�h�E8{b�F�[��N�I��"4�K3I�,Q(�� ������ʍrgK|T�F�y����m�A�oc���(5&�`�_�I���B�3�{@�-#?J�t��U,&|[ZR*k����Օm�$��!�~�~��Z��;�N�*l�/�!�1�8�[�pݠY�%������;q{Ŝ� �>�_	6��<��.S�*�m��]�V6���::�P��EE	N���W���q�c���7~r��h#��>=��q0<s2T>kJ&�I��La:ԧT������M�\G�^�a|�њ�2���;r'��������|��wu�}]����+D���Q&��֟�s�9���{2�'^/�8j!S��]uG5ÊRTW`�J�S��ʇ)ɉ��J�`K�8��l�s 572�E٪J�ym_�F��U�i�(=�4
qL�`pVG[3��`]p���NMD�v�n��ƪK�{`��7on�j�L� ���MN�ވ�^���y�����k��a�.:�=!M��t�ƺ���L���2)!ٚ��2�v�fݧ�'m`�C�0�W����j\g�S�@�L��ûH�e� Tt
�u��?@�ڇ��6�{�um#5\�e��p,vQ��u���ȆCI�~���ʨɟ�j�4XMԗ|6�Ի��+A3W�5��S�݆���U'���%Y(�?�9��<Tղ���	_�'��C���Kw>���m�mk�5�����o��CH3��"�X�\�R]S�d�[׏G~���A�e��}�"�>j�3�֓Sҳ4,O���n���چ�lw
F����wx?H� �1�v�p��9I,�JO֚ G��z�)Q���i��$��Y)�h��m�nV Ȗ��$̡�吓��f�}��1�Ə�|p��ϭI����$��e�A���-�k^��OLpN�O�'+���֡��'ŵ�	�Z&/8�X6��
����v!-�S������ݒx@K�"����f�bi���7�T�׆*̿_��7\�+u{�(�����%iZg$���:~��/e"zM����'����HT"qk�h��=��\�:���5����!����0���Q��1A���GZ�&�C��`������ߩ2i���c	z����*L
\i��0���4Q\�Q*����U5�i&�/��2p�X%`̮��@�LAx�!��'�r�.�*�.o6�gJq�'�z����@.�Y@aԂ�%��K.��S�u�G�L�6YBL�E�A��Jg�.�������`���	�;I��H� >�}��X��茸�����L��-�u�S����x!���|<?b�ܵJ'�Qc�� |��t�;�'Ul���m��0.���Y�eV�Ge '��	�.��Q�f�����I,��S�?�Ƴ�R��!�b�[��P^/H��S�e�TS쪜+V��p�u;	�P~�M\�rl?�	sĦj�<Yk\���i�s$c�h�+�3,��dr��	Q~�Q����x���bޠQ��r�F�g���)C^`o"a�ߵ�o�W��z.۱(n�pKun��?��d����<��(�8aRt����뵕�|��m�`��n�'��`�N��'�+����������1�?H�-ڍ�P�L���D�Ew�m6Ah�w��
|��FٜM-4�ߊN�۔a�Z�w��u%*Uy~F�E�`��0U�&���"wQ�T�E��U	���0:������WH��Ŕ�R1LcYP�u�����7r������,J�.����Rwe\�\+ڶu񄠍�(�d���0�X���\�P�N�P�W������6а�_��&b��Wd��2V����7l#�*�-�^�b���+�?����l� ث��!!˵�^WB��a�g�V�P��[���8�"���p�?l��p@ގ$�}O�4�u%�XL�X���䝼�E�4`S!u\hk�v
B���8�x[/��+V�kD/.���/]3}�ď�U�&̤� V}>��NI��O�LkÚ���a�M]"���#�A�b��	 ��I��ȣP��HՎp#��[�dtt������%��������
��Ap8���=Cߵ���}��RȊl��8��&�F��h�6%(o]�!`���`H�jeނbOj&ZQ�Lț��q?#�S�s��� T�F��X.��غ&D�hi��W�JL���>��2�u��y����ۇX��0��y*�ָ&s�=p9�2ܴ:�©�f���|�p8P�8���~3�x��`!�~SS b����*#���\`f�E�{{�"�^�,}�O��u
�,��@6{�` ,�7��^mdl.�Cr
��c���/)��@�N�o��K���u�s����E��������V�>��F�$䝘��kE�R_ ����
!�.�\.�R 3"�B�L+���q�I_M��t ��!�����I���I�^&�S��D=�8{�l>�H�Wb҈�� ����.��������C�ErY��Wi8�7�s��޴�}ܰek�͵�
�]#&���U~aD�'"�ަ��Y��Y��U�s��� A���4C�ah���o�y3�Lֲ�T�:	n�1�t����;���x֒Zh�$�RY�qq��,�[���@�ħB��$�F�~<��OWICL�uJ��-����3̳�u��9���}�z�Y�p��V�D����[��%�����4�V4/�X�.ݽ7�͟!:q�f�T�Y�$�uD��/��`���V�՜��]��'�o;�y<ƣ�T�Ʃ����K��$Mܖ��g �?|�gb��ҽ�|_��d����-�?���m%�f���zY�E�d�c����2���C��oCk��4Zr��]`��79��:�;ǈ��H�m�E�DG��{ߠ��W�6B<M`)*�PQ�ѱ ���0�,�����V %�����[�S�!�)c��ʩr}4�K7��B�ue��$G�xS¹��	c�Q^�	kǃ��)&�(y�6��l�4�nv��ŧ�Ň�[�D�a��R��̆��t�M8�����(�����z��BU�9�R]m�ٗ�R���d	Gm��m$d��D�!j����#
�ĠSoj��׉���|�����;��
��nl�?L��zehA��C�)��a��=�g�]����Em��#�Q��I�4�?�6]K	�eZ��Q� ]�;�0AM�WN9b���DE��S��@���"��{���&=0ۘń2�ߚ�˛V�W�s�q��m�z�VYQo�绅;� ���eM3?��V�l}���\���������	�Q滇���]�P��1�=_O,xqY�3=")�v5p%q�?�/�����M?G�,c��G��	��A�FƦ0U~�I5�K3oJ!tt�2 pr	��el-̞�g����r|>��}��؂�Z���Oc,��6�>ʋ�Мt:�pA�˂l;�`%�Z�ߎd�N4�p�
�\���� ��c������b��
 h�E��^�E��ŀ�iҙw�#A���6�K���e��/�����i���a ��3M/�q"Hh��&|u��o
��a/?���=�!�H��<�U�MN�w��8Gg�<��Rp�[��[�4?�p�!YT��d��d7���hRHVo��bQ�*,����F=�R��׀L4K!sPpiq�U1�I���N�Qx�!; �w]#hN�^q%��i1Yh�YoO`O�9}����5 ��'n�e:�q�{�[2A��f�4_G>~�/G�gRPnF����,�>�/��@�+���2*];p]�̮������ ���놅�ݺdx$3^���C��:�Q98�X���wk~��:�ϧ�����KJ1kR�lޑ��\"JG΄
�SR�o��]j����	.��-a�;�؍dl8��0w7K��B$�Rm֌8Ła�U����BG>��o��~+}�N,�8��%�Q�R1��U��b�~�� ���t7�I�f�ع� ���l���2��k�2
b����Y�&�
^�k�HW�����Y��g	@�� ��T�`E1��.G* !'���`u9:[rHdœ|^9���]2����$s6[�u���)�#3�I�[6�kD�M鿋�,��m�c	�0��G��c���9Z��:�M\���KZEy���^�w�]$�`t@{�A�Ӗ�����8
�">6��DT�3��\~9>��M��^:ƌ��|����~�\����*��Ѹ�@���7%�R���ȿ��$㈏��؜�L8�RW�
��Dc"�`�k1�O����B����f���/�ɗI�p����{k�n�ޢp�� �M���V��ɋr7�G�M�j%�H�b�J%�^��r�W�o��*�@V1��j��D�Dd��F]j��m�����p]QS������c[��)G�]�MqUW�hPg�n9�/7>֝	���gs.�Fte��ŪO�x�2/��='m�q��*�+@!�N��NA��9���"&��c3��'hn%����q�nf�gF�������h5P�
L��������nph4C+]�î
�H�i�vb����G���9���z)�N������-�h̷T��R`�@��?��gL^mr�ͣMi��+O�
�	���j��#=�TK�����+Nn~J�H�m�K���g9ߪ<(���`x�I���g�+�T��b�T�Ǣq!L�zr�� ��tC˅-k���U��)Bz����*�<�tR���+Sjt�0�d�Zp�Q�>[f�w��WA����[3{AG�^�6�%$�w�X+!q�@�g>K��;I	i��?�G�ui�pӿo��f*�Ɍ���ʺ^#()^�r�[E��Ǉz|�+~C\�L�ܼ��w����w��a���&���$�!��F���*�]��d/u�����e�QL��\�o��°���N�>�;���0K���ϳGՠ���մ��'�(��?�����q��X���Xc�����@���7��H"&[{G'��2�>��a��	�fWS���E�އ�Q��6*2;S�X��W�X7� �:�W�p˿ ������p���A�ļ�]߾8��/<������d-�,�*�����`)�P\T�Gu�̎�{G�Z�	��)��R O���'�3�+k!�nL�N�$/;��駏��	�=
�EW�W�V��)85��:�<�~���&����]`�@$5:�F�y�7�
)�e+��=G \
X���X|�A<�XLKɠ��4֪��B߲��<쇠̫�n���J�`�����^\�.J��}���U�!
O��|߾I&��v�;��p��1'Kb2+��� p%�]�~�t���(w��1���V\8�G�3�&`�#dm��[�;�MQWh%��l�1�@����,�xѻ"�w⛚ ��x6� *e���GD��-X��x�%#f8躟���{�Nn^� C��`�?dM5���	xT�`{0/*���#|�Q����iNj�p��k����>3��Q�h�Re=���7��@]|,J�������&�p�ê��5��S5r��X}��*�e�uf�^���WA� �Cs@T��ɷ����#s����*�j���(:�}�-6�ݖ`�V�t�a�5��Ve�)�Qj�uT�Pp�1U��L��v��WC��T'p��t{�2��)�?9_u��ʮ95��"�+�槳���c�!v�L�;��� ���s�ߤ�&��5���5�����>�d�,�s�D��IGq��D��MX���	�
S���}����gм7����M;8r��C`�{�*�&�2�;�c��'[�	֧U�]P��s�=�>��F��s"\'7jz78����1&����t&"Ҋ[7_��o�Rl+�r��j�Bǜ��y��v)_B7d����� ��"��X#.26v4��j#9I���Z(����]x�x� �?����X��:�n
^ʩ���$����>h�F;��OQQǀ�?u:b6�<!����U��'İ�$��@nC4o��RRz�T���Lp��*��X�e8�q�C����f�pN=} �����./�U�0�.rv-/���}S�ק>Ţ'ag�ڜL�QGt�����o��������:��H3gw� jp`�XB�������=N�Z)"p�u�h#ta������ڮ�n/�$T�FHv��[����q���?~�~	s���|�C�68��s�`�ȭ.s߫O"6�9 �ȱ K�@��2�JQ���Ĕ��U�z�CT���E0hpJ���I�BH~ ���9^T+�l6�#R8��1.��>#0W,�~�T+�#ȭ4�a��=�h{�]�d�i���������sAu[[X7lG��Ep�ĂX���3!�h��ɪ9(?�q��ҵv�1ПF�F�e�Fӗ�#�;b�7ƹtg�!�t���%�Q�Z/�N�6�$A�Q��Q�}�7L)_��i��$���8�p�#�面;������!�:3eף�%��I4R��yz�5�eRk��%k�Mͮ2���5�{'?��@�&f�H$�5?���c��T��� R� v�ʕ�����;l�rJ�*x�P���u]�K�e����(�"8�c�!=3A��n���J⋲��~:�OoڄaW��~!À���7_��d�v��� ]�m�P֕3�g(Nk�<���/��0r��<Q������u����hU�h�����(o�rN:���j���Wj/�h#M\���^U��Yb��(�La�zsi���l����;AL��؜)5�]��
%1,�F���Qp��і�S�ۓ�9ζ�YThDR���'{M�n.eA��éQ���ĥₐ��,�Ԛ����9lf�1�z�O��(�!2?�x�Y�[��7v*��@K��5%��⟥��(�L{>�8��O���m�L����	D7sW�����؁n\�V#���e�[��O�2�~A-UH�B��#�����(X������֕w�W���aN	5����xx�����ޯɎ�G�M)�K�qm�g�l
�V�d*k��{�i���/)'�v=,Y�$_�΂�DR%��Sm��v��V�?��r��,j��?�b��7I$J��)�Q�Lv�3��G���`v���	�w�Z9��c����PX�8&�ᣏ
��/�
�#��|"*�܉���=~�?LN疇��i%�������B �a��-nq������.n��_D����sr{�*�n`a%���ǮW���9g$OZ��PZ8�����}1P�	�5�B���_:E�t�����/���CD^:�%��J�=k+5���Q9���U~�M2�����d�7��}��oW�O,��2G��U8���x��x���x�N�a�Q0��,�����c��~��<{|����c�!'�Z
}��x�����Y��I=������L�߄eX����ˡ�*�BH�I��r�m�=y��gռ��xB�*�pX�;Ǥl��_�]��P�/�9���t�g�cd~��ُ����<���"����5�>+ߎ�<ac'��P�b^��a|~�%�g���%���/��>�J�N�b� ��گv.�>ҡb=��e���N<�Lw��I'`���C ?�[����i8B�Z�o��l`w��m��;$Ih���>lZ)�l�M���.����ǉ�I�� �	u��$���&�Q!��������:)�c���$�����o����O��&`a�#�����*��(�!��F�xm��x���^�ņx�T)����\U��n��;kB�vZf;�SL(pH�]�|��� ��]�u�q��e���.��UL�Iwc������(��p@�^��M�>�61ѩ����>n��3���;P��PQ�������,���b�l�J2S������g��R�����H�u��N�kL2�rt��7��"���c� �����:���z����-�˝uΗ�h���[[3#��K�l���5	�NB��m�n0z����{����c0��,��"zx_��o��2��@����}�.���um
�n������������_p&��I���mm�Ǯl1h,ת¿�J�V�����+ZZ�rw����FA��l��S���|X��D��	�҃;_A��B��G��?�Uʈ_,bY�8KW�V7���!?׀���\��v�X|�u�������;`�ui���f����fos���'�f���پ'���H�X��j�ь��{_�����4���Y�21j����A��d|�~����>+_�7����A�2C�t��#?:�����l�-�Q��l>O��'��B���k�� 8�������C�@��E�j�;�x�/��"W�"�6�k�%j��z���~����jt0<��P!�̐����x����C�?˨��ED�몘�v��0�OZ�O�k:���{���u�2�s2��l�D^�Sʏ�2���0k�k�JA�$(;4�A
���E�1\�/P�n�L+�6gB����;�,�����|�n8��j�U�ڂ�70�_��o�5�f��&:�.0t�A��S�<�S��* �Y�<JeӀH\�#5})t���8H�
wM����%�
�QC�z�Yd�ޢś"��8�O� �鳏M+�)8����)�j;D�I��/�i�ϝ$�r��6迡��P�w<m.�J�0��7��ks�	��-d��u����}�h�_�O����q�ہ��$S.[!6���U�Cn�v��i�ޅb��ߝ�PU|�z.~��%Hc��`Kz������KY�#[�N�3;�g�ͮ�p1��E�]Ȁ�^���%���´zqMgQ�4�'T�\Et&k��Ya�(cU(��Y ��=J��U1��J/��[����G�r��_z��|�v�.!0w��R�DJ �x�>=g��>|Qަ	zih�M`�k,��:%��X?�Ro���CՓys0�_o�W���܀�Y��?��js�����P���%�DK�'ª��'�Ը�#y�)��E�qX�6'�A� Qm�������j�.t,,�њ�?��H�����y����YSY�C���Jd��t��(Ķ�����ܸ�4~v?���[G�{�����ˈ�B�g�I���j�����\G}��sf��vl)�0z��8�=��֚Z���E��K��8F!�sx�x'l��*����&
��zVuP���`��SdB��#h���́�o,,X;Kg0ܻ�A: C�g���'��.���CP�&H�tЍ�~���s�Q�+������7�����R��v2�q_�	�\]q5���C����;1g�~P#���Z�5��NR�;gn�ə�s���4��Xы���2T<�$dd�m9%���}Q�2���<['��F���޳��ɓ�Tg��}�86�5�_I\�����#t%g?!B;��d�	7e�|(�*�`���?�b�]���9��-��6W�k�0����%;�8���ʑ�=+zy�n%2�{o���f��V��*�<�O(��r}si�i�a�؅�X�B�B���� [/��߁�J���kE����@��?��+�W4#�Zq�2Rda3Y���Ąr�De�L�c���K��y�7��'�G3�s��e1\��c��p�Y-*b#Y2��y��M�ZAOc��TW�jN��1��f?7 !�9�h�"�T�K�Ő��9�?H8Y��k����6���Xj��|����M?ꗤ��^�m��}�X��'�sf��m��!i�-֍`ݮ�� *����@�2�Z���d����'8�:9lGʿe�ӑ�@R�W�z7�t"�K�4y+��nuB�CP�#�ľ�A����������j+2�@��Kq�S>�A9��b��O�dG�K��+���6�!��5f*s2���4��l��I �N��-, �O}���G�{�M,N� �O臗�9'$4K��&��G��l�?�j~��vx��ٵ-#[�����������*��$��n5��CR��麘�]WQfEQ/����±,f��o��F��OЫ�-�`{$�(4�n��&e͡�.����Ue� ?3����
�_0!�:k������XH��yqz�' �{Nq���ru���HZ6�C<��E��K�?��]�MbPO�!�Q*wh�|��bd[\Y%��d�c������ ����n�$I�U=�������$# ��^r&0����E�*�7X��?F���pc,d»�n�z�W��L�K�mt?�O� �����H$r��hܳ���lQ������ma]�"�Nq%c��ywj���Ş�`��ػ�G�i�!F�?�A��y[�Rl�����^*�:)1� t��ݡ�-�{�!{������������� ��5�~Jk:�;�J�x�����"�7�K�Bz��v��+��%jɈ�I�}��@�;f���#�#�Eg�w=�b(���~Uf��IT��g�ޝm�s1�����k3��`v
����h�n�f&�"�
��X�J��u)�/#�ͼ�z���D�MqRn?���:Z���"��X��;�1㒑WG�XA�2%:�q/ ;��\���>��z�$��]�kJlk+4�m��h �2�Ӛ͌�âي���jX��kT`^�7���t5�F<D��Bh��5>�'e���M ���lNG/� ����~f��)T3HώkG���9�m��oB"}��9�Ҷ���A?�N�a�lb��`�~Q4�?7'�O�R}m|r9���S��Z�����D��9�LcM�`�Z HIgf,��2�80P�R�v��)Kd���O�6b.P��I+JO<(�t��q��eu��A��)&C�o_�Ø��r�!�%��$v��X�厇*hV0ͅO�>6I��A�>*��@�H6,ݎf�9����r��^�]JC��qd�%F�p��b����a>"/%��+�5�%�oS��O_�w�5���&�Q&"��>C4Ti~����F=
и]Ț���}�f�f�2Uu�����=�sl2�R�2TP|�B\w�(m�#u�n�0K�;��o<�2	v|:3���P�6�	 /���k��@Zl8�?����3܃v��U�/�ɝ�YJQ���܅N�����}kTs{�w�������g5�=����u�2�*�y��7�>'��U'�s��7(ù��g�9�ض�i�>���dhc@-2���T�����3QC�_N��x6��s�8��G'9@�A4�&SXs���`DDߊe��\&״���Y\]t����JZ�7��%�%��d�tf�jC����wGJ�]ろA�u���tH����_�f��'W���cEi9FH!1�%�|u��z"��.p�I��f"����F��C� 0��$��J��*�*�')k G�(��\_ �ܩ�m�����uF�U/��הe2���8�t�J���M����`�""�R߬����x���'�UAh�X�S�񗰳�"�qH-Ҝȸ	@�W�UD?xy�[�,�+�X����d�Z�"�A��缁�?�(}��!�Ga1��y>k��&���u�L�r
T�Co;�A97��S�NUk[>�٬!KU��+<��V~������=e���g,eib����5+j�O��
r	�I��W��q�31��"&�Bމ����W�,;��g	%�8q�,�&�p	Կ<ܸ�g�×g���w8C���=��k~Z���^N-�iܨ8�6�*�S�Oy�_
	Ng�q�˭JVh޸O�b(��6I
�mw�H/��Uq���u����&|���������T�Q��^�9��S{a���S]>g�)��L�%P����ޕ���߮��.�������3Ν�1+M{�T�������sba��IH}�ﾞ<FІp1��O��C�}+�g�$�TO���p��Z.��3WwᲺl
�y���YB@8�(�Q��20��E�:^�'�S̀&г
��k�W��+���7-��, e|��@f�2��otsA�	�ʹ��f�ӏ�öw��6,	��w���0��A���V�mi�d�HsJE��G�F��ԛyG��G�K��Ϭfϒ< �c�uNQ� c	rm�u���.9�u/��Ɖc���l����sU0o	g���Ič���ܹ��Φ���O�3����\H9��ƌ�=���|��k��+��S�Ys	�|���]�f�䥎�Q�.̄]�Q;��ho|�6�y�}"��Ծ����P��"��/^����s�U��@�ĸ	>��6��J	�w�of�x[��]@S���m�Q�Gq��2,_�
#�i�:|;�-;��ڱ�.RtFZ�0gCj�p�xrܣVn	�!̷D�����S�P3U�;N��H���`G��XE2Y��$�1x��Gb� ��<݌�}/eV	mG���W)D�eq��~�!�
'7�u�⦿��Ѿ��|��[fQ���೔�[��ҩ����^�I��Bl��̅�K�:a^e��$���+��
�"h�@.�h�
�,vߌb���-��O�\����j[�ǯ?ų\J�}n��?�ݤ�)>�d*�_x9��%�#J�4�ݔ2���[פ�����v�+6Q�4�>NL�����+�����%a��uwWgK��@��a��I�u�p���<MC�����5�P�wa"��;n��'K1�F@�jg�|�9�Yp�#7`�*�p�E$��O��X4�G�1��Ai`�;���[l���pir��b�SƉ��w5�yS��r��	22�@�8?e�BM��I�c�}�!a\�!��Z���^�D(�!�1��L"A��DC6�,���s��<�a�Pֵ �_��Q����,��p�J6� n��	_�ޑ/n,����K,X����#�^D��1�%E�ٓ���U�\��&	�s9�C^���6���$�~?=J�uJd�(�!(+i3@X�BP%��h����-#cj|y{��(/�'��9�c����l�K!� *�y4�g6�5Kh	.�q�0h�*֘�9bf������Q^�Y�f�j@��������t�r��͆w:�&�2�I4�!����yޯ���{�y��a��y�Y���J�4f�u���V���@k�`�����t�)��j�NT{���Xa�dxX=1�20���
%�e_I@��P�kqΕ
?$�Est](v�':i��J�-,ۙ����T��:�q�����zB]o�;��Sȉ����&��\�y�C
L)���4�-����������x��s@��d��ƎI����eiXO�:!�.$4��n�esL���q9!��������à��0
f��P0��{�{u)烰X��/��y�z�^\]�.N�_rB#[�"�� �mO�w}M �KI
�դ�cT���{Խ����^�]��`x�[L�������:��,!&�br�#gC�&P��l����y4����C�=Ҷ���ӈr��N��p��?�W>[�-�K�˞�=�>�P����M'i9VL���E��4j�_`Z�T��`���>�N�jF�>Mi����_�h1���٥]o�<UfE�w���w�����\P�����`��_�#�`�vw��z=i	>�����d]33��rA�jKT����c/E�Ct�}�(w�������(�=}����C5L[��R�}q.�C�	0�U5��:����ا�a|:n�6�MScq>��{ڒpښ��n_�;�X��3��:�c��߀�a�CY�i��ʡ�s�҈�0��8i:���y\��M�\{���T����bF{q��O�Z��	�j��4N�|��8��+.�͑�Q���<��+�pd�ʩ���w��SU��0���'�쎲�/[_ƌ�.�zT@����Cl�������֓�Y�5. (9ruq���=��,r�e���l�4:Y��E�q�Җ��F��"�0|�ĸ ~�ꖐS2�y��v�f&�������A���d�|I�@}�=kC
LW�\&�Ԍ�U��q46��(��Q}�_�����+�g�F�tj�A���i��O�-'h+�r4�B��X��k0]����-r/�!���g��4�{���O}VVl8�
檂
�&��:��;�
Y[]��Z+��H+�-l�HY�����l6�I���$��t,:�GM�qл[&�p�Dю������h���؝]+qtQ����ͩ!O`��!��鎯�A|�i�/�d�qGycU��x=�pӾ`���:.��4/��{�_R
��U��S�ou�b��oHԨW��r�cU==�"��{��n6�-��㨿22��W�ش��@��1Y���f��j�,m�C[0��v�Y]��5�'�-I�kh�.�݆-柭�䢳6R�s\�J�br�*��Y��l{�`�0Ko�pw(T,-܌E�������X�[���Q��J�5߻��=�M�z��YX7�g)�S�4;I�9W-C�Z).J�.�~��ruHx���hP��Gݓ����I����N����Pӗ����;�зݒ����z;���Nx����V`�n&�#,���@�����Q�dOcgފ�-��:���%�l��6\�93��o�S�ՠsp�%7�o������*G�2�w��(�%4�Hp���8��Gw��Dnjm�Ob��YW���4��^�U�+�)�^�.��B����Ô���C�ZR�2��D���[Pi��-Я'U㏛	� ��P�����~	��=��� h��V���!AN���"Z�*�J��2�v�I���T�;џ# �+'m?�«�����.�ᇖ9��3���[��4��r�.�4����a��d�$����Al��7� �Ⱥ�g�i=6�=$c����@ҽ���7�Y��-$4Wvl�nF�G�3��$�� _����Ȟ�6Q�׬i|��c�Z���'Vy2/���,Lc�߹��3Ai:g埶[2�@}��o�ef�F��3S�˶�"a~B�� X��f~xՔw,�*����)u��e��~H}>�A��]y�\��F�#���2y���Q�W��L�"��ג��h��=�;8�p���M?��(έU��"��m���`��f��n����>��O��������XGsF\����/f�ZF��z�Q8A���Zh{�8ֻu���h i�f�L��U�8J�L���,����d�|}^������Xm�=��3���3i=kL$�e��dx�L�v��Ⱦ/��d���pd?|�Hw���W��`��T�wl��=��p+�
�����W�g-$�l�`��=��qXf����Ҋ<3h��I-�� {�2�sW<�@�0׀�Ő۲�5
�B/��c8�����Ź=�V�L�"KdQ�]k�Y��h����le��˶Bt�Ek2�E�?3M�Q}��u�SɯE�/t�܅C"쟌���X>�P�$Ւ�T&xms����o�`�kvW{g�Y� �oȴ�yA&���CZ, �dO�+&� N-�4�8��κ������-o?���Gd�2P'���e^�����{��8O�H��ER4�ؤF19��"��޼� @�d��p�-^�ǰ�p[�l6��)yްh������Nǃ+�kK���j�Ԧ��QH-K��1�}�V(	뫪���V ������k4�\5�"�jX�z�ջwa��Y4�h (B���iN�p��R$֮�G��k�.��B�Ð�m��e�}t�J	���4��钯OB+j��{o����\�`$�nȡ[�I�}jlF5����tm B��r|��h���5��j k���)�,W'i��	o��P�n�o�TK"zTOr��3S�_ŝ[_!����f2�7{q_�*����x��;��2��h� ��6�=�+BI����h�c&�s���~+>��C�|�dR,uG�Y�t,�>�(�Ģ�ZQ�s����q���Nf�q����/d[���heݦ�/���/-RXe-+��[���^��כs�& �a��z�p8���u-��?�F-�ă�4� �H9x^���T?��]wT�{�B%22p�8��i�W�Q�	�m�1���:�F���`�A�L�Y!'4`�A ��OP��xw�Eb��t����O��i^���kP`��Gw���x�y���R�/���zu������da�� �(
u�8֎7ލY%ʝdS�
�ܦX��}`	A�RB��N>�5�`�:JdT��m!#T����ZM��9A�?$_����� ^�1,��,	e�o��:ו����IĿמ��^�W�����O��k��#��M;��>,�+�d���/3:�K))�|I�&��`��*�W�$���1�mY�^x�\�iR�����y���`q%�v�`	�1�_U�����>�ѼX<������-H}������p�l_5c�%P���3!���R��QF���a�}P�Kv$3骰�7$��c(�T5;lSn�D���&�+��7�Nt�%S�&H>�5�o��Ӆ}���<�7H&	iI�"��U�~(9`gz����é�3�	��0M�F�t���{��,ad�����\K
zG�#~���9F;ͮ9xζ
o����a	� ��
��7-f����^�Q�I��O����.z�4E�(�)	c?��%D�ԗ'49�%�����,"����.���HL���3-͟m1}X����2q[���xx��J�\[l"P������n���� ��g��%�f�O"��FY~Tɖ�=���� �؎%Z����ާ��%�O\�E ��B3��6,l��m�<:ڌ�qO��Ƕ^�!�Fwk�Q纕DM��`���e�mEN�@�<�9���[�;��	!����� N 9�'��6
(���SuI�BHϺ>chQ��mn|�z"�����ek�����'A���.qW#X�Yy筴���!�_�q����7W`,cZA��zc�s���a��cO���gY�U��������h.lAU�lx\Q��k�r�����DD�~�x�u@q �l�Q���B��>d#�ӫ��K�bߚWr��d\�?�h_�.��!KJ����̐������ ��5�P�2���g7C��7wh�p���R�b-VR�,����<�.�G���'_1դ�ף���Yk��������|n�N�^�'^��
�o��r��9��J�^v�[���y!~���lڗ� �j+9�
��큳q)Ï ���<����	n�5.�z���	�m��*5믾TJ�[�!	��Zp�B�c��K ��ua��J���?G4r��FBeܽ��ui �G�gO|���;~ǖv] v��Y�/�$�͝��_õW�'"β��-6h�nب���Na�;5�f�:ZQ&r���k���:�=�pk���I�a���l��z�=�p�_�q^�ٷf�0��V_��N��s|hi5�d҇ڐ�]:t�h���= ����^jio�ElG�P�g�Ć�"��9���`����S��J&]Y;�7�H��j�w�܋[a�10��"(y]�O?��_z�{o� ~6T�ח#�a��C�{��Qz��}a�������y\a
�0E`x�Ub1�>��ھŎJ�%�Hń�jA�ɰ6=�{J_#O]�Y�-90�-��:&����U)�����l�ov�b����r7G��'�E2���<_@�#�X�&�+M�w��4@��ǑY�p�p��6����U�?h��X�V��
꿐�I�C�nC0�JY��E	�U�� ��:=�8��9	y�њF��^M���>>��>g�9fNXk�����HV�߉��@�p(:`����y�0Q�� �܀R+F�S�mv�?�Ҟ��/aC9��U C�$A��qj+`�����!r�C���H�Nl�r�/
}�X�B>^����
+b�X^8[���c	�a���r�7�h�k�������#�:r���u�"]��+����[�lA'ȟf�)*�B�ë� �\��S@ }+fRC(�:�F	��~�$��S��)���)���j�ʹ����¹��Q��I�E�$�	�;��|��pW���YO�$�&Z:���G���1F>:pɺ��O�m"���� ��ۃȝ9�l	����GoŹ�F�ۡ�c�uN�.۰��z����2_C�c��)p������:���)�����v>��%R����aP�.|��?A����y�Oڛ�Pe2V�
��7�g)��pb�ww�4="�0
�;)����1����ն��p��u;7/��s�QI���'1�� W�� P��WOڼm�HZ1f�-�F~�4f2�������U�i�XmkL5TP�uZؔJAi�pm��ج~O�bo��RD02�hN昐��A�!8D�rX���c��)��HL�)�ծfHl�h�� �5#�E�����$�B.��aIxa.�=�Yi�񘪩]2��X�#�>�3�*cyo�Z�j$��Tp氈k%�z�nÙ�v	��	�_����}f�Tp�F�@)#
�~�j(k�B���ޚ{y/��m&2�OYf��(`��b\����k�=�zn�k��VEݣ'7�.a�T�3�YahC>2)>\������.p���\���Y�D� E��mQ+�@o8m���ʼ=�8WZW�����Y�_FwiB�=h�j�1����s?�����A��?5~a3�|�u������-�A�s�MP?1�{����ܪ����y*��h��?k����:�6��
�a�*T�ڧ�J��˺yYWp�_0�X|�L��d0{�Da��q78X�|�θ����6��c��@�D���� 51j6������?�q�SC����FS?����Q4fF��LC	�����EvZP>4ʌX��i��[ęL,?��zCdx�Q8jRs�x���2?K�����uBS��_`������s$bI�×�t�挵��BEU7Ӏ�J�Kڗֳ��&��u,T㉏��yq,}凿Ecr�k'1KY� t�{�=�![j��Żl�e�[�t`�L ��`�輦dZ%߉�:>Qq7E��\_8a ��-J�'{��f&��h��5����3�f��t��-��B�&c���SNY��q�#i���mS":�_�ɼ�W�O�/Ry����f��t��˻���S��j�aktJ��u?l?(7̴��c�����GsC!
�5&DH'�p�i��fi���㋨��6��B�&���6۳��-`2b\Z��a��>qA�4#}�d�&{��H�?�l�Z�Z��}�yb�2/��������q�@��#�f�-v�$#�6>��@�Fj�z]�v*�ĺ�$ؼ�! �wn�Dq���V��څn�Ù�^�H��U��;.85(�fḐw�#jԮt��?�����ta�ڕ�s~J�6���c}մna2ZK�  
r���U>�gg�C9@A�[&�a��!}|7��ke���b��׮4�÷T�f :RߑR�u*Cg|3v�������$��Tl2�$=��MX>7)%��^e�޼&��ת�^\��g0��tƮ׀��_�z_�.���3\�
��%��Rm�]�h�I�-G"�'�KD5YVn�j�c�٩���:� vUQ�w�ОH����,�����3������NX�՛�_�?Sh�p�P����TV�"p{�:-�`G���mQ�����=�`ܟ7V+�R���燔j^T�j��Y7T����\x8
�Uf�J��}K\Z����\O��GK��fC�\;���u�4B�h)�[mN�m��8�`.�w��bHX֨Q��i���re� r͉�����1��ژ}0��E�j�g�jj"��($��܏�}pƆ/��h	�X�jz�oT�a��-<��m%� �~R��$am���z\��~�	�u���R�6�����,�}�|ڒ�v��/�x�j�Q�G#�V�?�u+lp�Ks�E\GOrx��R�U8��ޔ�W��+�Z#_�=T�-v�n(}��h���O�[����l�T�7�8�j���蚹/ز��P�� GHe$���dEW���4�Gw�(RR׳�B����˄���ק�v�  ��1�t�0��7He�6E�	!���,�������jf;9��PF̕p�"w	�`��?���£���Tѣ�e5tı=���u��>�~��oMR+�����%�."�%���N�&��98 ��ȅu�����p�Hz���f���+�����z�l`"3�LG�%��$�M�R�|4���:@`���.�j�!���ƜG�;��C�k)N�x�!w �F�%���z4�W_K-�j��|C0\�45�إ���!�����f�JN7��1����ҏD궅XY������r."�B78����|X�#��gaL�=3��q�� ����db�1�(C*S�9Π01[��p&�"l�͛	��x}���t~C�]8|4���u��V��
q�O���`0�F2;��s$A�K2��tl�#�<|�T��y�*lEp�^	�����F��B�p�pH�`��ȓK��K5�t4�$��f�_��^	?S��H�@�{�M#i�M��w�T�!i�G<c��1ˉ�ԊJ�Xu��$�&Oiwח�J[�E�)[ʱ��%es��lW�P8��Ht��L��� N�eӿu�9-Et�^({B��i��qV�G��IX��W5����C�Xpk��C�V�Y�d�wEy���qJI>V������6�y>�1�
�U��M�	��02�`��m���Qa�AlA�Z�C	���N����|,�DП9���	���\L�^�O�م8�XV��\۔��E��8�o�e?�����[вw�� �	[��^e�kW87��jR��C�'�Э���c�J�0�/m����'0M>!?�2�B/0��e��<ڍCTQ0_��>�a�*#s����@� h��� �Io�p�`�,N�7����^�@�ry�WP&X*A7�Z���:i;'�M�<-��Gu���!q�!��K[X�fAV^����F��F������Q'3�ʹ~�DN�f^��z��תS@����m+��`��{w���يIq�_�Ul.S���cPp�#�z�r��]���c��ݷ�*���^�c�ﳔ�G*�e�����?��J#�]��\�i�rc�S�C��N`CP�s;�+V�mʟJ�N�砋�ȏ'�U@�D���Ne��n�>�^��4�W��".���c�iU��n����Nb�R����Bx3?��W��ԣ,�֊!~]TA��S:+�oS���H��mw��w�<�����z�g0�r7�B��8x|U�%on~�8mA��	.�	��Bi��� 00��N�s�n�|<�X�.��w��Z��O�ѩ=���YV�L���zm��Z�LK&G~7tf��R������\Մ����Ğ���\諢�w^j���;K��B��C�i�.�d+傍�O�-^
v�ME�s��J�E_,�B;���������$�=��a���� k�fb��εO�e�����&=�4Z�?�:�54�q���48��)W�B���=�wN�O;0���L����ϼ�M����C��@U:�C+-s��$Ql5��(�#R��z���H�n�i�(�3}8�-�j�c��rL��?(��"��߁9�w��_|r�1��zC�/W��Dp�z�"x,�����$9za��K���r�g����d������dl{z*��������Q6�����;
%ܒ@uU�y��|Sҕb��Z���"\Y�,�I���X�de�=���n�����thUw;�w ��+Hs�T/)����G"̧>Ix3a�cPE͕!�n�[ B�u���F�:�I���V�UQq~�.��*�t��;�F��q
��$��[K�$�%��M6"�?��;���Y�7q�ĉp���n���U�i����h�.�ʸ��!k��[x��w{S�~���J�6��,K�pv��o�r��^t�N��`�|���p����A'�D�ӣ>R��]S��^+CiPf��;vIJ,����t�$~�"��;�Z>�YKF���F�/?RB~�~a��?�{�^,���	RC�y9)�}�|S�b��e�U9	�]�Z�~�d҉t�m�����A�����bL��o�˱q3���Ɠx�L��a��� k����M&��^��@U����Ga�g���I�O��m�d��wL*h�=gؿ����N��_M�c5���hñ[�ռ�'��W����E���W�r�†xAi��5�K֎ծk����t�@J�9KNH�Q�w��,�.�0"C��3u�X7�,��fM��=K5���F/����EZ����tm��ﺚ�B�)]��XW/�)�SpRb>6�F��i..�uMX� ��^�'x���;[�Q�9x�%^t�D>����Q�2/�]ml)s�TЯ��r�'��C���rr�^k��Z K���MJ��q�h�Z>冯sf����)���} W�� �&"�L��]�^eB������44:���#4���I��hy�B]+��7�S~0��Ҟ����м}E��K��6E Piz)Y333�[��4 y��A�Ds�,�����g"�O/�(��x��y�xU�-���۫~�<Ynp�_FH �ȸI�{b��ÿ�=}|�R1~�K-����������)8���X �����	O˻z�A!Cu.�4�ǯ�E�7��-.,Ԥ4�tp�0A�@�L�
E\�w��p[��N�J5��r*�g�/rӔbkj�Z�ց���㠫ey�n6��<M�@� �SDLH�o��x����N'����{b��ϱ�!u�Hn���Ӝ����'{<��DQ�J�9o+
t���|چ��y���Gt=O�4_Ѡ;��^\i�h��{�g�l�7O��<���>��%_ ��##Q��?�^�&y=�^�4-,���(��]Br�Y��e��#�m0�{������.��}ݷ�pq�q�D���WV�c��P�$(��ϭ���[v�^�S�hZ]?+`�Rlp��4f.�{4��]���B�j��v�䮲��G�k�ל�� ���ڌ·����ӈz�^��LFG�w|'(��ܽ0ġ��)�n��Ϛ;/��?�����r�����@�c�l��^�.��[	���j�����|x�w�����G���E��I���0���-T�j�',.]��w.�_����n�Q�R��'VJՃX6a��"�*��Ve-��|9A�}��w�\�����V}A�ܽ a^f�f$�4��LB����$���k&$��# ���&�{Ig�w�B�XwZՖ�)��9]�δGί�49��~�:��	�%��$����7,��+��%9Hq�	%
�1�S��޴	�%�_�ld�0c�a�ο�z�&n�k���*�_ƚ�9����c	yG�il�#�l<O�ڎ���@em��,9� �j�E\4�+�k��=���|� ��������k���Ե:))ķ��,��t�o���<c`�kUɚ���	bH��<	,�|��R\)���[<4hs�.��_�d��{i��Q/?,����WQ9���;�Α+e�a�<Ǻ��%��f��>�!�	�T���65�0{�:+;�����^��. F��s�"��"�:����9� ��@*UB�֚�,!]�1\=ʧV�����)�n��,L瞨��,|=����;�t�z���p~��� TfHE���$��=��K�-�!^�X.��<�(�<]�A�.����>z�OF{|� �1�B��^&�������y�����n�E`�DY
������c�O\�q��rKؒ��	]��wO%-���v���P�؃wb�˪X7A���J�+�z�)�~ԝ�0g͸����8�9C�������K�?1A<�U$e���j����p<�U\� ��6ݭ�v[+�lxף�^�<�f�.�L� �w�W�wELc�k���;�r"�`���_����[$���-˭Q{H�����,����8�>�:�� ʌC�Ԋ�|�M�茂O%�1�M���d�§�N�?hB��n�M-� ���No7����{�>˃D�%m���wv+���\߾<].bHQ�?wٔD�J�?',�ġ��j\u��853�A٧_���F��fŋ����a��D�!�z[�\��h4㳠4��G�6|�`�fyz��U-�曽%�������߹���>���w��o�|����{A,2e���P�-��G��V��E��/�mb�\�'"��g4zh�^T��%�C�ڍ$���f�p[^��n�SH�H���ؤ^q|a;<��8b�~鹧8X������{�_�h[Rp�O���Mb�}�U��,J]M�Z�T��û��!�y��Q���).�
��v����(���T�z�`������ 
%=���Id8%�yգ��3¨)�%4����@�췬/�֟�[k�*Vxv��;�����pYǦ=��yu�b k�E,;y*�n.ʤ�bfm|Y�� �Z���xcar�?�@�Τ�qM��Q
8��.��C䅮vg4��s�̲<+�VM6���FN�d�'��7/�A^,��tŁ�I'��_�����22
��lS��
���z_Bߣmf�u������k� 	�P�ˌ��Z�wwM�����x�p�k��.��: ���'
���RK=��7��J�/�=��7}ۺ�˃�z�\��x7�&��S��ٟ� ufd7h���v�V��4�;�	��ICZ%iBM���@<8��7u�*[<�ņ�D���7���/D�u��_&7�J׆PDʽU�<�.0�βU�qKT]�1މ��&egز�6�Y���zX1aq���ݗ��sYEsT,��b>cC����5I�t�����r"��SɊ���tR�ȝI�aO�bOj�ӹЮk��V	�KV�����*@��uDnT�-��
tk� VU�qa{pE���VRQ� �S�%��w�.�7l[��Q'Z#��L~c���Nz`l������
����"�\o���0�8�^�����J���ŧ�;���̈́
�V��(e���W/�ʮ#�E���Z�e����,ۯB�	w�wU�V�s5��Da��-�^;�ŵ_&�mɏ��#R��Cd�9�����.����&��;p�_��®\�NE�0$ �D� �w��y��z�����"_�Wzѥ���D��L��|=��6\՜OnN����g��N���:d�o�z��];�0&2�?���/�k\�� ��Ƽ^%�"�(n�(������������v�<�����b{��;��9�̑�2jGX����Y�m��!�~"�?�R��e�ivW:2A%j�s�o.M�|�Bp��-�j�c�s"�s�7V�q��t�c�Y�3$��)��B�����^Ẁ���4B�a��g.T�j@4�P������Y�������K"^�d����q����+܁����g�&K�~Bv/�r��Gm;���/�9�u���,�@c,g��i��<�Q94uN�4��,J(��$\bF,��w��ǰ�F�.��M��QL�kfG�N��{��o��'}�$�HU�cz��<����D�\����D��z���ƾ�Y!��p�ɹL��'�QmM�V���Yh��F�)#Y�yL��@�i�vU�VkB����P��-& ������#��cim��Dj|�j�^q[:�c���3j�:��W&�N��4�ڝ�y~�i*H�� *��E��^9x'sj��_Q����V/���|r<)��6B���-!����pȄ_�y6���N��n¬�B@&׻���W�W�k�d��stP�T�+��5��~Q�����������(�ܗ~D�)Ȱ�w��V=Mpe�;�|T�"��Z�ۨP�� lk���{"���|��C� G`l������p2�?R2��Ҁ��u�oX���c�pVݤ�w��8
�y��è��Lʸ����&WL&�H9P�l9��-�uޮ�|;'6Q����o��~o�MK#5���Srw>��q#���N.���)u�;+��U��/!?�H�)k僧G���j��&>�)���k�׷ 5�l�tI��>�:��܉�}��}N+����X�!Ӽ04e��g��Iõ@�D��MAQi�x]�v0S�:�1�"��G����Y+dU`I[ֶ��/�R��MYgl��~�m*��aњ�����6�8�	g8�������yW$i�z�O�q^�۫�H���KG`�L���5vA��P6�|B��q�uN�U�T����]5��*`c���%z�U�&����
�����m��"��`�?�:����8�4Ny[p�g<��˦�4,�i��Q˙,z�צ�
���Ȣr30 ��r`��S"Z�5�D�2������=:�ҏqI�.��K���� �ّ!#�DJ����|4�⣹��G��
u��G���Y��o�GjX.'�#xa���$NV/������&���h:�^�%�h��ZBM��%<����OK6��
��2f^V���2�ٴ����[`�II�l���@Sr��	mx9`+᫬w�~S�?@�Q)��g�����j:��٤G~��A"�"�E�m�quP�h�HK�sJ R�q)��T��8	�.9)�C�yd�Є�8zWUtq��%��P�ؐ}�#�O�l�ghjӅ>.c��P�"r�S�t	n���mu�K�j�L�+��K"�
�[��v���%�GV����=��4����	y�#>J�V��0#�,Fո�1�m��cWΜ�]��zI�qm�6�_4��z/��X�c��.b��<+l�Xk����,H����0|�wՎ3��R���|��������h��քm����L ��J�[./_��%�_�T��4�ӑXO�rxs.��A͌b
y���Ih����(�3m5.�H,%��.��F�m�~e��6R&�m�:#���:V�M
���T'k��ߢ3/ަ�tffr�:('E�S�� P-��� N��ַJ�=�9���%�����M�7�P��V�}:Y����1�<�ʖݤ�~��%��y�v�i�x��7$r���Z倀��(��%���u�ц�]�4-p�BU_�_�M!�a����A���pU%�ѱ��܍,�R�~D�d�{�G=�m��ܧ]�j�ռ�鳽CL	�T�N6V�nbXIv���|ʥ"س���Hbz�uv-ƳUu.���T��:���&�	=<Q0�H���Uc�/��&�Wf��G��B�kA�'6����l�Al����B4x�XQ�_�V�8�
Z���О;&��T^�9�_���������z�?��7�����D����Y��tm���{8)RK�K�������Ƥ7��+|�9�l�ğ����B�h_iD"�O��㯻��zy�H�}.��@Y�> 9��@aW�.�6�����BBAV����X)�Xp�_�J7#��<<pp�]#�Їd/�4�h~T��A_۴&����{��RB `�IE�{�*�6�3�>����-��a�-�}��$���� �B�:r?�<�;�Ⱥ3��������&�����x����6����G�bn-s�㥤��
�GQ��h�:��M�l��ɰ��ĕ�-���������}��W%�h�}	�Z�=�ǚ��&�l.?SKe ���j�N����˙Wt�<�۶c�����KO�K��䳗>�I8�J�cUERe5��Xݖk �]�P�>�8!�kl�Ԍ+�'�Y��>h�F	e��Gu*56�1�h�!��.��,���`Y-��K0ԭ�(�#ti F���*#l|��t�Ϛ���愬ME-����I�������sՏh�5�G��8�c��6�Оr=T�s����ݦ��@�OO�5�y!4����# ����PT�����'�y 11RA�,�nxb*�L��<j̟I_.V��!YN��Ϲ#����/ot�rO�&�b�d(�a�|n6�s�k��F*���ZS%2�����B����&�B�.S�"G1�#���C�������?���r�\u��K�F"�ƃ7�i��tTS�	�V[+�{���t�3���kG�-"�X��Z�0�`���vY +L���fQYT���P�A�vu��� �Bb�������%~�2�=�5η�۫�PM��g�k��ߛ\��iU����+u�l�&O��G��/�[X�89t�~�L��T��e�!{���n
��z�4Tl%R5�*5���1 C>��?�ρ=x�~v1WG���;���572Uƹ.���=ۉ��>��Q���B9��M�Dq@O�P6/�P�Y��&B�S��bMCmJH�������t�g*�q�T7���<�+m�������S�9��Bѹ�|�O%���LBn�����&�<�|y����2����crD�Ta<�g�co�_=�Z�c)C_�xU�i�p6�0|�?8�|��0�xb�B���5�G��ס�U��,C�M v[rV2��fys\ޣ��fd*�@#�u�A��UU�P�2ˉҏ&�*����6ˬ����eNӕ$�8��-&������А��ԡ���T�4�[�12�����Q� *?"�|0$��JD�'������T��w���J�O�̭x���k���Ɵ��&��g{=Q��#����}N!��P�����Qw} jG�|����Ak���!-���,�*�q�׀{����R �c^<�,3rp�ı�f�Q��l�ꤤ��x���[�"yGM����w~�M�yt09(�daA{�`�]~ �ar���h�9��B>��A�F�&"2�y���I!�^�K���ы�7�A��5cP��li4�(�8�cЦ$�Ē�/6#
^�xx��Y����U���Y�^�D�\�L�	<�~��;V
���f?So�s��:W�[7�,�9g�Af2+�n֍��l~��?�h8�&�c�[��ZbC�l�m�V'��M�`����¡�O�<��?�0C��ㄶ��\2;�	�#��+=�d/jb�fYu�z^�J�Veث�
�U��Zҫ-Y{���(����K=�?	���A��;��2���]���Y��_�!�mz#|�p9�Js$��!�8�������m"�-�_Ϫ�fͰ������������Nxܕ�����Hhů
�`��iqol�Fz?��h�/4����:�T�ߜ�M��_�Ț(��e&4|������:'����:ڛ�"�%H��7�P�#'�'�Ğ)��Q���q��;��<6s���E]c/�;_�*d'��,��n���|��C�
k�o��T�C�z�zsW�n�Ac/�$K�=���1���ePC��� ����p�5㷛�
Xk8(`�`��҃�\�ZH�Kk 8�GY.�DKL{�rbf1����Idx0�]t�f#��UD�):�S9��s$�9�|a̱H���L�]��bMxH��|*��&�*n��}���-ov� ��s�1�/
]K���_i����e$��I�K�E�Z����*�@!z.1�M����J��$�C�`5�r���\ ôM+`��#v"�;EL���(�+u��;���K�d��I'�F��i��±�Vp~9���C��?&��'nVr�4���#,�)"���x���cҒJDyz���m䊏�ĩR�YL��C�(�6��X�i~Nf&v��E�b$�U�G�5�dg_=�ru��ړ>,�0�|�q)j��!��9�UH���^+H��>�+3G�C4�����򿃃�	zӳg��Ȕ�*��y��C�"����ݎ#����c�����5�8�'���:�����9n���D"J�t���>�u���{��l�j�gH����0T�r�\�ƶ*��uZ��m8j�j!��j��b����-�F�'�'�Z1�h�J�,��wg�
�Dn���I���N§	��0��*.�p��v{8�)QFtܰ�q7+��Xĸ�$���Q��V:�A���)T�y���l�I�����B=N4��m�"��3��$l����tB��ւ���}(;A\�K$H�%,0 �0i+*�bB�yAUCx�F�୾}w�Z���H�(#���y��ڙ�`f�CQ�����墆{f��}�oG%Z��,7;���^�g͙|?����G�\���C>If�E��N�i��9����o_bW��Ϳ�{��[g�,\���u��.�VeP;���H�W� ��T���[$���Q�E{�5���Zk�N�ud�(�F	�������Z��P�CC,�9y3)����U})�[8u�>�,�痠��.k�g��8M)u�B���W�ܥ�-y+q�y�*NP:�x�iY��i�"�	�E����ޱtT�so����zlӒ�,�����%w@f��c���ځ��������)�XE��Ӗ���5>��t�����Ϯ.z��K^�Q͞\C!�f�Yψ��
�D��������2cw�D�A���9��gZ��@3��㬻��ns^�p��!���z�� �XC�8xo�O��X�,�D/h���,<'�%?{�t��tÙ<�Ԫ��
�k&��[��a��<�z���S׉ޜDa;����c��X�W�c3?��)p�hPZ�.~ZTz��U�]�h����-//���gf�n�E��?[LNo���Z��ɕo�Fq	����\����>��e"S��!�,��G���&���yf��AYPe;�LQ;uL���]�7�<۾��\U�/�����Ln��F��B��qH�<�)��ķ�����O�E���I6�Y`��{9��h�t�]V��iY�3��W��l�!U�%�@M��v6��Y �@������nAC��T�,��Y1������M�[L���0�6�Xr���V���m��Q0�o
ݶ��E*C�!���]���^!g��w�����8#zn�Z�"�x��c�T���ڰ�X�hj=�X�x(���ci1�Wk�R#ugD+�'#��qn�������Gs���_�f��-��2)-gA���u��d��H���!�-qV����=3��]���kw}�`>�΃N��>6���Bt���!�����en|T��_��f~��;z߹C ~·4���@��&d� a���f>x��$ϫT	�����濅��w,���:B�.F��WA_���@�b.WQh�@�ΌR-X�����-(��;vU��Jm-����|%��;�/V]�T�&�4e�l\$M�pYl�h*�d��˔_��Ų��L9
yW�����Z��PͼH�А\��/�4����s�F���0���
����J��*�z	8���������H�h���\��{9d����+f�2����T��Ta �� 
8W�)�`S��y��  Ov��H427��h�϶ݤ��fJ�A�
{��B{U+������q���L�����c�hBf�=X61q���P"Ŧ~&E�}o76�c:�H��!U�$�����>��pQ��Z�RP)	{w� v�_�Yҁ���������d�,}�W�K݁�,2:$H>����2ъ�e�^��P[���k6�5cK�^�..���-��>8���U3�!vتu�ľ�����O��G�4��VP�FW�Q-�������<2SS��=z���͜5��1�,[:�b�^g�J��r0JՃ
G�c#��}l0?d��]&A �T��i�ۆ��̝'G{�肔Y��6�{vO7x!���ֳ�IǧE9K�g��+�1n��e���U6�M��Ea�I���&�w�`3G�����@C>6���Q�leIdpq��TLތ�v�t͸����b�$��9:hwS�����3�m��&���J��[�hi�	5XT��	�W �]8���d��we+wQ@P���QrU�""���G�,�MF�9��Q˰�o%d��Ct�"Y�*���˝�GrW���*cϴ��L�v�B=M6�p� l?>w�
�;qD��v�{�)��f��,�|\q�*�1qbָ��D����<�b٩��)\�9���lXv�#���.�pԴ��3`��=c�O`��
�d^�����C<y�~h���a`0o�=يƏ5�~�>g�
��$�����T޵���G����������g��Y
�H��[T�fR�û��0
	=�9�����7�d����o���8�)���N
���G�9X��\�ãذP�X���1�ƍ�x�Cot0`?cP�m=�*ş'$R Ufb*+iOx�ֆ�Ά�?vK/�|���,i�E�۽ϟX��Qݝ
��c������ٙn�w��4��Axc/�x��E�2I��O��\��dړD㺙t|m�8�ι�NOL��%[wp������l�q�*����؟����#��夙�w4��G)�V���_�8��o�3����V!@��5����A�"�h�jkJ�a�ݨJX3��e�eȧ���I���E�g6�*����r��Fd�&0��������˯V�7BZk�^�zfF�s�/�r-�62u��uL��r�#"��`J������/	{�+�Z!��+�T�Vu��vڀ���t������x���� �raޯ$6n45�aV�U��E^@0��XR	p�l#2���Q�M=^Wuf�V�v~�����*4����k��XJ��䰱�y�L�ˆ�ɂ/KR��6�[!������;���[84�K��,VE{���E�T���6G���P"�B{1�8Sw�n��A��j~�h�<1X�B�v,C��\��Y��l��f{�3WW�QY�!��"�pAT>�kp.��!*[�ίg|�������� lzAgt�W W�_b��eAF�)G~)��v�V���|��~��k�5�{0<�2�X;�=v��U0���z6Eo��kR�B���;����y4�[w�Bh�Ĳ��V�@%]�M��'}��1�3Fw�>�q�z�1k�N%��Y��$&���)VN�����s
)4B���kRl��=�y��J�����,j^�(�hTy2��K�T=F��1��o%��P�a�4�"qZkT���đ��3K̾Ϲ;�������]OR�j�~��a����I%Ϸ��+e��H��nay<��}��u
�����+��Z�S�����7������/WZ����8=5�rn�D���Ҙ��c$�h��m3��]� �͛[ϭF9�͊�0��ev	y̒�y��Q �q[�l��(������!Q�)-��]t�jk�B�%]��41V�4Ī�R9�ҝ̷�hU�lKl�#<��"}���|֐ܹS&���=r9ի�
D@ɺV���j��P��_.�ə�C�P�>{1d��W�WO��`�M�N�Ć=�s�G��k�>������xؖ�����+���a�t0�̑t'p�84���xe���at��e��S�+�5Y�e=F�Prǂ�����K0�i��ɐvjU��c��7#��� N@�<�_�|��V�|�j��'���i�ڴ�NN3����j�<&)��F��0�:Ӱ0=t�֛O� E��d�J�r���x�3MJk���	5��HpK����#���~�u����`ƛ�s��_V=�l�vdu!�i�G�Y��Yg�6��^���{���=hZ�y1�$�{�,�h�9͍ ��Yb�!��w!pB8,}���@�F'Ŗis'�8n�BV���Nl*M�B��7���D8& �zb��O���dœs:�E�������4'*�X���q�v����, �Ȅ��!�����4껤��1�Ѧ��6'H*ZX�7�/ԭC�seQ�#��	�HD<�M�Z�U��W�Z�- %�����z��\�C�%Z�K��!j֜�&��")j��OT���U�� Dn4X�o��������ـV�Y
���<Ĝ��mStz)�:H�S��≛!km{��������Q�/;��J�l������٤�nsU'���C����T[I��	L�#�(�S�0�n i����)�8�f� �D�n���G��s�C�_N�M��t���X,���J���ɯ?&����/�<��$��cqG�CDb u�y�	g׭�����P��Ѥ�� mu�Y�"
�c'd��qF,ճ��UrT�/�$�u�'�B�o���82-ϵm��ޥ��4�%T��+�y��U ��|��h���k�/Z�т�=�ˁ�H\$WrB!�y�jiM���-oj�3s���4|d��CI����A��]��é�MJXd� k*��ٻ��!�s�������`�9V��z�m��O�/�0�� Vj����{�<Qz���D�?A!#h�-mk�?�&�s�r*��P��S��ب������If�|�_��W�k%j�-mZX�3��T_0��!��B����b�N?�dw%#��-]H����.��h�Q��
3�Zk9�(��
v�l9L'(�$�f�@��?O�Xe
R|����q��_�W��A�b��DA�?9����mC�M�y:/�	S�)�Փ4���6όI�JV�t�X���D��'�[�L�-�=�5�(��58YE�*u�xhxƨF`aR�z.�O�-^��@ge��N��#�n'b��Ӈ�?u�oIE����`�t:^��%������o���]x	�=��Zw��!*�� ������|�!F-A��P����������!�[ߴ2�F��{ӏ|d{�Გ9heeχ�N�Y�c�=[\1�ZP��Q���siKW���e��{�3S�+��L�C��l��h�a`
�噌�p�#�ϹqCc�JaoΖ�~�`��'԰W���S��t�^Q��=m��r����	�N+��Hm��6Ũj�g�o?:����O��R�B�ě��M ��\8σ�bz��5���e��dyY�!���Sk�ϯP��E�ܥ���
5*�����/L��7��V�A�,y�L�FS�Cǝ��Ivk�9��*g�=4�FE"��
�@*?�7��Bl02S�7���������Zsb�e�m]����$�m���/ޒ���E���oR���� �$?4��3�k�yB
%���,�Yl}�����>����ݐE;�:�M��[�7Ia��ƽ��b�Y4q��~��4� .O���Z-��'~̅'-KW^��)W��2s�r�ZF8&>��,�mZ�@��dpK�~t�@P��ʪܜ�=��$ضw9��.6�ƾ�Y����`*��^BV���uO��D$�!�y���;��hJz��M�����>0�;�9��P�J���G�IX���r�b�-��s�L �#����,�}ȵ!j.�[7��LK[,��j�
�$�oÀ�{}�Ղ�q�_��G9:ļ3{|�'�BS -�0f	M�ʵk�-Z��e�����o�`��F����f*ɍy���A���@��T�%9�#9ZV��jc��ڿ2.K�j���-hD�+}_�}c�+�)ER�ǇL٦�	w��[�K��\,:u �P�=,1C��c�fl/�[�{o�ɇ��ٰ����c�yk��q��([&�'fN|'6�>|5��}��+���CR��!7xT(�"��0�j� 3�Β)�5�Y��iݕl0����M8Y�x���yUu�M��tO�~M76P�a)�� )�R4#4V����pYv�g��	 Q�=�G��h�Ʀ=���k�:��M�т��_ݝ�|X�O
f��(�f��� ��%�9W���ڃ����s��N��,M�%�͐{?�4$��K�^��F����Lz��q�V�?�>Fu�a!Zl�c���t���a��o(۩bc
�H�fS�������s�;��$~��Ą&����[��ν���G�&0B����/�]=�MVYn��e�p�}�^�
	Y\aY{.�S��/ěͧ|w�#Y���-�l��m�w��ݻB���zY�"U�Ne�|l��M��b��["��惑Vj���LP����<��Apk��-���J�;^;�l�Z����.H��P��_��P����\���b���nw	y^��f� v��3tZ৏�}�7	�0�hT��q�b��/�*z�l[�r��Y =��
���h	b�V9�+zS���b���2���	h���A')"�^�e�����������a�*�I�{�O���0���8����e:�y�dk1�3��u ?�:�k���Y��C��.ڬއbL��R2l`�C	�mc}l�g�z։����>���V_��ɨo�n{�h<fW!���t�b��rɮ�O���2���Lhݩ��q�BC�����#��7�
Wd������y�CS�5K�^���+�$�ǅFQ@�%�v�A��:U5"|�`dn�����yK5j\�
�z�+�8)��I�''�S���-P����a�$c�dy�<��m�=@�7��iK
[j�)�vc�%����_x���#��ldG&�-�@�M�
y���;�zD7��ϰ�Fht����,v&o�^3=b�be�Mw+XZ��v0Cl!�v�,pA˅7��m6���4/��}72��?��)�F�5qQ�M�]���ŵ���9p����d�8I���k<\���6͍�9�����[�@{#Lޮ�F��F*�Y�3���U�W �WTX�����=#�����"�y8v�\��Z�j���|5�ǂ�lD�t}�x\����#G�����r?�W�s��&��� j���̎Z!V��-x�L-	<I����c.z��U/�A3h(k+���0<���/�{���O�0@͝H�"��^v�@����Ef�����<�BZF��{���X[[9�˓���x�(�w�Q�o�|/�	�b��a�m̐m�T4�>~�v+](j�xK?	{�D�z�1��dӬD\���H+�R&b�;��4���>�aU�:%`����j��"�2ćJ�P��3uh���������_�uIh�5��"�G��֓�e��1@�a�R��72�*��z�Ď�͌6��i����< `ĺ�E��ȝ�4���GL�6^!��[�$os���	*�Vj�\Xy�2���\)T(бv?��l�x�sh���7f5�N��B�E~�)���'��;%�۰�Ab[��-Ǹ�{�q��ݘ�����z%x҅M!t庑����N1�|�DM$��� D�i�Ң��)l������:�8i$�R�h�ies�t,qa�׵mӉ�,� �礘�|(�� �˷��C;:��o�/���3�c<����
�<-*	��)�/>a��A=q��إ�;���uw�}��i<���Zw-]V91�S!�p(����0��`X'ɪ@�8I:��1E�a�i	�)���`�.և�> ��#�J04R|�X%2��ه���Kq����!�Ŝ�`�&R�N�kL�O�uo��9Z'��tn蟟dXP1����h>W�U�.�LL �,���y��f;�b�d��?�)���3` Yw�h��KG5t�iC!��"�[T`�tjń���ѓȷm�i%�H~@kc!6CP�)���z���*G���C�[v�b�5zp���@��;)�Z�o�X���\�	LZ~���h����ՂA.�q��Y�� 1�ЩNp~�5�B�d!��������e�:����:�-��'�]d�W�Q��"g�mBO~ㄜ|�N	F����g��^+[������ݺEev�S����:l�Gxx8�@(V�֬�*�g�[_lv��L�V�V}�~r5yܙ,��q�ؠ��'�R��/>PІ+M�'q��uiޖ��+!!t��a^�{���T[=�t֤$��}���ୃ�
���f$��yU�}K�lV1��i�D�����N�o�������<�"�nQ��a��y_]����CG�O�k">�i�N�� �G�_n?�}�����A2*����P̣r�rT��"�f*en�w�ޠq���e���V��fNvi��k鴒��\�q<�QP~j�>�i�#t|�)\�#�I�Xg�Ⱥ(���\��sU��TU�q����� �K%
n�D�䖷�S�=���# �-ˎ�!�V+IR���4:�5��^��Ւ�L���u@�k�R�\;��~���v����f���������:M�֤u������5|lCk��D��(zB돜@J�#D���=��a�Ġ>}�gx�CJB�u	�%��oD�����>l4���5�Ɂ�d2&�t���Ka�@�o?� �¦�7Y*൛h�}@�(^b�)�֍:Y���h�@<pW�����L�v�ۡ�P��!�Hvu"���1u9�҈�W'7�F�`q��W�e:g|��]x��9ӖBVY�������s#49N�>iͤ�|��`W��L�|5 �3�;�K Hj�Ê �eq�}c<
y_�{t��@��]���a龈NI�Yx��_4�6�5��<Ͳ$�!����KB�FY|�I&�Ȑ3�e�pj7��@m&=%+�? i_K�����@��e��D��[eq_��{v�Ŗ�B�:�팖c��	�D,
]&��q3��x��������|�h0�]��������������+�*��W\<k�҅PI�Ar�؈��J��u�Z����&{+�Q�����#7����{coW��e6����mM�i�֋̕'�K���cO5p�M�j�5ts�o�=��xֿ�5��yr�p)���vМWt��@���7��{���cvm������=�"�ܔ�|�Q����W�SMg��x����Za��F�7�rES߂����ny
p�79�u�J��f�66�J�>`�(�<w,�t$WN�tE�|r_�!bt���Ixi����P�B+u�͕�`lz�=j�bO��A�2xqs=�
������N4j+�zr�ڞX�O�eT�DE=���8��p�I](WX�EF "�Gf�\?����|�#�ߥ����D2���&�D��,�B�LS+μ����5�B�*N��=x��
��8��3J̷ծ� X;����aqq1$Iu�6H��T��1�\T�/�S�N�"�r9:����syT^敬��r�tOK��TD��i1��0��<�x��C�0K7)�e�#t�;�~ft1���{Rθ}nr���\�<��E�}4�4��4����0\
-u1'&P�J�m��E�;���AΗ�J���]!>X��UL�o��|�Ʀ��k���¦��/$.$���d�mx䫵� g���H�T.^hL"M�a�Е^y�&t'��w�<~�f�cx�"j_���G̝���B؅ 7�o��=V��RLrC����ط"]1ȴW~����j��]�!y��1�S�1G88;�^�>�:����>BI2�H�^Z�M��[
�Y�S��J�Ǽ�M�[W݈U�es&��殭�
��mgΓ�%w����VLZ�h���f�Ii5��غ�@��T�E7ώb����:% 贘�ߌ��L֧oD�C�ڦ�<�� N^p&��%H�-ʊ>����iB2
)�9�A\�	]WUuPeTȝ����eD�i�ȉ/'^`�)yb�Ė��s�����s��~�T$���S�J8�P�eL&����Q�j_{�X���g�z'� ����E68`��Ua�A��.�T�H��6�l���jB^�*�Ҧk����A���� v+�v\z���S��:�3E]%>feɲL���u?�}+��z@��s�P�?�.��Ր��o\�764������-��.��͟(���t�1��m���y̯[Lq Tx��2M*��p��������#�ۋJ��藿���� ��B"uQ*�T����35=U�����Q�.
Zj�@j?NG.���O֦(	�|��!1���ʧ 0&�,_��������i���:N�
����m\��h����bd��`ԬB�[]�01����~Y�c�߲�b=|�ds��� !6����5z{���Zb̲�&�"��7x#?�qa��c �/�n����J_̅;�HQ�a�f7y/ߧ�f-�/x�7�V��+ީwU�g� N �X���*�rMR��G�e�����5��z�ԟl��ά�n�Eg
:�5)a5��v�Q�g�0�n0dY�Ҥ����]�怡w��\�������G�Ҫ�L�8�RO|m6���ab�e��
{��1��e�/8²��|+���'}�6E.gHkM�lF>i����ֈ������[���0\�N�U���΍��	DP���d�HPi�:0,Xc�S��L�r��qx�í5
�W%I���Uv�֊����Y�4&��p������G#W���f�x�X���N&9-kdD
a��^N����T�hk�N��	JH���|(q~�g�,+�E�n������k6*p�uE���Q���D���x���:Nr�G����>cԉ?�b�y_{}�C*�\�th�$m""tW<[�z���������cw=����Ͷb�%�q����C���78컙���g�db[d?qS�{�e���9�-@t5![
����� �_6�x��v*��b$�#'�����.tSt�	&���9��*����Z�/�Hc]��.��UW���%':5-6F|�����*�$�e �Pم�7���M������5�Á][���L�.�8��P5��{���L�B�i���Ծrq6$mTQ/0]����6	�S�g���� N<(��?��;��p�[���Œ-2�3ff�|�~��1� ���d.{��9\�u�z��5[�Ji�����"z�Y��l���j��6L�����Eb0)=����:P��v9��ǈ�(��'�H.S�۶>e1	���}�ojK
�4McF������`��9�Wͻ�2@���!�pq�L���<��喍{���<�Y�*�	��~�"&�����h�-�V��& 胺�:KY����#_����(���E�C�j�3l~�-����EUU2S�"����@��﫢�/���HŢ�Q�~�Oo�hd��X������A ^`�ϕ@t9hfy�I�B�,j6\o��wW ���w{橆�������F��I��f�7:M��K.A��AȩG9�$�u�}Q��y�K�7��)[�VAЊHIh��X�����*��i���K�	��'
���`c+��	2)|5�?����dtc�l�jH��1�(Lɉ��C�AH>F����RMpc����v���N�W�M!�j�}Ou��ߺ�� �^��b�VK�gy���� ��ahzN;@�m%����q3x^���?;���n5H�r���e����;�7=Jv�'w�������ƻT��+6�D�h���8}�q8q������Z��HN��������٣���U��%��o2*�G73n#��ǑJ�칂,*Z$��E. n�^fEa��hZx�G� m�"tV�䌁��J�_*b1e�BOO$��w����:���ٞeg�'.زAw�"I���-���"G�������P�V�F����ۮ
?-�\2R������z$��j�����J�|ٗC%� p��
S��n���W�twr�r��溛LB��^/K	`�o�y�my��@�Qx��u���.Э㈌�1�`��~Ζ�m~�-]mc�}7����[��n��ä4=�H��З�V r��@���ѷ,��Nސ�8��z��ca���[��L�)�9��3�yW�t� 7�b	�שZ=�w_h�~k�OZ��#����D����6b��XW�
C���)3�a�T.X���N���PO���o�eyY�pXa��ese������k�%�ƋЖlD�G{{�yu�=�{��آ�mK`hw��v�Co��S��/�=91�p@虉\���UH��u���a"]y�V��}G�\�;@�k��.�
���}�%_?��tZOPE���?���1$iŻ�L2���iA��C߫�}ɲ%�w[�d4Cc�2�͋�=e��v E�R���e�6��7WUI������ ���/��2ێE3�Ȃ�A�vKi���w�ŝ��0ōn�Ǳ��(�U��[�[�Hf�w�J^�'K]�7����t�u�@�ĆH��'��锶��D̿�Z�7㝗v��5�W�/��ㆢj^T�.���d���/@�ʈ=D`7\�Dz[��q�}t��ڒ���p M��e�u)�jz!G띬AꝪ�`�@�����fi�ey#a����D8�~�r����r?S�k���jݨפm��\\)cy�2r{����QA�`I u�BG��?��*t�t[H/�M,�����Ǒζ���\����H�&F�K3�|<rds� 8��#R�h^��FZH�7�i#r��W ��/��6ƶbK�[�|�}�p:�(�CnJ�E	4аc��n�J?#�+qn4�4v�sT\����Ǔ=���*�s�{SHx1��`�ʸ:��L�*��)��XjKr�Q���Q�|i%v�S�9u
̐G�jJ>�E~E\�	����ʷ�T�n�-{w;���0�����9���7�jZf�2��L6����}G*>���x����-k6X	M"���@����E�~����/P��~�����J��m��F��+�i�v��u=�����۳�Uo��(N4C�ДaV9���➔>5�ƙy��t*��Ѕa�5�?J�ʫ�{��O�3MPQϼ��m_�rh&sb���f(=G�� �4�6��l��|��r���U��f���5�s�zFC����@y��e�Y����P���!"Wl��Y&�n�\mQU���u�XiW�@ԼO����ʆZ�p	n�{���l�I��M�(I�k[c�R��5&U���$�mt�a	(:��O����������J�xA�~K�cY�Ȟ�1�����À���S��ճ5{+��9lu�����6ҙ�꣢Y�>c�Z<eGp񛑃���	�pV*�����>����Y�ɶ/t?9<��Fo�J��7�J��u0{[��q�-S�A�1`�M�#.Mb==K}	+@�G@�wdt\��C$�-��X���U�@���:,�]�ا��tՄ��G�9RɰD�BT�>j�j�Q�������S�wi��dDB�)Q�����ؒ���A=0���cAi'�K��]P�W�O�ΐ���'��V��(׾�R�K�ܰ���[�~Yg��_J���&�3����C��ﰱȇ.�3�>8�l��D�mP�-�o:�g�P+�P�#��X˔��0�}� /��;W�,%��Q<@8���]��b�*W{�4�����8�`񦴡���;՗ʨ��P�s&���+�1�>(����@�b��	o��`s�[�:8��jd� 	V�W�#�_�nY)w�\�O&!щo�C'yK�k� ��Z��9�gdX%�Ę�� D�{ܸ���sk@�-��IϘ��O��d�����`aK���"H�PA4 � �&17���{��Tb�,�;\M����ڽ��=s�RU����y`��9���h�x������JE��J�:��!�^5����D��fj�*��-O�oɿG?�c����m|�/a�v'k]����ks"*F�Q��z����#��c�1D�m�oKG~�v_u��7l[�&�%b1:��?�S�4\E�֧���f�?t�>Cp2�ɀS��ҿR�����;)�'��tm�c����u��{�=5�_�ε�"_�B��u��_RL��sO����B=���\3����ؕ�B���H]�>�R�w��aL�'�4���4[�mn_�3?��% �k/X��79~	�ϒ_S��Q9�e���k*����"|��aC����i�1EBC�)J���l�Dtʬy���K&첼�j+�»�E\�h8���	���͝��q^��8�;
.��zQ�kjB�e����Ç���t�����>�YU(������x\��6;Gޒ��׾?��&��n���ڔ	���6�&&��(��C�4o&k��?���N>]� ��Y_Ƚ˃�!�Gl�0k#	I]��Q�j�hr�~�eC��2	.!Q�tX[������k�����H�D���*���;�n�Y���������64��}^��K����Qv�i���>��H[�Rcɧ�ܙ�@Õ��K]Fe�^vO�}-��)_�_��KP�m�.�DsIPz�)P盚
�eRM�C�k��I��4�Xn��ʫ�'�v��S����)2�7Ư�6�M�����P.��2�2w�ƍ�$YE�#y�1 Ɏ�N���	�9���v��f���Z泔#^\֙�E��,��L��Y��f�0�f?F��k��D��4R���=��O�Уe�}נ�R=����V��+��@������fƵ�
 �9i|�����G9�p%A�-�T�w��^կ�Q*����\�aJ&)G�����$��䩠��S��͹�焤��n�Ӹ ����Q��#M��$�W0�ݝ�«" �6�o��Zr�I��E��s��j���c����6��?u� ���1�*ud4�܊i1��붏��e].S]~�d9�\��Ꞟ��D>9%k& _����s�R�Ct&��mTj��]����Ae�Y_ת����R�h��0��}�J��l䨬���p��䲥�9 �eo�����@L�`�����"�=�[�ׯ��wѣ�7z�WnmM���k�4��s).�!X��a�M�ভM��b�D�LSM�Y�s��W��!g��`�0��ﻬ5(��CQ�y�u΀������n�M�;�V\hs�24Ql�h�s��fR1Hwk�tg̳��Qub�я����s_�^qW�#�7
/�إ�Ȯ�p��B����w�r$x�[��vO���B7�q
���f���Da��Beh۳&~X�����-^1� H���(c�˶� ����U�\f��4���ທ���~^�-B.�;"Q����MT�h��m�y�y��V��UU@l�eD�sˆ�@��r��鸩$��+h5�/_���*�i��RJ4�O�uO�Mb_���#�O��Ȏ�D�G��s���@ҔG��.���̉rI1���JsUcRE��g�1C�j�3W��ĲJ-j�M��[��
���Rc�ں��.��^ok�|��'1<@�	p�X�X�ᖱ�	�^�]x���h�sX���c��ք����;cS����Q>�F˴UK�<�
K��,TJ���|	��9�B�~EַC)�|!+�����l��K*5+<M��&W��G�:!f��\��f)�P܅��ձ�l�ͫ�Brjv`o?q�9Ns�W��̉��+��B�2K7��u�k�A�>��4�h� �k��<���+�)%d����s�����ۮ��s�º�ww��b	{�)C����T4�ol��I����u�e�ƨ��D)�=K��<�(m�э3�C�\JMA@��?;��n��4�x=o�_�.٧K�s	��puɢ	81?B��̛�Y;������c����lEp��d�v�mЂe�{������W�Rva"f6T|�q!_n�p���żS ��A��-|T����]�f�x9��a|�d�E7���H���q��>�+}�
Pg+�9
�5�Z�L���[#1dg\}�K����<@���o��O
tv ǳ��v��i�u��S�y�^��,[Ȩv(x�<�h�:v�5pɗ*���d� N�'��3�����f��n=�����b#ʓt'��� ��:P@K�z����b?����S����`K}�#n����qF�䯵�1`���Q�a�)9����]A|�a���[D+�E�)�Җ�n�$>������n->��_��UUxtu%��L�M޽�����m+pw��#���:�GӒCt������J��0]����xg*,"!��0���

O����Vk��E���[�;X�'M]z���f�_���f�25������E��N�&��?8���:�� �i
|�$j�bvt	�%�-�f���OVuS�n̂a�z���||�j���� ����a,g�$��W�Uw%��`�P�k��,�)C�p�����znH�e8c��An��z�]��g���Y{��[�(�xLj�	��|�K��T�i-_)nct��Zp����A8X���K��w}سu�UhQ�P�E���)c�����k;J�YH��Z	��5o`�̦.z�}2S�������ٲsOTۥ�����%���2SSq���'n	~�PBq����i@-�b�k���@��~��޲���&�;�,��sb`�?�j������0�ŗZ��)��F\��� v����1A��t��$3����6�n�(������	�&z+)[îJ�����q���n��f��W��^��xC ��%��<־,�1���l*�X͔���6�Y�	Y1�[7���x��%Fj�h�����;�$���f�qf$�kL?8�@뻧&�Fd[LF&|8��|O��$���b_�QV�8��7_��6D�]�Iڷ���:�=}�ZH��d�t�0�W�H\��+\�֋�2n d���o���T�9���{����G$;V��J�`Z�����v",rJxQB+�M�6�pV�=�A6�#��y�6AI�"�gJ*��u� O:�Qc&b맧�cHI���E��1�J����c����|����yӶ
�AYƭ�)����< ����7���ZC�p�N��jwv!���\��x�:�ԟ�Z�����he;I����{E�CP@=��5I����C��bǋ�9-&�%z�y�\[����Z	C3	3�,��V�9Pƞ^ܶ�,��-�k�')4��h�Z"HF�]`d��{#��"�#D0R8��G���Ef�z^P�7�?���X�C=?��>�Ј�������@�a�lo���f �="�6��&�ڹ9�C�#�d���k�#�k�ڗ+�Fn�����8i�d���K��\�"�t�u_U���x�~��3OO�K2�#6<�R�3�a��@'�S>���>��`�����
����i��P�HIr���l?����@��p��r��~� ��&mFJ7�ZU�=�M<�4��S���{M��T#�����ĆOZ������뚑3��g��R�oR"V��b���WBQB�u�H��Wr��#r{:s��M�#��@q�]�
M�$�t���X����Dz-ࡄ>�����M��q8��l�Z�♼{�Dv�l1^g]/Px�s��tD��꣫��A9�n��m�S�c[羻�v���]n�n�\�X�>Kܺ�I+��x�#������E�V7�u	����֘xӝa��P�VލJ�1Vҿ�)��Ҟ� ��Ty�B�Lv ����X����gU���}��5`Þwȏ��D���� �	ܔͣ��S�_�5lT��R�Ng1Q}"���7�}�:C�N���C�T��ue��[�Ŀ���pc�Z�[{`J�I+ \oW�n+$9���H��I\|�6��?B����;�쓏q!�\�]mi7�2�T� c�1�՚ }~|�jL����¶���~"寜�w[5���
�V�ق,8��&��/6�^��R���9h] �k����*O�p���*BGM�#��_�l� F5uu6�an�����m^����_yf���3��"���.�?���a@V��O�/�z31�8��?39p�5F)2W]���po�܏�[ȃ���z�/V1��T[�9�4�{�'�;�����A6"9��H;���Кw|���9�ŚX�����F��g�23 �b�����+G����۸;g+���*�t�q]���<��/Y�)��z?�gM�jB��h:eКq�;hw��liי2U%k	ynQw���L���b�,�0�rWu�;����	��+�$^�bg�$�+��L��tb�5`ǵ`��1Oޞ(97U��\���PJ��0���J�%�2�	�晕WS�vS�i�X�E�����5��Y���1OG@�;���T8��w�rWO`� r>��+s���s��DK��L����JV�ѯ�Ra�@��5�a/�~a�Y�"4���9:נR�3�Yu�%�R�h�$������e#0�&��C����9�	���|0���/o��N��8X:�[n�+I�b�t����B�N@�1 �XNw!@`����jeFb�e�e�
S��{,E�(�����A�Odu�-�HB�5�gh�]���^S�^5���:2�~(�R�pP\|�>� 4�CD�-�o��6�2 k�iݰ/ϲ�e+O���q������t����m}n�y+x�������KԱ��&'�M�����eS5/�'��$Ă0�"�t�	�(J�v��f�6P���7?p�8��jR�^߸�~��f�~���'����d=S��m>I�r���^rS�y�QXy��f8%��7�h��[�WS�gg~�� u����W�urd��ʺ���$_�r�Զ.1tV���pH��sq�V�({�z1����7�Bx�ʋ��=)��(ώh��|	��#�^�{�&���q�؀#��q]�6>>cIy>Y,����b�F	i�l�I<�		:\��dBh�4(�d�y�Y]�c�	�.G~�J;h�u3G�_0_4Wl} T���L�m6�;��D�t�Az��IY]�l^�8tα�Qo�sG�I���~���.��gwd�]�3��J;V��<Q��޺�M��.��ѧ�����4��!��n�>�4���Fq�z��4ԁ�!W0�zH 0��q%bM�Q�L�W[O�aD��7qwrv'�[����z4�������CxIj�(&��ԕ��19tX~^�_�/��B�栰:���#2�2�rF� ]/���р�a�%VP��du�����.iA,�;�;���Ay�����2a��Jzv!��\K�s�ę�/��k���#�'}�Vg�AZ�If�\O�%X�="c=c\NmF��ʧb��V�����ήt�*�(���%fY���1�<����'�}��UF�����!�դ���%2���.�B�X�B���[.�`��q�i*�&Ӌ���翹������.���Gﰁ���J��,y�V9h����ۃ/�
y��޸�&��.�4��{����;1�����#��I��9ox��"��\�8K/;,�L�:�@�_$�����ᦌ}�Q�S3����S��Z<g�'xRA���
WU��L)���\�!Y��n�rV���bd�W}��5�؄�T=�����nĲ��MO�S�����-�(�Y�E͖���;Q��&�
�-�#b����֫GS2�
G���FX0j�8쭓D󹁥Ѹ�B櫶o��Y�m�1Bgi*�`����u3x��Xd?��g�6��{ ������V/�v��Dk	��p:G����|c�R-��L��%�ń�m��׳&�D`�����ؓZl����j��A��r�<5~�٫��I9�	IW<0$L���d�
��c�y.޷ؖ��К�a�t�gu����ř�qa��N�����
���q {Kz�T+���@���G;h*YQ7%a�V���Tܠ��p����b���RO�I��אU����B���+s!���>�W�(�=�7|�P4��¡� }uӽ��z��Hz1W���������/� �$����{�� �����N[��6�z	��A{�=�Ĵq��R��KW9[XWb-��kڎ�m�v���(��\dg"�86�?g���xЂ���n���c
�������P�2o��A\H�������R�o��I �|�o^�|@��i$����!`�b���l��� �3�����ʅ��ZIQ�+�g!�$J��Gr��֌���?�i��T����W�A:���\�pu�6\"4�3�3Od[Ƃe�̔�
 ^��)V�tQ��s�kNq7���b|_>m��j�Կ�/6��@�������u9k-Tp���k���|�f��#�>��s�(����|�����O��(�e3P�_����m��=���V n���8�.��hU�\x�԰3���(v+M�����X�Lq0�K���^�H�.]�_���6��S����+�%��@Xbr*_n Av�?D��X �C~�b>��o�(�4f������#U�2�I�tq�i@�x��o?F"�;V�Ա_����,�
��L��i4f�m9qűFc8�:Ed�fe�o�&�|9����*�x�����0Z���~�u�i:*V�4�{��0�Z!-i��(|�����`�%D-�Ǘ��sR/���r��D+�����4���I!��m>��OI(ᣛ�m@�}��J��]괖�L鮷�j��Yd^؆]@"�^'�O�dB�)c��!`f�q*�/����%���qV���Ö�rM�l�ܙ!Z˅�δ�w
%��x{���$I@s����BcU��<��Ab�Y�A�H=�Φ��oq3[�q��Zl����u��5V+�@�!�G���l:�=��|�H{ʷ�U8p`�ʤ���Un��͟*��g	�"H��;�d����|����p�PY�8�5���:�n܏�)��}I��b-�"H���y���� �7�I.`��$^��]e������]ܝ� �v6�PS����>��P�1Rh%R�83�K)���pD3}"i����U"8!ؓm�!/mZ�'s��ǟ_�f���@�ێ�����@]��0e����Fl�����F0-��,җOIP|�9���j��+3���ۛ/�*)� S�f�ҋ]ʀ�)���A���Kդ��t�<�3HEQY�����ިu����J��;&Q���
�/�}VK�	��~��i�D�0���4�<S�u��x ��sֶC`����+A"­ҭq�n�ߛ-Ыc1[����-��f�&s�Ws4� ���? >�l�5�e�j�"���Ξ��m���7��F��ъ�<��r�j����c$�C�a�l�۫��"1��}��L����c�Kݘw��~XQ���B�V�{Hl�o�:%�9Z���
�q@!#��7�B�Ė�C�f�c�ء�x������e�:I@ݏY��cN���$U�D��-G���!5��O4�m�436����LC�Z�Gw�O��
��I�u���"����Ǥ�8̛�d��o��t}#�[quYa�#������AP�i��=�1O�6߭'@`&7E�K{��԰���ζ]U�lwj3ؿ:{o�t�ܸ{Ea��BlL�_���C��?�kp�߼/��)���M��X5d�c��u1_|�Jl؟2;?�1`4�Nn]����' Z����s��'h��*@��;��βu���01���j�m�^�W)�@�'2�)�IAM�/��>��_&�,��&�	W�D�0?)��&�&�3��N��d}���������e�hC�X7u^	�ME���`��j�;$I��^�������^���5��C^V�:kҹ6��Q
��Y��~kGD�怢������N�m_=ι�Z���ϻu��o�e!A�¸�*!�zfp�|�H�`7�+{�~K���ÞL��%���[�=pj͍ƼSZ�)b���[X�aܚ�K͍i7T��j�MЩ5�(�p��k_X@����a0R��k�dؘ4+��?���N����Ҏ��g��j�9%�$�GJ��&l� v�m�������>!Z��/�}�����f�Z-��Vj:|�c <6�9O2c5�qd�����Fm�r��1��Y�8��d�#����\��K�p���9��%�iG`d���<v`KKP.�X[Q��J��|7�u��5Q�}b��=�~`�]�v�JbhI�E�K!6X����9F{(�?B�ig�'LX*(��$�@?�J�D{������$�#U���	@��b�v�����0 f�/!��ǻ�p�͍4J���~3�7�Y����#0�6�U���gNPn<�$��"y��}u4�AWf�X06������7ӡ�saH��
*�`��F�5=�{aV
r�9�1LC�|���`����؂�^���>��P�d���f-"ܼ/�C2�л"��W0|�ݒ���'�*$-!_�O'�>;��pʪ*o�͵�.��I_��m�?�ً��XٯM���蕿:�^RO9�\4��s���o��	���j���P�����n@W�N�g�bo	�{ʈ��_I�[w�����Vu�`��qD8?�|V#������8h9�7񞪄񵢧,��sz����'1,�y�}5������[���h�W�����R. ��x�i���H1�)4~���ŵ|�(������᠏{
.���b 6�I�M�^����X�.��y{���յ)��%�v��/��30�1Ճpu���k�#*�&����h��=���P��>݄���2��w�:�t�����V~�A;���\���Q����h��)��є�}��`WC|%�J#q��-�ܶ@�+�V�Ѳ�`Y��"<yJ?���݀t������t�F��1|xR����X�z�)Z+&DܳaՌ/�cl����|)U5��%>;�� ��@��y|�I�����x)L�Bo�@����)ԓ�J�W4�S\���+*��8O�ň�S�A�d�iW��uc�Ը�(i��*�ҵȄ�/��ݺKKm�kݣ�N�1F�����vDw��u�P�/�Ǖ)� M׏ת �d�qu9�y_1M0�Z�#�����f��Z�U����I�'P��P�`O8)�G�Xg�1E����s�9K����Ф�0�o��͹`�CVY�`*a�q���Nt|h'3Z��&�z��O|R��5�Y�ֳ\�A�\��[Mq�q����9�2,�k�܊&���シ`ֵ���zXdxdbmg��`�b��ش�H�Ӏ��kK�3��f���l�T��l��ݜ?#�/LB3E��y��}3�6��w�3�2�v�,�ɘb����&���[@��6�(cr��)6ԅ��RX0�j�V]�1�^1�%�4ݮjq�+}C��z����!C(��6}Y)��u���?���G)8��\�O3w�3	m_��:7$��a@����~��OD;���w���u�(w��cwv����]�lO�tc�%BUo��DLc���(����[twA_��Tm5�(#	�����8��<�]�E���VL�B��I2�
r����~���N�(����4$ys��K����N�n�_1>rGa�}*t���|�́b��\v7�KB����Yr>--�+w *��% ��V8]V�cp{
N���#�V@p���G���b^}I���s��34B-m�4���o4��^������U�O���3��f�����E�<ٺ�Qlu8-8
Rd2�(*�Gw��I�A���6��i�p�𦋟l�'���x��	0�~�j� ߱�7���h��[��b��g�Sl�~d���/�n�,���_�v�O}�Gf��$�Tum[�HѨ�/�H���[O��D�M�.7ƤՆ�xt0�Ҏ��YTB��TK�
�9�0dXD��;�D�"v�R�&�@��cW�w�[k��b@U�R�m���;���u ���<�V,�hl f�"�5wδ�������_�%���길Z|�W�K�F�#R6f�
�IVtH�Q��%����]d�!%&H���{��!2��@��7`���<�@sUa��@�y��%W}����[�C�p���	�{��6�	P�r���.�����D���_�G���1B�5f'j8�Uu�2�M�x4v�0�����fmPk�|�rR�Q`
�
Ћ2f�������^Ē{�B��䰈�6�� A��L�1�E츦/�/�p2���p ʞo8�ut;�cP�/�QS|���� Ԉ0�u�^�T�4�/5̱������%���`��mP��Z��Em��Q����H ;�~�!O���Q��v;!�K
+��pDٕ��N�2Q�#��$��������	$W{gcרt����.�1��.ّ��}���I���i���9�"�Z�"<�8'���#kb�3��;o���<.)�Z��O�ئ��/T!ډԽ�������͎�BK_�q���x�,�|��ZRn�bRd?s���0��� 7��(|{���n�]WEN["w�c �Y|�����ě�"&�"Jj;�&UbR=�?�?{��'s�h��gź��������?3S��R"�����W��.Ƚ=݇xW����n��0Jv2��q�(o˚\+�H�� �b~\sUzR��6X�\X�FX'���(}�S9 9\�- ~E�eS�z����uXv������v`�&T[F+�����4(� 5�3U	6T�j��Jc)������{s
̶�+��}��,�'�;�F�l�s���1�8O��a�J���03�1�����0×��Z-r��D�3%	.q���.E�u���W�OvO2; w'lnF,�J�NzZo"[�[�h�`�n����^��O)�R���#����u�oB_Q��R�aF�td$���֚Rp�I��+�vjV?;���H�
�^><X	�v����=�KQ�M�q��:�c�ym�le�|�̴0��*����i3�m���N@"����"��ε��*��?ٍ:ޫ���3qd�}HՎdmJ�1�X`t!:t �'��p�OR�V��N���-�ū]W�f�i�L��g�X@4B[\�	%l[�X��r��u[M�eS������3�����o_�^']X�|F�pf���V��N���oH��:�����ZsG�KS!���C���"�'�"z�л���a�ERO�@�����|O����X�#�`yʊ6wp(�w>E�m�����n�{���]�5�Ku�\��H��
Г��3_P��N囆!�QI��J�\�h�.�n(#�U�8$���:��>Ƽ�}k[��]&!�z^[L�6_����V���e���< ��/���M�@j��՜�ᥟL+\�*e*�؆L�+����%�9.�oe�2�*���Do0��j-����Z�vdm��8�6���h��j�>2�º��_�x�D'�+e&Z� x>%�8�b��p���~W{�z��*�pUC�����2�%ݲ�f�[��\@��CF��%G�gS�*7�~�] kv��d��K�	#q��.�����7�������Tc-�>���o.�n	gT��]G��h7�)�`��Y���HRPJ��"���_)� n'ګB�7r@�8�5�{�-�(�T�#
`Ddw�匸���_#�k��� 1����� ��d���	/im_�|ӛ��.��o�@!��s�:)C��/	��}��&�^��ܼ��K �S�%B'o]i�����HBU�x����9��{����E13!�+-tg]���JD�"���Tի"������l�����5��Q[�{[��%�N|��u�"�s$t��r�S����>2nE�����-R��;>qrW�	�";����^?�c����	M6���V頡X�1_P>U��־��c_���j�.�!%���{��y���m��pX��Na?�bܞ4�v���P$^L�ۼ��tC=�9
����o��-���_�Sȯ���e+Q��ZmZ?�xry��㧷�� k�T ��΍�Џ����"ĴHK�ā�7��n�̓Ly�J�4��t�v��y�I~x���3�VJΑ�a��G���]��L�òY���-JY{z����ފ=z��k
fc�Dܕ���̺�dl��k5>]���G��`���~���>'I �q�@f���!�s�R�\9"��-1-ӑ
���P:�7Bu�멓	DW���:D RD92�5�Fҫ�o��M��6� �Z�F�i�q�
ԛz([,	��̌Q|'�����`�r�ؑ��ZA{[���X�/4��������*����M��Ϩt�i��`���uN��9�����T�����JP�П�#�$H��ӓ&2�ԁ�g/̈́��%dU� �N����It�Lw��3R�k�q)��Y�dxTTPH>��:��3�"\�'�}<>�E\�6#�;����Ax-} �`�on�&BU{e�c���}:6���hU���%�vM���+pQ���G����z���+(!Ay�o�Wӡȳ�c��D��3���i%p��r$'�1^I���)���4���I۰m]ꣿ?����Q��gqEN��@�;�vD;֊�_��4���0�j��#�;@t����*6��4s+b]�18��sD,�l��%��i�ֿ���u��ӫ; AZ��f������xƕ���.����������.8m��92=��E,b�|����($?�f�m���/�k�|h"�2{*�
��HqQ����ђ�o��[�L=���(�>=�� �d�m�t��ӪyA�8�%�q#���f����������u<Nq�B$eq���h�0�'R?���{���z��cH��Ѽ��Wm<�w�/�2)�)�q)a����;kR�>f���o�T7��.P��q��/�����!��¡��SsN���P6:9��S����)տ��~
;c A��\�ō��?��s4�E*��b?T��WT�-��Y���ƕ�e�}N���;��h�]�ʹ�3G;ƵA1v+�o���ժ'+m��R݉�蟪��YZ_���q�2��	�ڀ(��/H�����Is�V_����͗��{S��m(?�f#���:"/\��6V���>�民#6#w��{���E_�^�h��,[����8��|f�'V#��-`8���o�R��d���>����w���,�7�*�� ����
�9�Kw#Y=[�����T\�'5��Q�u�
�:�����K'w���⻶%>6�vP��@@�e!����v��B��9���wb�F�N���y�suȋ��b|�c�ef�P�w�U���T����^���iM��϶���J�{F��FEaͯ�<�b$�?{�+�����ҭ4�^���i�~Wno1�0�¶q������m��pW��Ԙ�d�.�TQnap�f/;߇p4�kTl%���'�4<ډ�[c���g]K��6aý&x4a��j�d�$	��X��6�ƹ\#���dh���l,����!�7P����O��?&�'��@�7Y���<E�=v�Q���ؙ>�Zu�*E4
l�S������mU��Y�� $����*R�b�4�U�h�*����:ݦ}� AC/T�ez������l����&��UڀD�?SܵT��;{.�-ː���7r���Q+�ު�T�v"��@73t������׎� 6K����y\�����]�N'7h>j���,p��?/=��!���YѰ<����=���zh·��RQ�7��i�P�_�,�g��'������7x:�3o�*�^�yjz�WSZ!0j[�� 4��I`Q���>�]�ɴ�O�:���U9�S6|�H�4����mQ����W�����E�,@�p�НC��G|���`�+�x;̊\����^C+)kTQ��R��Wkr���]i�&�ؤg�f��E<�h�g^�SRa��Ў�9�a�Daq*BPf�.)�uz�KƖ��Ap�GU�D���v��G�Ne�˳�8�3��΅A~������m�8 ��=���?��:�,�`������*H��qx~�Z����bL��W����9�[�����1�'Y<����K��R�M���R���{hB�[����[|�U��G
����An#Ms��d}c�� �֒�q��?0D�����X���o�v]/{�r�9�NX9�Mt�2�iB�k�͝*�i�̗�}�$�z��7���Jx����(�.��<Q����*J6���f����8#K鶡��]@�s$��u�7iSH�t��%�@6}�=x�����#A�6Z�e��r��/�|w�#
ʹ-bjw�;��y+�_��ҍ�j���B��*Z������R͙>�6X�g&����H���>0����Y :좓rU��J�a&��$d��f�7��H�[^�+�IM`f/��xU1瘸����Sk��#|�R#+X�����9��a�-��_WB�������R:A3���ț�[D4�ģr|�g<�1��[$`���[B�^����@�Wa܃U�rR�a�X}+��X��ΐ	�Tn�t�cZ����t�`��A�*��F�@�:��X��It�,�0hZ0�����N�V�M���\/l���O>F$�D@K�rX���R�0���H�t_���ȍ���m^2KN�����P�nF����w�7I+܄�+�ik摌@�w�]d2��Ⱥ)>֝��#2��$]�z,��0�vB&���-�A¾7	�h�	�9����h ��!�.�t��~�l�ܚ�
�(�n��A,���H����و�4Ń��lN���T���P���O�O�L�������4�d��ߤ�>��!~��m|֝��8�o Z�9-6zU����H�FЀ�{��<f&$�Y��@���8���gΛp�n~J��|���T��9�Z��b���6��y�ˤ���(��\D��[}��a}Zw}�	Z.��& �p�����_)���C�Y�㻛A.�-�*��}��}%�����U|�)grR�Z���	$�ƑTE'"֐-��+�'�sG�^�=h*�ۗ�ߣ���k�6-�c՛'�Iе� ��p�KJW���Z�v�H�4���x;M���΅[-�ȃ�|�~���2
�oS�;����̱޳�`z��)s�!��C��~m���}#����)ʸ9��M�(��)�\�O���]Q4QVFÙ��H�I'����"�w:�6e��ŷ�zh��F[=��Wq��TM��̚R�D0sgMXR��Ǖ:��}pX�V�>�|29	ާ.%��j�����!w}��͠�7�� *#E'��.�n�.g�Y[�u���h�!-���)��#��!n5�&�
��F�S��#ٕ�)�H�A�e�G���J;��2~/4/��6C�+C�FH��JР�4�tŀ���>M�߂f��@�I���D�OI5r�� ��|%\�;�!�h0���Ξ��k״f�i ���߃��SZQ^n!�x��j���{�+= t��Ҙ�i>hA��.Vօ+c~�o���B4Cy�6n�IAP��J E18���_EW��|�U	Թ#��s��|/>On��=��d-a8wL}n�R8<�rԥ���쎓�O!�]����98���+�q>��X\�MR[������ҏ�1��Cz�\�(X�\�������,�?�A���^�����=�0\�
��oG5}nA�N���ǽ!� �	7[[���D�ʤ���V��O.�O���M����(��h��%��ϔ��0B�⺠�q��`��ĺB��� �^Ҿ\
&Y�
�\[T���BF+��\$U�h��.���O"�vbG�PM2�j؞[l���K"`HI��W� 'cpYm�Ʉ��>9:Y����V��.7�������o�B@�[�h�6�s�	�"jw�z}�m�p*�V��p1<h�ز=��4n-NB&Jx7����/�ӧ|
�z���Ik��n�e�qƞnvm��af�1P�54\'o�j���L�*K+\�0r��J����ǁ���E���af�b��κ�0��*���bi�&�[f�T=<ܖ�o6�;�����}������4B�`C�O���x���z!�x'@��2�	�w��%�-2J�YS9ŢL�Z�=�~EZ^�RC>A��-�2j=8G�2��zg1��G����m��Jc���~�����8'��7�|��ifZJ2��s IS�MJ�B5�������@2��<���t��K���l5*$�[���K��ߒ�5>`��#��.� DUaN��M����
8�]h��}���d�[������?@Ȣ�5☑C��e<V���|O��� �h#."$Tڠ���`��o�p�k�g;�M���;C2Lػz����0{BAE&�
r��iS�p9��Ґ���_eM $�׉ת&[�D*
���eg9_���f.�+c4�_�Mn)�#�%?m�����sk���`�=u ���Hz��kr`�c��D.�p\�>����ջ��|LzȚ�w�(
�.Hc�mn��m�m�{6�lGc�T���l���a�k�� �1�5�}9XҘ�7.gJ(�����0V���-|f"�a_�P�wL�~���4&�]��],�Q�p��Mxԃ���/�	۬�����.�bJ�|����#%E��P���7�|�ǜ>(�*�Q/uY_�z�w�]��D�޸���P���	J--M�1�	�c�S�2t?<����\�q'��dY�s��x��wms���Hc�`_���?�U	�� �����Yɞ�Pυxf���٨�KT3W�8#�D�W�E\�ξ^�(�j�����pSM)î��$_�P9<.v�Gv4���`�ViI�Vj��to!��g�g�zq���f��O�?-��Y�7��_-��%���V͞�7�I{���[��S�"�qi�� �*0z���0��kmB��y�) H`�˚�����9ı%��&<��w�%�1Gr�����Gj���W�eF�vi���|4 3[����ܦq����ӿ\�u�� t�;�vS�x����,���B$ȁ�s��PO�������my��;��%���g��%һ��#*�%9�Һ�� �'L,�^��B4L���ǿє28��疬$u�8�����^n�0�g k�oO.s�n�{�?gc]����==S����4��B��W?�!}���&���r*c�8��!p�$�)�'�f�R�/�AE@���p�G�0�wD����*��
_��a�A+����\�Ep�q5��m��*7�̏O
o�i7��2��C�)��zD��k�g�"�!U g��ѯj�,����x�}�<��@Zs����$�ˬw��Wc��B�I;t��:���s+pP�ǯ�ܶj�n�ѻ�����y˥_�`]Q��쌹.YD�r$GI�V�Z��b/u nZ�+�S��/qg樲��Iw�9ָc&��qV?&&�'
b�����W�?Sc[,b���| ����B{�5x��C/!���']�� AtZ�o�:��o��������Q����I����;d�M����&�t渢S.ᵆ1	iYajm��zzG�;w���t���Gl\43~_�ǡ��I��"���ϫ�q�W0\D���@͗�`��5]SY-/s�Ѝ�H��4���	b$��k�N��f�,��GCU�(z?�w}6�I����\9;���_�dM��k�O%Fz3��(�N*#z�"�G�8}ϭjZ�l��u��aYW�C���*�w,��RܿC(y����x�ˏ�q{�a AQ��k�H�/.Q�E�͕���@j_�v1t���h���(�� �-�����I�`H���b_�yT΂���O��� �O:)
$��>H6��Ɲ�vGE�Ԏ��9>6�ή�"y��]hE�t$3��^
NJ�K��!�l����1��Ϻ
����u�J���W�]x���9۸����/J����yT0}g��i��;�IB�M��I�~��VE���ax��2>Y�\h;��&7�zmC�^7Q:�*@0W������z�wo�o�7��HR�n�#$�p7QS8��tF�H����b_������4/�^L�/�� T�ѩ���xgz�Ó��q�
s:`�h���Y"��f��K�'�@O���FMaz��S���5��]Q��W�t��2�<Km�;��Ԧ� �G����[�e�@�b�X�N�i+q�sh������ءHQNE6U��#|98�.���ܳ|���$��5s佌�vK��X`Έ���?N�b������/1̕
N�izs����D�ukrMt-��E�I�f|,7��E��Yu$�LN2<�h_]�1�e~��0+�|�"7lgJp�8�vp�xw%����iW�ŕ�ww�T��u[ 6�$����k�v���=o��֨H"fn�W�����bOi�Y	�,4-%!˫J�I|Zu:1� my�}Vs�üS�E��<u��r�~�a��nu� �ߙ�m����f�{����X,Mn���'6�/q�^p�����ؖM^;�����Y�%x� Kt�����W�3
���<F��Ėً��� p=�����b���1Q*�:O*������ Su@Wɛ�W�g�r3�����9�3����@�S�*N�yM������L/s�w�H\~n6N?�KR=y�C(W��qy��-E�&���I���YҮ���o�\94��<].�]�>��:3 {Z����J��Un���>��"�-Ow�%+�"���/C�_����7.~�1�ء�f%�a�\�ҝI�c�]轞;�zIwR��Xk�w��UPZV}�Z���%5S��P��;�)�"F@V�܇T3R�r L�ƭ?�>'�qߴjɻ�|���E�&�ۆڙx�9/,]/���[Z��bH�u&q�ȃQrʺ�J��T#c��M�s.x�;XC'bל������/RKs�2%Z�J�2#_���G�3k�9���~�j��{O�k�7[��
*A���72O����\���V�v�i����v��E���U6u�D!+d���߃d�&�Q�����'��|_td��.gh���P�`ȣ�̮\ڃ�{�-����IJ?�ǧ��r�o\��8�
�M ؍��Up<�a,�&}ވ�w�R�\�:��D�5�q�Z�N��XZ�H�(Y��&���`nt�2�5YT�;���xc�����ܖ�����������a��r�D�ӏOM�q1G� r�b��,����ɛ�	�ݗ#s���m���קKT�ƨ׺�E�Y�clfp *�>�T8�;hS�vY�s%�znp0
���[j�Oq��܂��V`��g��n	L�\��;C��Di����-���6W*������$�mg0�!X�_mU��uTaV�s/M&��#�X��Mtmrcc"�l�x�qwD��O	W�"���˷v����{]��4�@��\�&l�"���Vm��x(%xVo�+����bc��>^b�ɲ���1ف�m��
>���A總`���.�N�'��H������(��Ci]��	5�6�& q�L�֤����O� {V
�{Ҝ6q|��X���o��[�-}�%h0R&�>`��D^�ԣŲq�����1���Ɩ�<G·�/�P�	�k�����L��!��MF;�ڽ�\SƵ�N�v�p�E��).�&��wt�M��9/�[z)oz6r,���(<�����y4����m �`[���s�$�f5���c���@
�:�չ�BD����Z"�����)#z�_-	�u���1'� �hZl�^G�7�e���f��P�H�Y�3d�3�eZ�a�}yL���X�T�Y:�^kWގ�GM��=��m,�S,>�ؾ�|�;j��c��i�P;� �ձ�zb�O��;�oL��^����z�׵H����q�\aUC�ayS2�=��Ae�NU���]���s4⛙�h�Oꦔ@k�� �Y�0iOν˖�K�n��^�5�wN\�h9zXE0�י��^����yT)������� ���ݠ2ꅓ�Q^i\�̉fs��D��ױA��~
@���Rw�ɀ��c0��яF\<$Y��1r����%X5��W�M�8/��e���H�o]D�����e����.��v<����	��n�~TdH�:ӧ��:������`�3��x�,E���\�&����� �|�;�+D��y�O�x�3��@
��>�Ԗ�*�g;X�$��P�v��g�Fov���-w�hp��m"#T߱6�������i@ -�|~'c4M�h �=�Q��:�̘�)�l�����oW���j��n��T�mp(X���	c����QuX��}j�|z�*��l1�ex�p!��\}.����\\%�M��Z:<j=^�0��Z�����1���]/�V�E��Lԥ���f�`߾��GJ"�Z����X����Ű���W���̱�bk@'�I#�G�W[���?��7y��n���A^���2�y|�"��Dի��W�mǏB�Nn��k�d�Sb΃��@!A���[��V�ɫak7Rh�~ ޜʏv��H�ң҉�D�ka������qR��q���������FC_\�����n�]�R�pV�1�9����)����.u���	i�k��'+1jŮ�2z�A��[d�*^� c�ύP�����z��V��nÀ�+�;,(��<�~�R>�UT�fj�u��V���:�: (�y�6C2�x��4~��=i#2�ܖz)���C�齟���bp�+hX���@����/a����F F�̒�d��l��Uv�9����O�4O��tY���<�-��G�u`�&��d�Od�ʫ@"������eC���ž��ZY�v'q�y�`]��>���d���������D�)� �f�^���u�B�s��a�=o�!F{�|�r�E�υ��U-; _����qu��M#k�ve��d �*cG��������d�� ����9��s���^�;#ͲD�2�O$�I�����i�gQ�~��j܄Q��(�kJ����	�r]l�-�V ��mϹ�џ�%yy���"�t�jͅ�BDZ�ݣ+'�?��5�gCr���ԕ�J�x{��iǠb:��R)���^��eW۳��
a�V��*�0�	��y�j�4,���NN[j�-�3J���ݟn=��;R���&0�R�ږ��'%��L���!�A���3���x�IR�ft�h�qA8�hlgɇ���J
QL��h�g���g��Q�C�@��6��1W1��wD��m�PF�r�hU~��v�3�΂��
��[��K]3�	$��P��{�.Ӿ���!,k���9�\�v�*Y��Ϳ��MW�K�8��t�O�����5����\{6|��.����ƣ�N�o^�b����;���Ibm��U^bo�Eݻ%�b��w[�b_�xU{Ց,�b]��g����.�7��y��{��>� ŊF�rS���/����Z��Ꭾ��;��E��LԆ��z��|([�LWk�(�[�l�/��d�.Ѳ*�x��q*�4A���S�̩���%p���Qv;s8�)���;=zFt<����%��s�l(sv#++vy�oz.>��\9e�-����^��c��A�c�����J�#��H�� ~|4KꚖ1n��xB'��ux<� �E o:eA>6?��VE��+݄��}Z�K�$���ki����)9<C@�<��R�{1}���}�D��Iu]WQI!z� h^4W֒���V�霐�l��� 
%���}J�eq���
���Tr��n_��dO�^��o��_�DXP�X�_�7����)��_���M��1:��[P�lx� �Vt�-����ð;��r��%�0t|l̥l2���\�mCgyVe��B�)Z����a�&�E�\I�f���C��ڢ1�<v��m�η����m#R���������2�w��.?�0f��Ak��ӭ<
�b2y�J�]mP�XQ5���*N��n�|��^h?7w�[�&A�,+7ga&n�U��ϻ���2��X��:�p�+��۸f�|&��dԡ�82
`�H=@xc��X�r���$	Ef`�E��j*��X������
f��}��+l�1��T�Z,�4��W6��.ϪfAI�]�~/�)d���d*?� e@�RC.*Z_��K'"�D�cT�X=�W�誥|��9C� �������r� tFӅ�)�1Ďĺ-˸;5�7��g\N<���4~�;i5��h��F�Փq_�%/k��=va�����ᯕ�X�E������3�G4��hl<�5r��s��A���^�5�{3z���l�=oK��o�P�Q�O�Ӆ0��ݤ��%�� �q([��1�ݯR�ǯ)��&Y�.�����/�zDl��sBs�5׶���)��O�0�d?<hG�+��3��a��t)�R#��	�D���=ϸ}
Z|��Tü�u�!��Q�)W'�Q�s���8�[���}=KE�r1���w�ɳ0����]{Y9c�6���+_���/�$s�e�T*�IEo�UF�Ë?�g�Q��Ͱ���2�"���>�<��K� ~3��ՙ�y��5e@a�K�j@��%��@�m���[���㴋���G��y�,�wN5)+������?��4��u ���l�4��>T�~�<+	���<al���s�#@n�4�T�W�3��p�z��ܞ���ׂ w��pmUrQ�{��e�M���y3��df�߳s��0<<"#�%�����A�m&�W���B�e� B
!t��V��'N�@�/���B&F���ӌ��&�L|���
��"��Z��.��p
��e�ȯ�^�i���ڪ�WJ��X���۴�
��9N��=��c��I�.��z��r���A��*���
��� �_w��(��p��{=��1��s�X�f46텼����!�
ȿ���7������=(��Dů08���>��7��ф�����7���-oG�|�2����І�.���@ù��k�g�2Sc�Kӟ����ƅ�D`���1�j���D��h�}��",$[r�:��d6�'�����ZA�f����ZY�/9u]�����d���A5�'d��C��#Mشxb�p��^y)�Ǡu�BӪA�����.7x+�rP���޺6�s'ˏ�+�Ȱ�Qge��J(D������r����Po�S`��іR6���r���;w�E���+������*�ɿ�ۈ��1�x��c	���I� ~}� =y�^��" 㩑�Z0)���55.X�oOʿ4;��͏��%%��׹�gdl	V���H1���'��i⒢N�z��Wm�G�c��-�||��v����6�CP2�:>\���ч}z�g�}P2�}����R��^���������w��,����趐�3ᔋ�fN&�L��v($J����Ŏu�u�E"ʅ�2x�TDs�x�_W�uk���@k�}��Y Ga�$�(y���"�Nx+\�f��25v�Fy�����}�o���=	�pс��U�ǳC��5�=�XJ��:`�������ʀ�-�& B����*þ���
�q@�-_�W�f�	�!�7܆I�ըokk�q����3���7 {�  �;� �f�| �:���ͱv�N� V�Qۚ�1�nY���<�.��{1����L�O��j����?�>�1��3|b��x�&1���$2��+(��̂�����>r��}��O�_e�i2�`SX(q̨��O�۬z�LU��:
�@�]:l�~�I�13�+TV�|�>�F��ݼ�������J�3M^��iu��h֍Ddc]�� �yg��H���81�*KM`(� >�7ɑǅF[�-�nM8e�����j1�MV|�G�����E�и���h����,�=�r^�*��̝������ڍ3\*e�%�Z�ո�q��籀~QM5�p�;��QH����1`Ì�X8�V���[��s�?e�����b	�Pb���˛nR7<���)Sb��A"uF��O��X��>�(���ER��2���[�f�ΚO�c�n��.��bkx.k���ɱ�Z��<�#g�c6$�o�t�(���� ]?����͐X�5^¾�_���r��R.�fݻL�?�j�aj����M��uv�
(kTAI;�
����-�
��L �����<��P�Iʒ��/�N�[��tC�#E���mt�P��iݔ�"i��/�]����?�n�ݜI� Ąp��6�q�h�7�Gme]!dtV~��������d�(�Ru�o�m�D�bRJ�o��_&�����]lm0���`��_�:z\s�SSVRc��p?��)F{�=`��h���w`4�p�,׊�T. ��5E���)�O�����tKg�f� '~�SB�˚�������k���q~1�<'j�HHGB���tQ�y{������*n >��ˎ���c�@��+f�V�y��[����b�{>��pZb�ag{���t�$\�ŦB��W�2��&���55=!Kɔ�� ]��(�!�e.G�>�N4キ~e��)�`���nAu��Y����㋲�`��L��#����Y,��O�d��HOx��j�R��Oэ]�b:�u|��J�-�R��r5����mTʀ����,�9�{�T�܌�A-'�d����e�;
��"��}t���7�y$[�p㗎 �[���(
�y�3e�����=�$O�9�/���ϓ��"چ#]Vq�u&Yk�ohx��h�&�.];8��anf��J��oҦ}�^���9���aЯG�y��h��(�~d5|��a�e9��y#+��YG��#>X+��1Bֱ�{E�O���S�4��H��2\���_a3{��z,�ݱg@*��5������LxR�{z��z���&�5��Wt鰿��e-ϣ�%Y�d)u9���u�g�Q='�͹��@��L���|�I��aI���2ɒ���X��|��U��Z�	�F�����uZ�7=���bw��m���J�p��_o��&�K�4�B�pa��Y�}1p7�Q���Y����9����CQ;(!���k�����S*����.���٤��<M�kl.N&�^�g|õ��d����I�1T��1[�[�}�ӄ�bP��z�V/�ќ�v�g\�f��!�t��m�����Qy82��"[6����G-��W2�ӈ=V����}����@!{���h�Z3�^�7(�Z,\5ܠ�N�ٝ�n>��)ڰ4�,�y�f��+b�v��w��"0{��Q/`��>^	x�sZ����4MO���} �$��"J�L�A4�p�#����xiчJMxv�O׾�ћ�\eӮ���(�_��^0�h]%�a��Aƅ�O
��٢�΃�e`�gZN�b�L h�6�$����g�p�׽	L���dՖS���zٮB˸=�TTx���k�T	cP��i�R�/���?�>\�T<�8�E�9��}X_d��𨠛�b}�\��¸� ���7��#+U9��\���D|Ǚ�8�'X:<�^�,�J--Wp�m`	 A`�Ll��▃r�-��6�ȇ8u��
�!j��a˴�ꡓ�پ#@aA��Z�y��`�3���N���N
ԯ�&[a3�_��)\�/1�Zb�}�k!��o��'�7֒j����Gks�K�1H��	�n<��:�éj�Q��%P���	�3�O\����Ȉ�;�#�������J���^
���揯���ij�2��\��zU��Ɖ�U��L�͜gw����u%E
:C,��?ZkϮ�Y�-
%��wni���`uO����e���^�����d#a-_�|4��m�1���1'|�1�Wτ�溜�u~
���KX$�B� ��J�n�ÍB	��*0@Hy� 5����H���-{B��g�6 �t�c8��v�%��5����)n����2b&uR����X�J*�c�3䩳w�%���/�.&�A���'��&����׶�zQ]��˩���q���e���P���.�f�y��B8|6�/��}!�k�q��9:�a+*��<�>��DM^��,���v���0S�y�ʡT?��QӍ8��v��,�58TB��fn\Ņ�jI_�Zu�z�9�@�]2�P��S��)��MnWv�H��� �H��C�x��+<�s9n�Uݧ�҂p��?����L�v�ސUE��O\m�52h������[�WE�h 9養!]I��{�k�c�Ԗ���4�?3��^K2AFh���IE���T>�4����RVf��(u����zϜ{��2��6�5�K��잿I�X �������0�I�[ʺ���Q~V3 ����V�141��N�r�� �ŤND�l��Xc�YGpR��ߓ�W�Y\K�\B9��ˌYT���][\o�T'L��j��\�_dqo��
:�~c�Y��mԠ����~9��k�u�)J���tJV)���枔����۝g/8��#���%�$�Xsh�Z��@�z����C��үW^�W/No`#�X`�jk5������Z����ð�A��g�^���y䅘t2���7�VY��ُ���&�Y(o��`g�W::�+h-MNdv���T�^n��:�LӲ,��c���R�}�kp�����͆��`�9<�^��J3�1�~���~��;;|�)�mE[v��&f�B1��Rȩ.�$�	��:4��c6Y��b�޴�D�kG�B�I��n�,t9��-��-&����(������٪b�S�#�c�u�-�v^�ٖku�3��XaL��(��[�!\px�0�$ɠZ=�&��q`�.�*7G����Y�x�REu~Hi��dÿ쀈-tF�NBn��w��?I��2P��P^G=�:��-�~ ��0�����*�&%\���a�H�i@5'1�A}J����$�w���񫈼�1��F��5����a�� ۜ�����S�{
����jD}R�%��:nZ��B�f`�{�j��ׁR/҇ӗU�`�����ML�Z��\6s�j�$l�jr w��{��lZW>���=��K�.a�0|����ᇅ:n��p� ��Ͼ��*�7�� �����"��J���"$�9����/��܂6�^�4gV^�:�<zO>�
� V@�ObM�������zUaR�e���m���"���r0,�J;�`�Sv�M����2�5�4�HԨ��h��t͞���8���s�):�콺E|apD;�z��\��VF��<0���U�p'p1�������� 'Àd@��ÑA3F�P}�T���97�c���+`}ǐ�����vz�0<	,���Z{7/s	W߱�CecnqI����/�ot�,�\Ƀi��ǆWw�K�H�\�2���_��(�{�P�<c��@F�)~�8y-�����d���������!8 �u�b[���V���b ]�A���i��Nd�5-$�������WҐ$"f�e�/>z��cRƟ*����0V��N��p�����P}`l ����� e�Y$����`����H�ۚ)�x֜�f�G�'�D0q^Q�i�Jzł�q{��+{7�*#� �X�j�3N�X��L�IK�L9�Lj1ۇ�ټb��&~�d��~]y�4k�v���0��9V����&�\֐.^R2F �;l�'Pi��'@�����Ve�G�J�~����0Jg��<�ɯ�1�Y��6o^R�r�-@�^?���)xZ��=&�0ÿ��i�,i:l�#L=y�	��
��͛��Hl��.
��I^d�=���_X�#RƩ���FrU�e������F[^�����<}��lp9�띌��^D�'m'E;����JȌ�pF��%�i/e�i5R�MŒ��� �N�2q�����K�p����.����A#�!r!ҥ�D,��i1��Gk�/�6/G���_���}d���)=$-��:N��2�H_ah'.#N��:Z�'�O��C����;��_��j�sh�G�-�U�L���uY���3"�:f�7-GTN�C���!�>�U�f_�o�U�M�BH�zXD��a��h���;B�׍EM����S�[�5���=+�9Fm��v��<�����DZ"���������Ta�pը��π�����G讙TdW���#`�G���U���ę����m�. ��t3#�l�Z��O��!9#J}������x�6��"
O��}��P�Oe$M}wb���38�{Y ��$�4�()h7#M�ug i���M\�"3�1ҘU]�!�(+�ь��Q���tµ�.�.>���wC��j�'2����^5ʸ�8k��]W�E�R(t�����*�'��g�S
]v���񍈼ヮ6��A����8�A~�N��S�芆����AO��Z�c�[5e�(��?���D��4�4*<���LM�*�$f;aX��
E��e�6��� ���[C��=q�+�<�#qZ�d�
�7Ou^N#��g<@���mpK�N����spw�R"�oȆ#�h9�%���q�����O�w�y����z���z��}�sLxq<�(�@�~��:/���v�1��%��ѿg���j�4�U�	G:c�?=���M1O����Y �?�/BSp�͙����ߛH�f���ahǠ�Ug��c�s�#P�U�#���AƼ�8�w^=������g�ꤙg��`~X 
��vcP�?T\��ל$>׋�n8��g��ki�f�Y)���8M��$z~違?/W�q6G,��'�!�s�����8��i�{y�w�h��uu����e���E�1��,縗�'����pH>5� �6Sl@�r�5�g�:�߁,�G�s�����aK���T�Boǧӫ�H�3��m �Bp��9��Vc����V� �$'��Hv{jl
�+n򭄻~�ܴrKs p�9A��]�f�|+R�,����JD*���O(`^�B(�Q<&�oVA?�m|�a #aX��8�.��p�,%/&�X��nL��W�=E;t��7�6�Ŧq�,�!�S{���rb�Ȃ�C�hr���G�g�,)ԫ���,5r�ֆ�ӴAJ{!��= �*W��Ê{�MGͦ��,�A�˰Huu�op�M�)Nok�vݹ�=
)Y;����z��Y��bG�U�,��wj�� ����q˨��D��5k��X��i`����|��/m�]ǯ h��2��ˋ=^�%݈='��L�M�+td���,iI4����ȁO|�ʣ��Ao��Ԑg�%
(T���}�̾��Qx��cI!�ɝ���͟�>���^��Dк�7[u|�gW�(�������<��=k�ZsF�O%-�bA�ؕ�	'S�)�5o�%D�.���C*�Ivk�T�Y[�`��R���ŵQ�G�v��9`>P�:0hoA��J���p�)�W��:�����%��0j���4Y��j��-�
�8�S��~�	g�Kh�D=��Ib(ܸ[�����D˄3}�u��;�a�k��U��v��5�4�t��n$"O�E��Q����U��th~h��f01�}XM�U��V$L���	5�쥲+� 	�x݉bÁ Qf]�m&�H�d3~&��y�C���^I[��'��������bf#'�2�E�d'��$��q��Po��rj *6�Z��=Y�~o�H�.i�tX�6�n��*�9�ewB�v��,��:귰�x}K%)Gt	�vT?�JVBsܥ����p�#��\�D���l{�{��E|�������s�M��J`i2x�Mĸ�
m�u0'�J��P��u;G6����T���)h��E+�\S����{K�g0�h�!X/D�籟>o�r�s��˩����2��;F�����k�sm���Q�x=���:������l��&�1�O�x=���iD��mN
JKRD�GY*�A�J�C	�׾�D�N|�j�ܫ��,�Sl�]{�&!�4��	�gOm? ~P��e� ��$���Y���2?�T�r��͛��nקf���}S��I�_�nN� B�S��b� �\�+uH�@x�>���N��D��&t���� ��-���>���g�����F����&��]�$��@�~;eg?��-|��`b�n5�X�@B��{#�2|�T�%T�P�KDo����H俢�9�����5]�S����b��K�9��o(����zc"i$���
L����4�����/]��묓��N���x$c��&�⪰������D1k�u��>TU�������Hey�:��ʲS ���ڮP�L�!7�s�.Q��I@�Tx�Tkc�� ��է����I�n��t�w^�Y���7�d�[���44y�gl��Q�l&Uh�:������Y�{`�P��Kxt���(u���\��
�)߾�15R쏫wt�h�υh���������G+iE��4"��\��3<�k<�k,�,�éa5�$�&+�������,g�&<��Qw�C�_&������7勘J�'_��2�܋ªt;֒�ʄ��zͦUr����^6+�Y�®"����ܙke�7T>�}�H��bNB��H|��J��g�<��㌀,7����ay˓.��m��}�?�Z�M�[�G���������OM rSg�ksp��-K?v�OT��I5��?�s��E���qwD�^��I̹1�����~º�+dz"�q��p�tZ��4��ÜgN7w�KN|M_Q
��A R8lF"��7*~�ݽ	`�/Y���=�q������K������$"�5t����d���-����vZ��BO+����#��(�{��{���3Rހ���{�Ow�X�V/��?3�������b�Ҟ���Đ4Vu1���	\MHO�z�?��z��������Ǧ|'k+.�7�����=��²wq���Fv�6x{4�%S�7>,5m���S"�0�ҧ�]Z�kү�	r��X��k�F&Q�CY�%�@���<�'�~����Q�E@����¡��PV���j�3���l����F��U������o�Ȩ����?��Y8�~�m��'�&Z`4�N''����՘jÊz��=��GYbMؿz��ӵ.q�V��
��37�_G�#���+``֎�YRpu��U8/#1:5�3�+�V��-�c�BݽԅG�9�W>'�U���C�q]-Q�Qsa��W�̔�U�<�;M6�b�<��E��������J�L���ʌ��,�U��hGp�����~�;/Ȃ�T^_˟	��dQ�V���v݉ {*V�C���|��11xM��.Əs�<<�e���T_���~�5��Պm�����l��;N�� Zu�nf ;2i���%?��z[Qܡ߼�H�O9�e8�V��	�Q0�ꒋ��6�
�}��D7x���$E��ܯ����9���ذ��.��ڹ���Q�$�5 �Ԛ���ĝ�+;�=O甔5��O�l8�p}��*�x�;S7Cj�+۠#Ę���	|G4��j��� }��+Zm�V�**n��;�M;�3�Dvh�e���=B��|OU�vb~/�%=1J*,�l:��c�s�D�s�趱/�A-�J��>o�9�;��$ſ�>����{�&3���} �X�����^Z\ޒ�=�����+������.����v{��7��;��F��b\h[�i[�/�	�������%��n:��<�.Y()�L�ھ$�����5��C�QtG�\E���ځ@_��qgW�@�M<��DRa��׼�����M�. �I��͆��XAW�L����"� �d�;����~($��YN94�	�>h���v,V�z+�xv�D�	��%�6^��(��n�r�o������wo8~B��i�����)znr�oU��8�v�
��b�.3�K����Lمn������p�t�~2��xٻ��S�=D-�t��"0]aqj|S�o����u-�)��lt�� d�@���_ph\;*v�����u���3˦�rX��əR��0�<)2R`���'��t1�k���e9m�v�������/�5�]�h��7-84��a�~Ʉa���6�JFT���� ��LP�ْ�꥖�(��;բ��?ha�H��AN�����	�yn����j��i��XLtnN��0,�-�� ��~��a�s̭�\��&yCP�Rb�mCp����2YI�Ο�Ҙan�R$(��@+�/���f��pr �eeͺ߄]�Xi"y�{~�F�]�n��jBS���	!��e\�du�VKxpI��~�A"R;��;�۸����7Q�4�ʢ�ە�t�$�ׅ���*0c�f�F3��B�� ��"�k1 D�j[�$�,M�jgh9����*��m˽�Z	?T��s��-bp�=B7�0���%�ŋO�?e6�����cP=D�+�wĝ�cm�b���$"1�+���;������_2c�������m00�0�8��F���L6�yc_U(�J@�*��Xk4�j#��&l��0 �H�h��w�zB��0Ƥ\��s��X���Ŭ��j������#4I�ѹ���{)>�Z�ĺb&!E�x�3�E��A������=��t~�z�]�)-#F�h�=؀��)��UU2Lۚ�rl7B�a�u���Ƣ���4u9�'�)���5_u���8���~nbB�:�˕��iQ|~Mj�IK{l�5����q�@�
���G���cC��t��A�a��;�&S{bc���݁gt�T���Cw��x�}gH�� �on�\r��A�%^�{#��F&�S������5���y쥻�Ĩ��!9�EI���7��Nc������%�I�ޝ� �]�w�r�}VLoYvPִm\b�E�e����-^#H\"��R8�r��Q����>8����bL[�l=Z�,s���z�C���o�0��g���!k~�~��"Z�u�������8%8��F',B8��t8�@N)=��#F�z-V�5���������&"ET��ֶ+�մ#�9��F4�_[@���O	����m}%�͘�?\�=j[�)}$��:g�QÐ�a[��>�Y:��MX�1v�J��ģ>T�	C�2�kB�\�3�y�S�
=1�xw�V�O�;p:�@�G�@❰w܁�u3S��}��!g�[�T�,}��Đ0�:c��)kAN��\0��mhA�X��PGYjG��������9lEZ�%mKQ\J�[���J�x����j
�+H�N�q;-�E�?djM#ԧ���R ��[6�
���7C\4�����Q�O=�f8�s��<�=���{a�F�tۑ�BW�8�> ���r�8�Q�ͼJ�-�$ ӆ%��m#C��X���^Str]�����d�x��ɾ���d��E��C�w  .��C������|x\��n��+�X:{@u8�]�����;���tycq�㿶qgny�q?.u�[%v�%��]��Q�O�R�
�мSK��o�׳!��[����h3���$�Z��~b���F��ᒭ5��WD�p�7��gȑ!�V*!H�	?(H��������S5���'Zm[i���w���
E��<O� ���.���w� �{���I2E��I�.mQ��1��j�����.�b̯�z��(�X�E��߻|�b�kh
�sP;���	%|p�0��s�+��Y������}_�L��mt�Ȍ�� ΢��Q����l�/�1��ٯ�6}�dl�	������e���%�I��ч����V���%T^��;QS�I�l"�O�D�k��\������6Bi�A�=���*J�5~�xU�0:S����	
E������O�OM@�R��.TY%X��M�Ч ��b�i��?!�O[dJ�P �=c_�5���4�"�=x��'�R3 ��2������8��h�Z���mI=��'uyV�k�*P�۫����E�#��ZO�ӿF���%�VP������?����x
�cȣ���w������J=��%\wt�p��I u�&�]M�Ϯ�ɚ��v�#���Z��<P}��+R�h��?"=c��a_�<LAh�E�)$y��&����%k��5�#�G�A��=�f��1T'W�/���4���.���"��CH���D�b�ž��T0���v�Nx'~�����Ǿ�,}�2�U԰���������#����,a*���ϔQ�-g�H)s��M���3S[BZ?2`�ݐH�t�Da��X�c2A_@�IX�C�Fz�����>3���UC��Y�
m���rIK*�`H�ך�&}�v��r�֭���Q�vKŉ��qW��9ZAvF�X''��-f.��T�p�3,�0��辫X|E���m�Q��w���OߟF�I��F%�"r0��R���vѠ��x,	؊�ɹ�<�2�z$޲ԋ)m�^$/֓��S�#Ûk�e��"���(4�Ӿ%S�������W!r'aq��~]]`/HN����=�y��s�z>��s�x^7�@��-�|���L:tH�(��Q⑾��~ʆ���)cK��8��X��ϩ��$;��I���g��a�w��Q"�*����h����c#�͆A�z��U���B����O�Q���^LotHE�����m�5ӌL���Q*��xe���x��
 0�lu����$����l�/��u�g#kj�j���j6��܅�H�f��Hjo��+2ܻ�B��u�eςHv�����g$ol�@]W}6���<k��%?t!�"������Q�3)�O����z�P�;�M/"��ݪ9��#�&(�p����8U�L��[��g����$%nfM�y���6�)����Ě6�CS7��1����� ���FH�A�m��d�XO=Wj��}�[��T��C}�����By�
�2��;=�uCv^��r��w�ʧ{_���(Y��s���ц�6ԘEq)�b�"75c�9�IY�y�9�jkGl����c
��;�B��q�b���_�2�����WEU����S(Cu&��ژ�lhQo:�D�/���3Ҁ�ߪ�����^�	:@`�nD��TJW�/c�sЫ�ω��w��#����F�zq�� �9}c�h�� �$'�{�>^]M"aJab�q,��aBl�ᆭ�!d��E�SNk�>��Pz��j�"��L���.���Md�	�X&�"��kFU�ɘ�ȝ74��f��oYe�c�Ӄ������<ym�=��\��v��~�s�Ǯ\�ߋ���U(W@��) .-��yԗ�������W�d��;�ZD?��N���w\����u���8�;�JpA�8J	S7{��?A��Z�1�q�f�pDk��M�{�=�����&i�N��K���R��Ѱf|�Ӳ��BPt���ZbD�%�P�9m�>��v��Ydv�-�5n��-ze����8���R��a�=�b�A"\Tҭa�́��3Ѣ��2��$k����R8�8�����Pd�T0扈��ւ��"R�c���b'��\��oio�3��;�7Ʃ��>Ɂ��*7�+ <�>`��1fKbaY������D��Ω����3���+EY�V�o�ct����g�x/�B���X��l��nA���籏�y6�����I�+;V�ݚa��d �g�Lg��
�zji�4�����x"� A~$9�v�f���	��� ʼ�Bmv��eN���Մ�����T!�j��D���»U� �͘�
("]�{,z^f���n��a,r2ɥ7���xFb��9L0Y_&.�>U &N8,.���y3�E�8`@3����2�JȥZ���1��[�v5z�5tT��D���o���]��A\|;v�iQ���'Z�7��ҒwG�zHXz�L��c�����J���x��ܾ_-����% ��B w\I�Ra�D�Vr
�0��h�wt����e��5����Mx$��_�SwS���2Tt������p��h��ѳ:���p�y�:�H�F!�v�@��P��:��g~���ɋ�Bpz���fi"����ڑ� ��c|0�<��Q��;wx��D��6[�{]��:� �
%�� 0ϖ��g++��K'./z�P0 �x��5�FE�2�$Z�v�� ���L�"!;E0ee�T�\��Z���6��O -]s�*j+��`z�)!��b�����a^.ڮ߿7j�`�Do�Oٟ|����9��ْ�,XM���$;�o����n];�GQ�**P�@�`�"6���zh�@�n�s�U��Qc�+XJȻ:k�[|�+1�Yj����������M�ß���V�g�g�����۠F�:����R��
w�(��B�.6�T_IRL:�d��GKdf��U�_ᾅq�bI
nE��}h��6E�u��F�����NL픙�}y[�jtu�Ô�B������:�8���`�G�؋q{��b[���ld'���⁄�����W����!����(�l)�|X��P��Q��7����۾�$22lC��,a��6�R��{/m�+9@~��Z��\���@�
���g��$l���;&�S�A��!�T^��|��+�<!=_��X��ܳ�kG����������-<�Z1�[)nA��ʬ�w��Ûl����`����[ꁨJ{�끈�[��݄��c�k��v�)�;w^���9�c��ǽ�Kf�"C�Eׯ��2k}g��K��"���4F�AJ�a��`�4��)Nv�:w�L�����K�H��|��L C��4g�2�D(䋗i���F^&��}	$���Bjo�z���T[��2��~<Km�ճ�U6��	з�mv�Yd���������Z��~�3�X�6��^�~���AM@łjT��ߵ_����l��n�Su>������]�fVD.n��ȃ�ؽm͛�8;Ai9�h���5�7c�f:!���' _m얅ɚϢ1�iSy���C&�j�Km��9`ӎ9B~�����c~uNW,���-I�c9x�9�������-���5���[z��<
� ��f��X)�
��N(49�ixU]F�� ���I(��RpKg���k�1��e)��xp{���a̠����K�{/I6[>��n�5��h8`���&�/g�����tg-�Tj�6�}E.N�1uD���F�� ����=�gp ���U8����Y����_i�L�g��9��#�L)�p0p�#��h\;Q
�3qC`��o��J��\>�kL��j;�*�o�`p���� K���O9�5���S�	�Xiq�{Z_F#Xĭ?2yIWfY.�W�yA>�d���+Ɣc��-NSc�T=�h5j-K8�ANR��^���k��#AP���H�JkFz}��ȃ������m��Yˁ&9'���O{���m�5Q�d��r(�h0�-v|�M�&n�ҋ�1\�́�Sj3:�?Y�D���g������@[C�
�'$�a�+�aD��r]o^����<.���6�rE�4�@L�[�ņ��ħ޷������-�	)I�G�k��;�������
`�lD�F�-���� �+��-�x�U	��M���H%lo7��%gZ8��Jbj����zt���;���b_( ��H�%�o��6��k�r��ې�>b�)����f)�l���h�R����!p��#�����P�Ĥ�/�P���yIw�ę_D�B�؃�9[��Vb,m��f �G��I�$o���iN����<�&�}|�~*�I�A�M*@�Vo�z_�Hl=�-&P�.߬�o��6�%���,gq`E�����j�dπ��ȧ��`��R�3�-�#� j ���������MD4Ët��S����װ@���%��d �!�9�SR����S�lf1�+8j8�Ev+��!7��~!����CB�BT���3�0o-C`V����+�*�~!���F�����jEbCD��������ܷ
�rwRh�(�p�樯��m��/.�&$0���������$�D2f�'#�t$ũ���z��(WeeZ�OJ2���b�m7���z��)�z��ꡱ*P�&�ϳ� k ��aw�ǎ[��%�MGa&f=����˙t"�"3~@��p�����;��z�u#�f{3��ۤ��Twp�����~�P@�Jw�M�����C
�W�͸i�D��j��jl��	HI�k:�jƋ��v���fS}�b�&:B?����)���BpP(�RA���hX�Q�
$Ժw�{�L���R������шi陓v<����� :[K����J����B�J�/ ��U�q���M:Ɋ�|�bC~8�<�e |g2Al����D�<0�z�!�K;�z�W�̪���IF鴄#���4�eD;J#}����0�&��H0b��~�	<᭒�W�(��5A�Ѹ���[g9RS�,��ܤ����OV����->iXX0T�
��m�>3�f��k��FL!`�����Ĺ���iɝ�qOl�))�����X������%���̶O3\#���a�bz�c%rWz�>�ޭ$ƪ^�P!�!�����xU��&��q�Zӌ���e���2��4����o?�:^�jx�/���+j���߮�KY����k�e���n�83]�;�Z�K�K��6Ky)�Sk��s&���ެ��I.�F���}��	��(r��i�H^�0J
V5E¯]�Qw���M�JH�H��S)�@>�Jj�[���%��Z�Y��'�{�Ș�"^�� e�4Nuc�[�9`,1�3������V�s-*뛅�5�x�����T�R���ںUN�r�e���-]X��.7�o�R0��
v��5?o/:
.L��\�Q�y�qdBM��..�W�`�gw-�e;y�E@{?X���#���l��H����ǧ�]�k�M��/Pu� =�`�U�"ڴ�� ��ȃ>d�J�p^a[��!F�w$��s�'��|+��ut�-}������d(��03r����Ύ��1���.�ª��T9է��e���t0�ɱzL�51bX~p�'�ꀉMw���e/7t����D����d"�%h=�	һ�^A�ET>Nci�*P76�		?�]�>��K;��E���@T���o,�+����|ͱ���[!�0ׯ��B��>�<^��(?�\ ��/��س�x��r�}X���P֔�(T���Znd��"Z&�G� )�{��Gc(c\�w�}�F�ְ��qִ��8+�h�&^���A�c%`*�9跲��=�c|=�x4��W�v�f�a6������!8�l �@����)�U��柴��v]����Hf��P��$��~2��%o����	O�����wZ?q�s���]� >�Me�������d�Ao���в���6���I�4w}幵OJ���٪!�άw��l�)�ɉ�V�n�+4��}:l�P�,4m�1�2r1u]�C��GbkAi�P����_ײ��*��F���5U�������)���~���~�F/�fQf=x��'w|�3�{�U.��oլ^�k�ZCڼ�B����(����$�*��*��w������^ia\�IjO����4��S������W�m��I��d���3���􀡡��p]ĥ8��Z�8>bWK���W>��X�JC�;�(u�,��ѫDyn�o��%&8z���*ߎ����Z��2`̌��PC(�?��w�KD5�hfW�l�;O�������j]���WY���m��+�_-���Åĉ�3�@,�V+���c^ܕ���f6�[7�6b�f�瓘:�A���t��C�>@�}GV�2Q����� �@�ԕ �ľ�w7"�ma��~C�*�q�i���.w|�;�a�?<��c�+u�E�x�ˠ��	���!���u�/}��{���BP��N/�_�>)��=�]̏�\�� ĵ�9n_��#a�3[{�qa\X����ӧA0�#�%�����r��u<�ݝ:W/�q�ۍW�k�͡~,&S�ʈ"ꅟ�	��h�}��ju*s�c��`:r����� F4�]	xf�[K7P|��6�l�h;  W?lIg�����p���!�%�ԃC����
�*������Ϗ9sGn�\�39eь��u�����ՙI�^�[��^�}��H|.R/��_��0N��&\�����?պ��+զ9�b�u�!�~��0�����M�Td��2H^>��=���j�;��4w%���j����`f�A��l�y��e���eX����������??\�Zp����|���ݝ!��ջ��-cjb��c?G�Q�dݴ�CS�PuMp{Z(6yQU��� �a�X;���xg
��:��D{�sP�ˈ8DT��Q'vǅ���U㽓��E��q�%�1@��ͻ3|,�t��H�4$��hʭ��@`��ƕ�N��X�cȔ���[���.���E�Fa�j%X�]lrKt�'8�ڤ����
�7̡�����Q�]N%o�)S��ޅd�%|#]X7QIߵ͘�툪f�y>�w�DC�Ɂ�8R��]ESmà�|@��j�\݋?�1�]9/�A���1Kv1��6�8�n��a�`Sꕭ�S\r�Q����S��C�S@�~�p0b������69 =����p����|d^�Ǘ�o;uW�;5�t�W�4;i)�WO�9�Mhz�ו4]�h_�X�!��֎�?cŮ�o�q�_.��ݣi��W�����E�|�?BE򨤍���q�M���GGr�#�_�~��9F��B�GA�S�8)�xۑ�U�*,#�-�Q�I��v"A���nq��vf�y�Z����3�t�bȮc�#:��]&T���j;G�+�]OO�6�>�03M0��rDڽG��*,���1o����'���&�ԡ�2�M��z+z��>#8�e�e�F��
��<���mh sq�o�H?ƅ��U� �A�3��һNՕj6� :�!��2���o2�m(.M����a�y�Ӂ�>C��B6������-�I�㦥�
O׬eT��M8�3/HB"j�F7]8��\Kn�����Q�Z��P0��5�)�i�Q@$F]��H����F�*.��{?�_G�;�&��QSu�Ƕ?XAW��A"ȶ9\v��q_���i}`��Q��'�#&O����u��m�4��G���*>��ٶB���T�Xu��ԗ�������ZkRn�y��'�I�*f^���AI����|��g;�<[/{	�2��2{�rJ)��m=�Tn��x���5�1(�$h��k/�|_��izBm�Qvs,��[O�P'[#���PV�8&�^C�l°`En�2���'amL���`~O���#y��nvdM�����+��Y��8f�`�5/]B�|�Y�.nf�U��'��D+�1J�Hι���a���t�n7����%M�g�T���I����R���4��.��7{�b��ڴ|����Zi�uD�}���i��!@ʒ�UEo�"	���Ps��u����:�Bg�ף�\�5�Ѽ�JoU�H>���H����&����ֹ�=MK[6�\2I:�%�)�خ7~?���X��Ԍs
8e����TyLd��Bˋ������В㴬���m�0S����ad®�����R`&�PMr[� Z?�����F	:�{�kج `�@	��I������g���=�T�/��"Oh��F;��[$qw��[�ƒ�욥�Oq�et�P���/ʡ�d����#nw�X&���M���G����ܮ$��8#jW��Pt�?��ˮ�,�Y%�~�w���Foܚ��7�C��f�D��kZ����I�]k$��R����i�T�Ap^��w�L�UȽ௹��Ѫ���b��d�YŢꦾ��r8�bq8D��t<^Uj%���/E�pঠπ���r����J��Wy���>";�ݕdl�ٻ���eR-'�Q��S
�/mfV����9ђ�����2�g�O�i��-��^E�s�����q0�\�_�k��e�1U�b)ژ)u&/���h(�ys;�h~��op٣G��z!&���FdK�V��V���t�A�8�Vmy<�8�6��#i>=Jǟ�hW���#=o�2D;��2�����ߟ"���I��B;�k�x T��͘��w�2mב�W���M`�\�hD�O@�C��Y��Ĺ�I`��N\8;��,�u���>o�;�l/w:��.g���xȓ�У���F[Ry� �=�]�Z]+�C�V�����)�S	&�}�9�x��k.0�����If�;�d�[�ȥܧ�4w�ҿ9�:�����BNP�]F��!�;��W�������*��0\��E׍o�mU箚�����S�5��h��%v6���4Ja��fJǐ4��6���r�a�!W/pJh(YA�����%�@�:���}���slTn��K��,�]K�X�q�^O�fQ���C��1F�a<�ѯ{y�t�m�w�$TM� �ˏ��@��3I�y�x� M�J���aVlzHP/;�x�Z���?�>�w���V��t����I`�������kn"n9�ȃ�'�Ud�����2vq;�ɿ��D�>��I�A<��O�ޡ�����*�zQ��?w�C��bv}-��l��T [1��|g�i�m��A�N�T��8�%����b���E!�@GUr�<���O+%����+��t���}�B�$un����JL.ڵ����`22�����ܼBmY���%l�A&%��X}�ϠM�'�嫢�����*.X��I�F���Z�_����M�y��7����޸�[
}�W������Qܞϯ�<�HοF.��g|�8<��,��T/�*��E: ˲�Ԃ���ӡ��s�2�ƕ'�ܗ,�$�%�*?ysB"c%��.���<!�JȢp;����]�0��@/����܋9O;�HD,��6Qrl[vI[A�v`���V���.�Z�\�IѰiz������U��"\~��zP��VbV��X����ȓ�e��3�$�PnN�ت6L��������2��t��?�ş�/����m�)A4͡h�����d��d;T4vW��ͷ�^,Ac�D��2��&�<�z$���_*`4�? B�
������"�:b��8�jC3������d���T��0B���#/���� �A`�'DK9���1-T[T1������#�&ސO�〹}�B6UP5-����W좱�雁�0��Dh�JS���gS~��01N�͎�G����L��;>���q:��ɴ,=S/��j�䲐Γ[]s��ۅ0�1���f�H�Nأ*�_��*�l����!�Pp��)�B��Wؐ�/�U9C�bo�/��JP�iUs�X�tp���P"4��"�!�=
�}�0S~8��,��oj��w����kE�O�ϕL|��#��4�3�v
]����/UJ���gl&MD}b3:� :���;�X)�+��M�z�O}=%w���'�M�K�vGS��u���O���&=Q��'�1�ǈo�?AN3���������Z�l}�P,���	�E��NI�}�"2Ĵ@;���m����2J�E��pk��ۼ,!N����s�A�'JVK��}�#�	��Z��DP�(���H�7��S����Z)iK���hp|�i���f���"��ưSP��a|/z��
��N��/YMN:f!w��)��C4&���rt��0mg�;^���ӧ�[�t�A3�ad/��p��ˁМ��h�\�q�h8�Z�$��7���E�g�J���C%�d����6�ِ��E3���_�|Z��9�\��¼��¤��μVA9�@QfB+8 c̲6�d�Z�2�']�I�6�c�n�ČޖH�8�0��P�M���%���a��v!:��,;�Ek�wpH12�6��l����bԤpfj��ݳ)�&D��7���U�-*��Ol�w�/w	��vg���9t zzɑ��(���ҍ�z�)uQ��M�i*۾�Z�#^���ߕ)>�*�6Џ�����6��W�~7��i3�c������_�N/Dk��0����Wl8n朳jɵɝ�$S�Hc�_�'^��x��	f��d�����W��PٿO�i{���wD6���y�T�����&��+�?u8O1���x?��
+���J�	������.�,�^� ��-��[O<�s���(��3e�!���Sp`��zJ>uv�����y�nm���(��(���.I�t���#T���;��8��枥�Y�>�D���A���h佼3e9�<W�� ��h (���ce����zB��;��{V7����S��:t-2���y�%�`u0�򨴣p�U���$��k@d�I����A���Q2��a�@�0F�U`�,�����u���9Ր��@�>�a>�r}
9�.�f�F�vKt�/c�~7E)�n��D�c�b.�	���VWs`H�c��L���eU{CeS2Q�u�n�a���w�8�ߎ�C���&��8���"���FYQڹ���H�����3#\^W ;��lД)��@��	ʶ���:�)3�zt��?� Voʤ�|��z�4��ҹRU�܉��5�gE:�<h�\f�<���3�z�U\z��!ǒ_iH�Me=@�C��(�BQ����H�_���g�p��e���#:0�8�ֹ�l�1��2��qɼMA�s��\՛F{>�#0e?^�n��G��~���ǣӍ�:1�dY&,�f�R�r�p��(X]��jd��Ą���+��K�b;ڎ&	zM���Y�S�-wz�!m�b��qk�vD�mdբb���l��T*|�P�P��H͡+�@��Y?i�N/�Yq��w�s}·A�Ϩ$����s���=����8{��)���|(7Lذ��3D��g�4` J�%���bQ�?���۟o� Ym�,ƫ���EY7��XO(h��p��[�ꥵ�X!�#���T��!w����O5ҩ��{�FD����7��0'�V��E�H��l�Y:*�CuU
U��t$�w.=�[����p�uj�h#)���U�T J���s,8B�M3mj/_]�b����x���S�m��"�Sz��L��#����_�C��Б�'lM������b�ӓmm�[W/:�Z=-3�z�7d��#��B�fr1o��	x�����~�o0�Jh�����j-K��!��v�;
���¬X�j ��=��,��eK�� �УQV���DV�������9�Bd�� ���E�8"���돲�Q��F&,����nǒ	A���!A�hL�������E$/��m��C�V������g��όtN���
{a� I�N��r����Kr{̸|L�ޕ����^r�(������\O?yK}O�����䆈��9��oEj��|�8�k��cd��L��A�;u;�}�t�}�w�#i�����J�Y��f'ʭ��S���ꖶ#�Om0���B ��gBn#��9�˳�?� �+�dV�a�������9� �͝4�f�e��;
�
'���/%�|tf��p�%�+����ɑ:���2��&�P�P�7�,���!%�2������"#�[c�5�C	Ee���3" ����Ug�'I��S��;��iXv�d���:�D�L�����3
�/�����۹z��1�,�:�k�]nP�S��	��S�R3剏N�}��!�~0�o�7��'�(��"�e�R�)qYQ��VWǚ�>�a�Ļv����6z��G�]e�6щ%�O���[�~���r���j{+-�>�<X�J�/��VXSO�o]Գy&���O��� �+������l1�R�a'�?ׅ`���N%���
g�k��'�F�� ���,���<(�l��!$ʜ	_!́�$̯j�dq9}�隣} ٕ�|�AHP���H����񫍍��cFK��/�����V�buK�(}��3����As7<0Jf.Y�� �M���Q���k i<�X�'8�%K�Ȯ
�~۠enNZ��/���/R��,���dis��I���O��4M��02p���d7��1�ϙo+M7�ƾ������(0cW��5x�������jJ$C��4��f��ç�'g�{�h�T�E��Lꝗ���D�G�v�Dj��f[�cъѢ]b���QD��̪��E�L�1��e��Ή��u'���);��*���l ��-;�)�>�ӂ��=��Q78f��X�0I���[�%=h�B�Kt����s�{㉾���C�yZ9=�Ա_H��j��Pnr.��q�;�hr��4�!�P"�r�[s�fK�A����b�j�{S������̦���aGѺAя�f"�|gky���m�v'�Q�'F��nIǦ�{��Wx���]������W#!���YĜ���g�ेz�����b���l+����]�*��'��J�~���:b�U'�i�����{���Lބ��
���ݚ<��>Ռ;rE�5[�j��|*p)�XMO#��+���p�T3}���=����0�l>IH��{�[��Æt�b�L\��T�e�H��,��R��kHGh�D�i�Oͼ��]l�����)�?�;B�@���$˩1�y����M�Yy��u�M���̡����>|b��������ч<@K~�'A��|��{Ń��|X;�wd$v��>����	� '�N�@ɮ6�2���s5u���z�����kV#x�� w�q%�x
��	Y�d���%�JM�p0	L����p��4P�U2�Y����bKe�d�B��}H�]�q1m�`�]j��J�k�$����I��?Sl����5,b� 	�3���gm���I��F��1�]'Ք�!8|��:�oIJ����0�l�;Lw���Mx��9�N�'��J�=�ɂa��P�\�F�`J@ r��S�=�>��1����P���@t�c�%�>�*A��}����w�x��:���_}�>%�o��zM{R$�!��{Or�jx �6��ݾD���C����K?��YHMKy~� ��Q�/�\�^�A>�V���)yE��T�<QUK(E��4�nx�ȳ�n�_'ץŁ�7$^"��a����{E�9 2��po�!����J�j����h�8��	V��hLĥ/ՎD�Z�ǿjZ�;��C��AH�$�Ս���'F֢l>K�G��cG3�E�+6��������	[B<�,Fa����38�����,���)��8*�\�H���2y|B���qw���!L�Vnσ����A �,�U��n3O�l�����3RJ%9F�@�S��La�l)y�6��=l.ZD#�❤ޫO�{ĿV�M�OT�n�s{����c� bY�V�ی��`?mn���$B4 ���!B�-��ݻ�� S�9�]��@����;��nv�F[">!�(_�/��$��
r,RС�r�z�A�$��5�=Q���N_.ݿ�H���b������E9�7!�%�T���zkܯO$X��b%S�1PC+ϳ4�ϸ����� ��e
�)���ƚ�su���C��5x�{
�'Rr�yg��W𐷩/�)���&�����و�%بy��ܐ��9X�Z��ƍ6j�ڳ�K�PU��֓�$k�Y�x,�A�&���Cr�k7L�$JcQ�`LNW���{���Y](���@MI��7�C@H�A��B<��Bӱ�(�ZK9��CH�;��ִ�jq��J
$�8ן�ࡋ���w"6=���O]��5_���V�H�t��	d���I#�5gcu˙i�<\��~ݫN�A�C$}���a�<ށ*�թÝ0IPp|��J-r��\��b8����W�����+�F�{gCR�~�p�l��sM�Y6�E�%�}�����dY=� ��!T踚c-s(�m%L̚���������e��~B ߝ��b�<x(gXy(= 9�)���}�ɸ.�me�0�|�153�[���s�Omq���D�ޣ߾����Ow�V�l �m}�%�
�X�v,^wc���oB��F�ﶮ�1�sN�i���u���!X/%�ut޻���K�vܥ�����V�M'���1�%����t��!���U����O�g}�=�]L ��ݧ2��Qᱱ���U�_`|� �\j�w�dl���g����&�a?�.m�Ha{P�Ǔk�2�ľ�Wz���L�i̮���{�۶��u}"�E[@8�7v�K%0 	`8&X�n�"j� *ޮ���ͷa?TX^����̋������*�G�4�,�MF.��X�!�hѰ\��pd��	 Q�3�_���nC5!�NQ8n����D�R�,6�]v��b��A7$#���G�c�Q���^�x+��^,Ӟ��M%���	Nc�<�y�YET3��4������х2�����cݏ5­�yN�g_a��.3r	L�q�uS�,���q'��|f��@�G� ���4���0�! `�����0c�q�E��7��=ӏ�C���[����*�`�������
����)�������>\�`��0���D�Q�N(�`�D	��(���"�T���г����h��g&��L�|���}�:d�09���LFR�X�=�_�H�C,VW�z^ _Z���=���Kes}Y�pҭFFz�M�钰V���R����v�%�#�ؖ�d�1����h���E��UI���Wh���Fd̀��RJ"�J��7<N+��<'}K��"GЍ�\F�*�P|�?�T�<�����C��!����?�+�gY:VzWξ�����bUt��&���|j��T{˔i�K��"=�dH���M�*xs�ه�g�Q��� �#��b �M�aHɋFs���:��٥fɣ�-�[�f���.-���/�g�!�?�9�\y�Z�ѹQ���J����MgC���S�"�-;�W!Q.�,�O0y�*����lF�>J�C=���h4�)%����1\�������r��V��r��a��0m<�nw��v'{��@���9�~?w>��2��f%����B�-�yH,�4�1�%�[8؈��I�S�&��zá��C�7y��%�{�:���<��E'Bɾ�´1J2Ё#���@~�	`}~�\�I� �)<�;�g��&1y� x���<�qkaB�d�*Ǐ��Xh� �㌎�I��mk�1�$T0�C`��N6�F�Gqd� '�$K;��ߪ ��F(�t��V��#�T���9PCL�Y�Zu�U�N��m�z5�ה}���w=�cl�m����M�b�
�8��gMG�C���@yK�T�hB��֫/a:��,I|8v���M�Z���%��'sƱт�PX�U"�G��h�ҫ�&E7��
H�U}����
�r6���5��/B�*�
�'��F��;���AL�]�U����Sp��T���5mԃ�gui��"����d�&~>����,����0W�읡��P��P���ן8�N�u�����š%,d�
c���hOt� ��6�+i��w/�VyT"|�<��)[xM��~�!�O��ky14�T�L�
���1$�^["�R�@C�9n�m�<r]��H�L#g_^4�27:wWK&������s�� Hs�N�?۾��!�	>�����g�PW�EO�+��A�+昞C�.@Ó��*�KC�*�Q�RI�&��N�O�:��Xx�ל�7�F*��|D����䎪Xjܷ��tt�|Ds��d�:}0��w+��2e �g5�������3K&�8Q�c+,��
uX7�b��%_/�������+�%8�}[����Qқ+{'?gi�I�1"32��Qfees�H��5�D}�(��FO�H�U�r���{�?�e��f��QR�a��%��Az�X���#��А�����EΔL	`k򅂢Ҙ�3�A�=���� g
����	����Yd�Fb�W	���c٬���%+P�	��ĺ`Npʵ���y�u/p!� q��t�$��������,�a+k9^)���~>�P�U4����t�z��I���IYZ��wi��9�B��V���'��H&.7�6~BA�!���i�2�L+RF���V#��Ƃ�R�r�/-:z�"��Q ������$]�.�n����tj|3aR5ϔq���p�p{���7���A�ƣ��me���~!-;���<�sǛ�� �׎Z&=��U��v4�%�hOF�hNN��~��u9��$��?馮&���!�j���l�c:C���i⩿ҍ˛�n�]�,�Å蛨`Ջ���}r�\Y�̱]0T��d�R_
 �{6��w�l�D�x�n����b�Y��B��9�I����}�N�}��{����h]1D��ez÷�ZK^3�^��ӝ �0k�ԭe0�m��챦�%�� t<�� ��K����
֮+~�bX~$�Xߗ�l7��#V�gm�@C���(����hU-8QY�(�^+���-�h�'�����n��`������%KآR�-��+ٽe���䠷�$k�ђ���k ��JD&-�Ƌ٪L��L�i�z�O�l} ��{�"*�=�"�T���4*�����;�ߛES���`�2�H�ؙ�_�NI_/Q��$xD�*�"��:��v�����9��u�ou��Vˬ $����nFD���&N[}9�Ro'q�|7�6�
�ʦ��-���n{��&�	et�����/ar��P�<�;�MW�#��sՑ����B�H��ЎR?�R7�59��!/`?�)\���i�'5�]I(�����ر�Mi?(�2t�P˫�=���1��l�m��o(<`n��ր�q�Ma�2��20��F�F(�*�v#dEtdٽ̈�|�����j� ��~��Ts��M���XN�O]V,Ph��ę id�Zq�J%��Չ�}�2$�̛ �����c����/`����J��]� �	XAs�zOK�`�]�7�@��v���dd�0hu�9�U���Lj��;����^��΀f(P?�x�����A.��JB��c��Q��O��j�H�x@�C��<�����adO����*s�5��N|\���g#s�k8ȧy�'��}H�lH����ñ��C&S-7�5[�t0Ď;�m\	YS��1��mB1OQ�t��=c?�}�Q#��նa�ۥ����+h͊��i:�Pql3��>3�	6�C���c���n�\
���b��{���HE xȌD����8�w� ��Y�ʷ�XA�W�+a+�p�A
��x~�r$$W5�_�����DdR(&��j^B�%�_���2��f�_^�ɢ��t�e�pq���kן��y:lB����lZJ�99���܆s̱��+��j܂�7@�Ow ����`Ox�+/;i�{#�j���^g�P)<�x%�a
K�1��(K�k�g���u��X��z�Rj����ٛI��- �Y�}�����I�C����2g�mx	�^`ִ]��+.�⦥ZPD�J����~�0>B�ê�3�:k�=Y�>&�g8镝L)^�OmD+��VU��^G�d<LSb���n���ũ������z��	�D�1��]"���Tf�Y�.��#�� ��F�Y���*�\�������[,�#j'[������:R<f,�ř��f,q�T`��u��J*P����� *��l;����qu������m��Il^�sF�*��_�P)26^� Q]|�g���'�ܝr}W8�5��,�s��E��@�>)Ss��QO)�7�f �O�
��i����7V��π���?�Y�t�l���{��z��;�����B�GA�׏nD�����iTX��`�jV��5Fǁ�M�a���C�(V��x�\qg��Y�{sU��-�l�l���r�bLf8/u&Bz�nMg�i՛��3u  '�dH�g]���_��1h$U�!��P$��Ԝ���OVyS4m'_3�/{Ɛ	X't5U�ks
�C>0�=�M���-+A�ODm��W�݌ܻhC{W���tG ׎�GB�+��3BX�@���s�C1l��;��`��N_Kx�t:�+�G��q.�%f�@$}�x��/��%���cL��n&��XۼS"��R�6\)��;��i���ݔe�=W>�*�c.v�W�\uq���>i'K�i���Z��W�(VjD�y7B�y��M
���f��������H�ۖP��;���ޖeJ��(�->���xW����oq}�լ&�/Q0�Qʱ}K��e��<X �qY��mo���r`̊���)��piWZ]��j�A	n��@�T9ŕG��ʃ]���iCCBԽ9�G[���瀹?��P	f�5���0-̨��O^v�K�����+�`�Q�E�3͈B�ŲGlQ��ըk�I��as�'���4Y�bw۱W�}�V���Y��/2�}�#/�ZBS��������?Y�}��^79 ����~�q3�t��q� �m��HYNA�@��C1;+�M�Z`;@yX��ꙩ0�"wx�>]��۬��[|�VJ�x� 3��4� '��E�'X(B j���ꇗA[W�(�/�zO�K�IķG�s�_U8��@ ��}�kd�3��aq��e+}[��qz�xs��ݖ%��6��<��(A�]�Ղn�lK4#��8�ut�Q \���E^�y���m�k����\x��Y�ȆI��)[�������\�_yY]ͽ�U�W{��rj�S)�s��R4�1_�嬭�Wh�o�BwfB|pў��o��D�CK��@N���U���d��B��V1Em�
��toL<�A����_���i4}Fy�-e���4�!t5�3� Gn�֜���Ɵ�-LPVqad���,���d���z�U0$�ZO �5��������W�(��A��e�N��J�Լe����G�	h�N�H� ������T��?�b�('s���H���(:� )�I0�"�o�FL�;H��Z��E���˝nU�PQ�B���Nc[	�x4�\wA~ ��h�,���+YWhQ4��bu�7��L� �� aUh%��U�͡J�^�ϥɇ�����9�B��<u~�B�43c$������-o��V�2��v��ҋS�n����7��6 �+�b�Y;(���0:w}�������̐/�f��W��c���ti���U�8���2Z�,�=��ꋫ��P��bu����܁:܂,�z�� �G#��T�
�j��7t�:ѝF�}>,=�DT~�+�L~��~8��DҴ�����o����K U\���Y��׋�-n�2�$-P�V".�ڊ�5�� �򵢒j1Y-׈�q�~��\e�<φ�J��Q�{��+X2�;
!��C�»��?h;Hb>�F#(�O�?�1--ߓ��s:6X��;��@�ʏ������G$]�I�z�2!G$�=�^M?/�r=�*�
�gS���{j�~_ٞ��މ�jz�%x���7���7����e����ʢ�}�L����{3 ����T��OոY/3_��3L�K�6f��G�vA�|�m��;�Y|��oD}}�q�Pm�j�=ӭ��6��y�Wj�;j�8e�jt�w]�n僾Oߏ�e� ���e!�gF"M0W�	��NY+��ʵɢ�Q�����l�&vkja��[���H �NAL(1S��b���"���O{3���<&�ղ�"�(>ֽ��"+"��1
�NW�?��M}DI�����	h�g���]'��/&�E�AQ�`8��N9f�]|�	:-kL���=T���+�Ζ�2�9�2��ޣ�Ou(b,�@��@�+�u*�Q��\�а3�6�k0�:
dz�q-휮&���ߐ��:�k�kY�O�CEY�I4��C�0"����2X�ꎿ�ګ�BB+�f�Oj�u�wS��}�v(Ѓ��2&�3V�3mȹq��� �:�i+\�=��1����yH���Ko
��/��S��|J��>���Hfzs���+��!c:�g+Ρ�샜�t�2����jx���A�o,#B�\�~"m���₸��>D�O4� `�����n[��<tOքp%'*0�֬�e�#^�k-.5������I�b�W�+������iK�.�Z/f�?��qN��r�%-{	���Tt0���o�<(��]"㳡�Xx�J�3�ڒ%��0H��K�)(�R��YZ>�
?�蜐�aH�����g��=W���ًhz����P��Xt"�
�&�W՘���ROG�� ������W2��](	�^�8����V��f�W����6��Z���r��Y�5��O��  �e��Ď%�h�c�9 �=��3����ؿ��~s]�p���%Ca��6�}&!��z�]�y�yT`�����D!ߊ�6� �B�U�Y��A�#�P,a��A�e@�l���<f~w���xS�	E����N���h��Si��;��0��}͠��t�N�@�a�b� S�;�1��d���X!;���J���X���v̫���@��Q�KJ�
�fg?�G
�8�:�p:8UD�y�f�e?�eH�tm�=�e�F�{SD�D��f�j��)$Kٚ:��З��Y�ku���.rCL��c�I2���-�,�n��Z����$&KR�b��p�bc�l�1���Es�Z�`�+ky����t�p�f�3��m6��w�ԁO^��݄��>���.�[i\wT�q!cSX�H�(���bc�?��8L��4�/i}�N%���Ӏg��[pRϣ��u9c�#�i�A�P?A�32U��h�O�! ��*����Đ%hm8��6�!�|�����70��4��ɔ��1��v�f�ykLghv�}�mg�Q��m��2P�>���ly	���(���������k�x�:�Yg�AE؟Լ�@�-짊��X��x���H�
�&;�+Mx_�iگ��Ov����1����M鷚asZ+\�9�F�2.p*������U��X3�-��+�:MX�S�<����ޛ2vt����h6�q���z R���`�^}R�t��So���E+ ��b��o��d�v��rG�� l�Q�V�RJ����O��;V���>����]	U�B3<0R��"��(4Ӏ��.&߂t^&}lr�Zn)u�b�4|�+�s0��(xLL@x>�����X�5a^��k��D�9xh�IʓR��u�����6��*��v�+s]׫��hZ��W�xj]/m�	�۱ܚ��j�7FQ��ih%
��
�~����z{#��:��AQ}[�e� y�:�g�4�P��y,Kf��:����˶(8YH�rU�����M�������<֤`X)�}]w,t�����ɍ)��A2fgш�n0c1Ij��Y�K���Q���|B�<Z�j��+�T�`�ya��B��CB�
e�@55�%��/��/˖�K�PP�.O�tp놕�H�Ds���˩�.n��t����e��N�s�l�eQ�D{�q���R��q����)��%+fr,�{0�$�`�0��4< ��N��Mop�ڋG�����YI�2�n!|�-��s�Ֆ���r���55��Bó/u`�#A"3w�;F����� ����{;�0��Y%������j�2J�4jF~���^Ȍ:��A&��h�/�eS��P���t���\�d�!���7'|�`�!{�K����T,�c�!8I��DUe|З�Xil��*M�#��(ބ�7ӷ�xL-{�L��5�u�y!B�>�V���AYN�R��R˵�*���ڃV����-���hM��Ǚ�RR���K��yo<�;�CbRW�lV�-W(� ft�*@m�jp�:�r��*��~�wȞQ$ z}o_��(rDKv��������>��]@H��ۙ����K�������=&'c�V�2��zuPp|V�-;�G0CP�T���s�P��	��(�����D��E�����+M�7@d�긚c��[ـ�)!ⴏ?��sm9n=��/i8t7�?u�+���X~�{1�V4��|��Q��­�e�
X�䴎A��B��[�?N\��m��#q�-�=�F�Z��	�O�A^�U5/���2*k�$ORE�e���V ����+WJA;�G�Â$v�dl\�I0�t�Mr�Z�oK��+�[)�dj[��^5�"K����zL=�t�R(��ŰSĎ`�q��Y{���˒�W�Y�6�C�]� �0|�u�Ȕ9�(?z9&���[?�ї��.W�K�ȵp}����`�F�_˥qI���i�t|�clX&�@*��]O�U��}�˨�,��2�\�}2z4� m=�|�e![x[5���_V��c�j�̯CS@�\h�v�m�	�O���X��T."��}�Kq�>m�\2g��;b13'S��`=�H-OS�:�3��k�L0��T�SY�����ڼ
+rA4�����N�U��N�M���b��=�Fp-�T|XJF�꾚w�����C�_]i��oR;?����N�:�����'�U�w y@�R�w�N�$�@\lr]���7���/�����¤�����k������?�a����1D9�-�4��wT���_ww1}��M+)� ��X�E�h����Y�Kc�F�ݐ�ԣ�{�΃N�=�1���;Ŷ��}A0P�8���X����3�c�x=�̗}k�;QK��(;#�n__��Y).�÷|!�,�D��p�N��kz4��T�ej��T�(�؀m��7TiPƩH*u>, [���X�:��T�p y>�ʗ_�{Z��!)8mI9�r�G�5���T�=�k6�@M��8
�]LgX���W�a��^%r���j��r�#4���:=W�!��Dz��&r�
����4c��t':ue�K��M�J��^'�c?��Es�#��Ϳ5��e����2:��QKB"N�.�S���	����h�����an	IB�K��[�f7ێ�4�A�҃��@V�%���V�#^.�=o�'#!b�ẏ ����k��#��Hk2�z�}�Hi08���a>������I>�x�eX@R�K����sY�	��7s�e/1�V^s��M�
\��t��o���]5n����6��wՔ[E���z8��W�8����{��+}oS410�C|bA�C��x���#�tn��n���lX�Q�J���U���Q��)z!����D�r/4��-���C�ٽ�c���S�&n�N�(8�N�:�F*7:���`@W"ʃ��>�iOL��/�Kt���z���C~��R�_�>(��;̲�s��ԃ�Z� �QU	�+�$��c;eqj>C���Bn�G��7�m��:��F2a��������Х��#$d�Z��e{h�e�z�*4���0(tu���T�I��fʎ!�Se�K�H�7C���c�%z�p�Y5�%>v��|���1��ǰ��{�/^ᝈ��/����ęZz���@�w�_�b'���A��*�k|V�+�x���w�{Z�rғ��ɳ�)Ea�7����>�KV��^z�o�Z�c��Fqy��c�� ��Q��nd`��Bw8q��E��Kʹg×x��3 V������,w�(��i#�﮶Nh���{b&O^���L��ީҺR�K"wY.�S%������\YH�,CSt/d�iD�ɓ��X���Θ}�1_�p��3�����F�m?��2��x��wU��	쑋�1��Y?3�'`��%*"^�&}��#U{̨�޴��Lڌ)K��h+ͯ�C>x�E"[���G�#GQ�݁u/�Bv<
��:�~�,��V�nW�>��N� &m W��I�f�a�e-�������#��[���"�_��w{|�ǡ��5�#��uA��f�`�M���+i�"�x���X�]����x�B�=aG�ƺڇ��Sn����nT�E�$9$���"TBOZ�yE6A]Q8bL�%"��u��8��5��j�В{/�=k������+�v�'�g���kktH�)��~nN1���u�!��Ⱥ�� f��°��1D�suG���*�p�tAɫ�d�PM���ϛ��^�.��堰�gm���:o�`9�h%=nV�Ug!�&B�Q&�&�&LŃ3M�.2�۽���� �0�!�='�=C�s�R�!�;�'8Ԉ�.���j�9�SO�`۬:��lɀ���y�3�Fk�\O�ah���5%�5[y\]�w�Ӥ{Ӹ��&�����J�0�����B��:CWx���=��<�f���s_��n�/v7M+v݋�VT@ީ��-��ۓ/r�N�#��E9�w0�n�̠j66��c�A��SC�"���
��j�����q۶�0��pӈ���Z��a�7ȴ��F�����޵���ǈl���cK鑩�����%��[w��E� 0�16�a:<�M��?La�tQ�z��ɏ�K��º]ߟOd$*h�LC���ݔ��Z�e�=w�ي ��(���4ďs/lM�p���B�Pɝ9��|���q����	l���V�[�S�a�!�0;��^	�W?�1��1�1���D �`H�#y����5���ĺU���J�¼��G.b�����6��.��Eb�!uL¢\����0�EP��0��Kt!�-V�n'�Z�_6�.�O�7��!�E:�?���.�D%R���mdgD�BUط1��Py�L�G�J� ut���i�Y�*�5��'z�挺a�Di����+̺���g$�I=k�Ja�����ƌ��>����Z��aQ�Br����>A�p
h 6p?�sԲ��=�q�j�r�̜"<���k-�r*�%>���l��R/�A�%E_�`�DknՅf7�ͨ[�u�u<�#7%���mX����2��V(b�,y�,E\�
��F�@*C1�;)0BFC�KU��S���迲�nB'�ss6m3����rZ�p�;�C}҅��Q�xǶ�Ҍ�"���m���ETz�ev��V�b�޵�\��!��2$�&�ȕi�;�h�gaDJ������9l"Z4
�\�����z&��ߍH�b�8�ݐ����oh�=�B���}"���Pq}�cVs}<�(��fفF:י���^�:7�����x��k��1ƥ��c6�AL��-"TEg�����9� i�z/�{��/�*���h9q��D�{����>35V��Ng��|�jӫ�6��e���2�=��Ѯpd�cH; �[���lD$��e�+.G�9���E*}C^��ħ����v��p�M+�O,���`�-MQ��9�
oLbZ����1N�]�H�q�JnX�G��*�=�'1�%|Z\2��(0ɬ���5v.����
������M/�*�
�����I}���[�$�<�+��V9(�� 3"�0�t� �4�N_s�F���qD�\Y���h_]�_���HՉ^K���1�]�t�7�AL��}Gc�#f���U�`��`�W��6�q٘O�r�BꖩJ/�S^��e�7�V���nU���v���;�N�.	ToY#�� Sn9G�i��#��d���z��T|�1r��3&)�5�i�#M��0s����(<�{�FD��<d�m	{��vt�o�$U?�c<VӘ*�O-�A_�9�Nr��G���ڢw>Ǘ�r�me�(B{7G![n���h��������PP�� ��po��d��G�:s���T��/��v��U�[�R�3a��آ�	:�{s�j4!Jz&0M At�V�s�0�Kar�w����"[KE{a�C>�6$���.x�%I\�����:$ڬ�!/�����!ړ����/�Ŕ�C(C�(��.�3�N�*��)_��\�|q�d�}��t��v�0�PSWͰ=�]�&?�1sL��ص}s$Jh.�$ŏ��4z����6��-8�P��y'��L����y�Z�ټE�FE;쬀D���A�f�4U֜ݵY�"ޫ��
�	T�!�`���x�ϩ����Ҋ6�pozԯ�.7#�֨~�!�ڬ�0JSob�V9U>?.�W��B��ߘOFfb��/�Z8���)6�.��F�+���~L�s�,�f�t��Hg��`U��	�U��e�9��z5�%j������)�?�� ǅ|jX�}�c��۳s҈���%�E]"$�*��3�#�����'I�^C�?�N��7+���X����x]������5mT9J�����k�aY�s��I� �����j��M�e���� k\P�0\�]�y \ߧN B������	nJ��%�q!b[��6�r�K�&�v��E��-0[��m���<눐��� X��3�q���Sҏ��K�c���"p`���GH#:g���B��-U%P�R-�~�:���ڙ�������z8&�s�����(.uoJ/��R�M�B�+H�L7�OsYC.��7�xA�w��`�YṲ����th)�;Y�=�������\� �="�壄�a��
�N��/��`>����\%ʇcm��ZO�wd12o9t��_��o���QT������S�*�:<���e�n\
�aV+��SUZ�dV}%��0����Ꮱ�����s�6�:M2��~����l�sE�3��)�\�����b����C��N�ݛ�����$�rƏ�σN0Ԧ��D���n� Iˤ�֭Ņ�*���F���Kh׉E�>������=8'Gd�0c�v%�6���Pe��ś�+�R��,���T4WY�Cw�}̵�GQ`�%.�.g�R���4�x��?� �����_��lיD`b�d��*��b~�IUc�˝nIC��G\8U��w�7�S};D�Ac&<�n-#���������\�k���9A�	�T ګ
ONU񎝾��8�Ij�J� }����R� `z34qD?���\m���m���5$y��u����Ə^6C��5�ۃ|k�-r��n���xoz��G��Y�K��z9+�lǂuH���!ť��*�v��XI�k�t.��-ڌ�X�ck�j ����|��Մڏ����q������b�	�#�#z?O��]�Q�[.K޿��t��ϓ;�z0ڄ&�O��;���5�y��dj��Բ��`��L�Z!�\���{yA�y���f62�#������f|��KB���ʝ�/��//���pM�٧���p@/3ѧ�Ֆ�W�«��ń�\�Wp�3p��T�IG!9�kW��	8�]Z���.ɯg�&���"���O��,��{
Wĉ��������It�����6�����%��m�����=.�z`��U̮��4��[P����i�*m(>������..��=;с�/�h�5�t/l9φFD�()��y6W���0Qۤ�w�h�ih�]#ދ
�6���ej=G�nB���P��0v�3���y3}]~�[	�cN����L�W���e���3�0O�F�J�ou�DD�y#�x�]��_ݳ1B%{�߿=��maOM�_�лJe��U"���'��������G6�]��#A���%�BW�7s_��b����`��-pÚ��O���";@���& ��7E ��t�|�ӏ��]6L�0'I�/�%zhC�Y;r<�g�]�*0%�G�~ٟ���ar�
Y9�M�8��U�YW��	W�:�zq��	p#��k�a�s��Y�]�o*w3:�݊S����
�$9b��9<�Ж�ɣ���y�����\m�sf�>j�� 0KEPjiű��hG �s�x�gL�,��U�c�qH,�?����\�L;�i��u_��c��U%�g1���8���KlCz��j.�u��`& �\ ,[j�Y����Q�W�pk��Y^Ȃ��]���%w�䯒�AMxrIm�)�:c�a�~l�[�A��(#�H�;���l0�*�6�w.6Խ�l
	���Y���Q��٬釢tq)h�\׷ �09R7�6�}"
�a ��=�ϋ~/���g��3\�L"8�w���<d������g�b@��YT�S�H ��b1�J�A}��s���=9�x�4���!6:]�}`�v�N�3R	=o�Y���E��b+��Vb��ne��7.��7�l ��W��@���5v�����C�� ����#�g�jFȽpOF�?v�Lil� Fp�#��э�3���䧺�o��1�k,v'왘qI��Z�1ό�i���?���S�����~0�kۑ����۲fg2Ǵ���@�!�_à����&˙��9���N_�� �g�A�ꜱ��
�9��!�zYY>��P�١��$�c1�T��,�	;:���nbS/X˗����,�M�^px�������P�8:��ܬ�G�u�Wܙ=�V���%��|�|&�z�\�6�s��p�t}+ĢY*$<O��}���������Ʌn���b�چ��H�e�q>y̨$��P/ 㣲R���;�4C�Vt$�h�aJ1�|�:��D0�I�8,�5�
9���r�Jȯ�Q�([�Δ7?mY�Ϣ���Jkû~l��<�L���jS�Q�s���0���^;%�!�XNl��Mb.�W �`���~��>�H�����Bj�����j�_������l~'95e�N��	��mU��2����7$L�U(O~��d*��%��Bo(�ҡt�|<)!���l,���տF��Xa��f�®�7#���h�(���a��C�f
3��V'��x�z�����Gpb ��%�we?�Rû� NC-��j�Mg��Z	x�ohq�2 #���(�v�+�����
��=�-3�_���!��=�����?"�Y>Xz�v���L�˓�+?�`~7^U�NDu��?&�8�ۙ��Nk���'����~##hY/����<�`\�˛y��iYɫ!j)��a"l�BL�iT&АD�
���ad��H����d�[����]��ݬ��%K���7���0�̆d)���`ӟk%h��er5�
7��Ιa/Վ�v�{�f�9q	�CXz���/�t���[��{U&�(~n�$ەa3�63B
(6А����-o��1�:�Հt���(T����-�T����]VU������w��q��D/�q_ݙy~pJ��첎�$7a�B'D_��;<�]kQ���p(6�2��jq���=��������f:�b�C��`�o���("����'K�\�Mf\k�RM�/ж������}��� ��Sn�OR��r�8;;»m�]��r��x�@�-��%�%в@Er\�__!����nQ�ꁔ:Q����� r �35 G�L�w~,�q���o��)l1�()x��c#S�6\��If�|6�Ο���	�~�a�e9�a#��%!M[��,&F�z�OE�N�2��n�c��b��|�hz����`U�-��E~�qr��a�,�:-�q��ɝEO���$Ǖ~x����>���N�R5���~T�INj��t�lQ�n����}�T,U���r0�m�E�l3���,�� �m��Br:'B!E�I�r��l4�g�:ʒ_]8�~�/jԳ��J\ɞj�_r_ԭA�vYj����1[�<���T���x�s|>�F~,��q}��A�w'�o���]V�:�6ﴗ�;uG>Wڴ�LeC�����-'dz1�5֑e�i���8&}f]r�.rL��)�lJ��a|�G"$B�s3��M|��{)I��H)dͯ.��/������/�e����ͣ����(8;;G�1��%���*m0�����:*@��˰M!k�z��]!r����i������ )�J�b` �T��e�}ù��<�S�Ӄˀ&0 P���U��2�<�(�ύOV�п���:�ˮ�0�8hp�,~�"s�w��[W�3t�'��]���^��{P9�$?m3�{��kv����o"Y��	�!w"a�xe�'�"ω`Ԥi�8@�VU7�5O��%�;W�4�B�������$Iw���u���u�>Fv��D�¹�08R}�4�dBU��M,��u\��I �[�Q�w�O?��������Y�^[�1��`�Z&ɇ\��ߖ��z�n8vD��U铓}�u��/9O�(�Pw�V^#��Jl1�T=,}0�<��d=�o��bKB�,l_iE�2�)��4�1�ުShdZR݈p������Y�M^W*�ìЬ����_F�� r�R�UL�.�uK���+�������&��$j|���S	]����;Y<߼3������&�������0�t��Bx��,9��=�����Pژ�A��wX�=��'��7����3k@�����4]���:���dF������4ŋ�'����������2Hl����/<�+%��V�'A9�G	���ɽ�����"�ʾ�K�8O �։�f�y��f����7����^�2�+��
�h�1��x�ô����ĕay����Z�:EQ��\�hc잒d��R���f̿���L��~6Ϻ�F��vc���{��D�a�&[��(n�l����봥�����T&��J�a{Ӳ򵓰Ǩ�1}7{Kʂ�Ƃ"�k_��ך�$XA� �U��]�
Qm�Yo�R"�a�ś٬qmK�Zz^�	��5X�q"�z��F gZ�\&�<��V��9����~��Bd�ة�*k)do.��g�k���f_���Oj��xS��Ц�&g'�ekj|C����]
4*�Eoi�S�p�L��P������݉;W��"��h�����,�HF��x�z�)I��阕���xWc�C6FZ��������賋���ύm����S�
�2��;^X��s��͑��,�����J ��
�V������)��$�o��������(���� _Ϳ�$�p��i�!#��qi�Q���R�,���C �>M��D�S�U͂�W1mn �oi,�H�Z�Gq�O����=��q�[K��.+ح��2,pȍۦ�SWh�J��2K�bs�È�]��]E~SSv<RM�浑��
��j4N�?�k�'��$�w.�\�I_]��k��sgȣIw��>P`T�_ϝ�?m��p�ۄf��ъC�5B�섺�pؿ�~s�����Rxz�������t�Z�:- `�%�[�oN����gB�P��0�������^Ǘ��PBL���N2ہ�8�z6��Jm�vCH�ĩ"��{ܹ��Q�NP�R�j��J*�l?Fq[� �����Ľ��88���Y��z�+�9��Yx�!춏 �wj��P����	]�TPl�1����ٙ�%�H>�t��k����rY��9�&7��}�wӧY���}fa��6��*h(,�gVgdfo���?�͢P���	"�"B�2l;�+�SeP�f����y^���h����z�������d�47��r���4}W�Ypz!AA����*׼u 
&0�zDػ��4��p�ʀ�"�eǽH����7�;&-���K�����t[������@��.��bC��Ҝ��jWԕ�JIE��:=��T� %S�����_l-�H35wL�/׻��i�f����<S�����C��b
�@�rO����/�����J�u��M|Pl�~�SIœՕ��>�MI/��j�%�x����,^g��ܞ�{�.�vw{��=O��&��>\��ky۩?-�-�uJ��lL�5l�䥡����j�wз8sC�۞sēv ���?�*3�Tw2a�t5�O���$�OпHDX�39\9^I�N9��d;�n��V�;�ꩢ[��OI�s��#z��d��J'�P����+N }l�*�u��F�La8+:��RޔyA萾*Q�fK#�5�%!9�\�1��<�!1�P)GV��*+�φ�x��'Czg)�q?��N�����i���ij.�ǿ�/"��@0#�<�u�r�7@���B�,��w���t��|�����ϑ^�^��5&�_�0�Fs��+��-=�f�s��&8�D�҈TC�T	�`�Ǉ��M�ӊ�Q�e�ۯ���Dť)T �MH���cd�_�%R	han�g���N�K'�Cqݗп���l��Վ�/�0=C�f���W��m�aP����~!w�ZJ7��68�G���Kep��AK͕G�l E� �����@�����q�l��ƫš%�8mHB�_��D��e���o��ڙ	)VzOH�������K���#E��V����-��k��j�D��wi7Y�x���?����cp,�`�f �Y7���$��Ex�LO�xV_�ԁ�(g�
���	���D~[�j/�Y�
�V�x��KEϕ������������ ��O���E�	'M��cӷ��~�b�{Yd��Gbx�I�d	N����E��y��BK6��ӒI�7��R�=���x���@/DD���r�YNV�\��Y��-ǣ��oNxp��	[�� yI}$�wv4/�c�:�e���k\���� �N4Z,�PHz-��[�	;D�(�EO;��[h��]��z�=^�sS��J�e:
��v��3Ub��JU$���`p�p���,9%v���Y���댣yCΟ \��)Y�ޙ���8���:�X��6SF>��î���E�j���ͦ*f�e�/Mw�ϣ�������QK�C�BP2Z�o���m�,E+��vh��^�����,���s��3�{�V ��̍P�cd�/:���Mz���1S�����Ƥz�b��f����������[
d�IvuN:�{nv ����nf����7�vc�x����7O�z�n������Y2%3�O���TO�-c5B"Ǥ���J(}QW9�VX���'���m�y���}��1��*�|6vs�O��ܒP�O04���Z��p�6�ؤ���x]ȴ�M��R���|t���	�K�a��U��#2�Xܚ{��5��7"}p���k*��R�틱�	J�D��8�b�XֲA�9�s�7��&JXۖ9Sj`<DD@�/��4�v9h�<
|s�3~�Rp�q,�^��4f�_���s��U�¸4E7A����b^�04(�E�!�aO!�NHH<o?ͳ��}�-�����T�s9u W �)�I�ڶ��au��F�����(.��SD�� k��]�3�j�����"�j\j0�������2��x�](c�ydZ]�Fm�6h���ZM0,<Ag�}�����Dnq� R��;�y�8��"����K�+��M �H���z)`��C���J���/����d�\$gYF\�Q�{�'o
0��X#��/�D��/�L�,�c��Ouz�G~�"^	
�rq�S�@���3��S��1+����j�z��$��9Ӷ*�6�'c&�zl��[���~Z(Sqp�7-y���k�n1���ƤE{�,��#�C��G���22��߰0O?գ����!�؃��*	�� )��(l~�6Ht�&��r����j�툞kG-xF��X`V�����X��ǎ��M�8>�V�G�v]˳��EM��i!�q��&;�kҠ�)����Z��QV��ѓ_���$3|�(Y���M�4�_x�+�%vu=�N�!�r��[A��̸�EU9FQ��X�uC\��\��aC�x��9}ѻ�����
˟��O{Brnjm�Gq�>�=e���YřB�<W�z���vW���{A��6њ�kt؀�i�܃��h��c��܉3�n�S�c���ć"�Sc��S�o�٢�g��^?/�a	kӰ+�tވ��A/�XF.�ܖ�g���Ķ")H�4��f���:����q1��(F�Z��?��#^�r��]X()��FD�7�48>�p뭮ȞQ���D�W1��g��b#q"�y٦w�30��Wat�&���<��f7𐊉����!H\��e�n1Ls�s�Y�h�ӏF*�,d$#��� Gg�#W2��+�NM�5T�qC�����;�-@,K���^����v�ۦ���ݴ]'��4�� ���+�O:�|�����_��綦���(�
0��6���W��% ��@�-�"���@�SJ����A�Yx�f�q��B]�x��x��0�cwU~�P�b���-�8m/!��M}��#�D��Ǵ�'�M�=Xe��%7)��ǉ��T�"�<�����}�oMLx7�TqsV�j�:�N5�R��j�B��_=�koU�u���ڶ]IXx��q�nz�xI���-�aJG��Lj������e�¥�
 5o�1�Q��B帎z��w���~`�Ӳ�<�	ͨN=eoK�"�!B����)F0�E�Z$Q���|���`H/�~|�u{G�-��=�k�|���I��fk��L���_�rm&�UWY����R�*�T]��؄ϰTO���_��Qŵm�����	�!����4��;q��Y��_�*�@��������*`����c:�t�ɣ���սT�P�?J�sӲj��,����ړI5��zB����n��E�Qq�"-��Y�n��؊Zz����֠I}��G���_*^����M�*�n�Pj�&=o���qkv0:q�
	��-�~�=�8j\a3�M�Q&�/Tb�AEoͽt�rl6'Q^�y�dB�ﰰy`�c6�:h��� p����b�S�t��)]
�J�x7��97}�Ϯ��,�;�C�z������<��$��Ba�����I��G,K~�l�
@ca�a�Q��τ�ط��5�Ǯ���sW`,��Z �ͩ���q�=2� 1W��a�p�����&���R�LD,�g�H�-^�����h��O%��	q˖�9�E�gf��؛��̠�ٞieZ
��0��dC���n�g���9���E�g��r'�Z[�����g#�<���՛p�t��Z�`߰s�w������s�&{7�u�^�!Q��>��̈́aX0F�#-��<�(8)�va-ĕ�R�M��r��u��),5��ocwg�4�����L*��j�5�;�:6��V���;��*�=�<�� '��ӛ�M_�Eث�)�s��h�_����#B��p�.݇:s�D{J�$�-� ��� �Q��y�u5`=�0�h�������K�p��c��<?��pS(Ѭ��# �M�-n�\{*��̇��;,˪T\XޝΣ4��G��H*F��t�.�\O$$qꪖ��5�	뚗�e�/(��V�!(Q�����R	��߯�rէO�摥w/_ěZ ;��c�`���'yhQ}�Y�l�2���9����b���w��۬�%BR*(������;��_#�^HxAO�����nu��f�uq�g9K*6�Xe��"��!l�:l{��MXG��K����Pe����a%�n������,4�-$�/��a��d2�i�u���㒞XҤ-,��>}������9^��rz`�6�2I|�Q��teK����|;�f-V����T�r�7:��j�@��X��W����s�J�D�3�9�q�}i�}�̪�02"��P��esp?��ڻ�b� �q�,<�ð�E�v�ɩ4�+��c��SK6�|G���/`���C�� ʣ��4�(�&6%�����g���t��>(��O>[��n���#��@��4�Sy�U��5���M���|$V�џ�yb�"�GE�u4ۖ�n����i0�2Dq�g�:�%AW��Be�X]�)u&�2]m�E�<����/RM�")�hB&���M����g��j���U x�Вȹf{{���=X�1S����c䅽)vZ�<2׽h��>�b
�2>F�oa�s��>Ӧj��t��z�Eή��Ŭ­��I*4�'QB�NIε%����P>�;K��y��� =\� 1�^y���0.����o�_�@�� v��)G/�F��]����݌�'�S��xѷ�v�pXr9����RBj��W����۫�O����H�N���Ao]��#�Ƚ�	O*_y�_0�Jov�\�������u�l��#�-�;��ޅ�fϿ�0�!����3����]�xr�!�J�� ӵ�{�����à>�+���%!�{�0�i���f2��L�:;�b�]�1����{�}	�>$j�}Oa%��m��������l<��v��)��=
���	S3��pi��[�?8�'��0����P�4ѐ�n��B3����{ �X�8R��������	\9��\{Z�ԢL��n3m"���s��Ŷ.���\V��'ip0������W^;'<��V�vrW!]��G�1�)$�?���g�F啴E��!��g��`p����!A]��,�[t���iM�cj���%���Õ��'(!s]i`n���%�����TU�K8/c�J�`�kcPe�L�)�a�P,���n>,�Vd���4�����3��Oq����X��ƀs0��N�baw�xذ����B��]�2� �
d���enKE�+�CG�lB��������w�)�%�M蛖 �jg�	3�L�ߚX��rw1:�k�.�(�^ѼH� �hf �B�ּ�;�3�V�H�^�Tf���7ܚ����!�뽑��IՆ����eFt�����ɶ1U�����c���lʔ�e� .���x�<"���̒fY�&Db��fG�{ɽ�#�+���{�>Ʒ#��f��E���BRdD�`��Y���d�Ȧ��p!�XZ�`H����@/!�?�^)&[��z� �<��boa=������"�cg&�x;��7� �]�����D�Eo��2��L��UJ7�IZ��I�q��W9�4�7�=5�0�f�$�*k̿�N@���y�о��O8h�>:�#?l@��5�w�QX�s���!�i�Qr9_�ϟ" ���Y��	�y���S[�#�6���
�a����
8��K�-CkJ��kW�� �6���}�4!�f5��r1z��8�aq�,���%�@.���[*6���}�z���1c����¢Āp��d��o���|�(�bj�7�/��Ұ�΢�r�5����PR��[U"�8K���/a��IM�[�g�h�N����/�&���e0g)���Y�޲���_��"ս]���_�k� iI���qɥk�~y��2&�;�T���:����ξL�{
B|y��a�����$�~�u�Pf'E�fd3#���l��0%����O�h�w��]��7���x�JD�k�Z� �J�8��v�b���c�[,as-�8�:��yo䩚0&EB� -	���C�M܈��x�U�߽����	����.T�q�P��L�{&�g�t� f����z/
��%R 8M��)��EZ�Ͳw�
}�W����s�z�����Y/ĬW�Z��^�;8��Es"{�i3q�ƕ[��
���Q�2ie�e�L�����U��?r.�߄;`k	��8Y�ד/�Hsc�n��u�nf_S�`��.�E6k˓����ḲX��rG{h�Z��鮣\�˹���	Q�ן�|Ln4V�~sn}d�)�c�R̥+΂K�ޖW��B���)G$jm�V�Dsd��e��6AVS���J�UdQ��Ņ�6�+0���\�9I6�ـ�EI�ï)�=���>���n���t_�����7��w�Q�� H�y�,��Nu�5|��ֲ�����.JV �E�]��5��ꢎ ��&���մ��i3�@?x�_�B�,�z�	�?ԝ{�B��]�H#A��Y��}4'�d���"�UTu���0a�kB�������u�kk�P��)�1��C�Yuv�㥲L�!-�x��wޝ -�jd��l���R�qL(��o���l�
����;)��s8�cxB�� gT����]_ђ�<Y򠃜_��o��soPȈVb1٭�Y��6�M������C/�M~�O䔛fh���f����+M�v/N
�p|N�~ɞ�}�Ynmو������
y���0A\G"��r��_�U� �yp�!���iL��R��IH�̪4���=�ꨶw���Wbk�{����{2M��'*�dW�m����WŨ3 ,Ɲ.�r�dT�򖡐U�H���-<�5�թ�*��Kh0�_K�[xp��w0yXg4��p��)�a�N#㓓ցb���m<b[�#!�~��F�5�3���l���/�9��xJ]�{�󄕳����!��O�7�Vg���!p]lV���|��*i�Y.FI�� �ܢi��˞����:P;�n�+��h���y�бt��PN�k�Q5w��Չ�~�Q�xK�^f���շ f�S*�h�~:{6���������5�n&L��m��:�����_>Y6�#J �6��<��9P~�s��"�v\ʃ�V�1[�Y8��d����{z���$]���	>�?���_�T��A�up�}l5�e��m�����+������*n�nķ���.p����*����ʹ����o$���S�s9���"��3}�f0���U �`���S�u��4�)�����j�/*��K�Y���Y�p��� 9���d�#���<��0	�ɟ{Z�*�܄ ��vo��C4هtgU�ȥ;H�Z��K�rWQ"	]E�n	�����"4a����i��$�Q��w�߃c�c�ڦd�^2��.�Θ3�#@0�'i-�
�~��?Ќ�b_��7��8�¿��s|-�T��B���}@��O�ӧ癀����ʛ����!�����Ux���i��ô	<�!̖z��y	�7��y�Y�m�(�2�,+v|~�}Z�4\n� P�|)��2Ʈ�= �s������Wİ��܎���e�)��9HHY桘HiolȣNS״��	�I ���WYT�ފU�	7����#�s�ޏp�����d���Y�cʃ �B�o��ˏ��lA�wpD�t@c�2^^S�d2w�pD	`��Oӑ�>���Gm�vE��>E��xrR`�m�#�dO-ሱLlѳe-���2{��@j�π�UY��T�Fz�@w?��O��pY�w)i�n���
. �<'�3S�����g?���l_C�::no��n�;�\EF	�﵈[~��������e+����8 o�.�y0��4I��U9�4�p����9E�Y;d���'����cg�p���ǹ�k�C��U8�09엽V��Z� ���?VyH�J����y����]����1�t}S9��NPw��\�8�
�1� _��	���*1��>*���w��q�D2�.�#�$4+b	�_���N1i^�Nu/]M�� �Pt��^��y�i����Y�b���zE�n��O�o̈́q���.o8�S=?���4�'�j������VR?�����@�k[ݶQ�l3W)�^�K���<H�=;AV�{��ėQ�tj�Q��$ZM(\#'������6F�<�=�&��zr:�}9.ē�Ӂb�{�x\R��Er��ڀ�f��r��z�!05O����$�bF'�5������\��xa\�h�H%���� �ZQE����d��������+�z�s4n���ҙXb��/W�W�Bҗ��ק�Zb<�������И�.7iF#ܚ7}����EL�B2Wʘ?��J����V^���	}�kv"��%���}Њx�(������L�MT.h����l�%��I:S��U����o����Z�(������C#��.���ܔ�Z��B�iz����h;�õ_o�g5�q.�S7��fP `mw����)5�0xt�/c�?�(Y��D2�v�Ɲ�A�`�F��G]�0�B�<��pi�=� �\�G�~��W�>����R�T �!"Cq���b�����ʮ��D�u�FҐ�b��4�ύ�5���.�q�Q#�5޿`�I�D����%@5��Xi�/��8�w�խQѾM؎���!Ó��}��H٭^��I�
�g���%5��pDy��^Az�xj=��d��@b����ۥ'����k�x���~����l4�~��#R�Tn��w���p�dˎ� Jn蟄#1��w?��Ѡ��mC� L9.��9nȍ5�ֽ�:~k�!{P�4KҠ�Nδ��K*qυ**���g5�RgY{�p8V���7�MA��2����3B%=`�>��V�G�¥�<�X����s�R�_T��b��8CnW�:6��:�|�Q�mn�媑��k<L@��ȣ2c#�����z�{{. �A(m5�<h)�{���v��wK�?C�G���.��RAͺ�jq?[��s�F���,9y��`0�^��.%��.lA��O��Z2V�e��SS��y!�*��58yDAw�J�yf�DY�p��6�3ҹnb������h�ũ2�"_y1I{�����vޙ����*��✈��I�C��ҙL_�Q����s5�'ҡ���7Xx��`�7����6���R`�8R�� �e��zz�wz)wY,	u1�F~٦�94+��ߜa1��[)۞& %���f�"r�y�16�xl�����X�E�|��'=u�SS���u,Q�d�g����7ݒY�s����o�o��y�qx�R���[���*c���9�Mץ�K�Y���O�%�3�\�H�r��* �&��4��{Ёz�X�ş��*��Ƀ9G\q���6q-p�C����rO�Tp���&��877ࣦ����@2��`�7o��C�B�Ç��МhQ_�L�+c�g��.��+=�W�f۝-���<�1R^�� Rݰ����J&,=	G��n
Q�Ί4	��_D:���C���!��zx|� mS1N'I�|i�ވZ���=�d���6'�K`��no�s���t�'�<eE8`�c�c�P,[�����]G�L?�
�ЂQ(P�䕒����?_/G���/�5��W�$|!�>�ӊY����	B�c2f�C$ׂ�W���n~�.�{�bw�餛��"�y �FƜzZs�u�@]�=>X�{��2S��L9Ī����'��F1�Q��dA�i�fc�C�;i��R�?F 0�aD��BK�K��s8ֳl�w���=��%�������/�c����9&��6��j�Q��D��Z�ӭ�h���2lf����p�.��j��Z��]@/3ޫA� ���7�π Ln�Q��s�U%�����j����x�!�����|bѾ쩮8���������JX
H@�0m����cB�c��|i�\4�p/Izz�����d/gdA�dK����V�	���'�8��|�h�]�R�1�����vAih���y@���1d����C	�d̋�9'�}�Ks�7� 8	dH#��k��.��ᧅ�.Q��������/��75ωF�6���Q�j{�!��4y-�%z��Kߚ��bĩj�t��W6i|�K�kU�%eEjp/Z�6��Q!:�r�鍻�EPefZr�u3s��3�P��5�ԍ�5��o��Tr�s��/�Ca�q��l�*f�prN8��S�\�z�ׂ|:��A��;Ko'�f\� 	19AjI�i��MsR��^G�eq���<-��d�I6��5i��Vþ�d\�N�dw�3v�Ǘ�_����*��w<-�3<��jn&�3ն��+T��Ь����'�·�ȑ����p��^ȟ񽋖1����g^�3)�{���/���M ��9+E�����ى���2�B��h���\��[�`���R�_�r�^U.�0�s���*�~@�a�,j����;zuO�誃�@�(�7܏���h��6XD���k�n�u�B� ������%�i���XZ�[{&�To�,W'�y[�7�4H������[e�zy�hO6Y��B�����Aua0���a�-3��Qb{)0 ��n�1�7��l8Fl���Z!b��'3��!� !J�2�#	\j.WF��j~���4��C���V�n�p[�p�ԕ)�V��Gd\g�\TEȂ�0��c�/���3�׀����@;�\{oܽEډUq�]L�N�*&;����z�mF�yw\�g�tz�>c�c!�Xj#פ5�mN^R:��ɥ��#�(�����=J�$�lʶ��;o��Ŧf����^[�6Ã�}Iq�O`�C�ݪ�aV�b�J�iN5����~מ��K�xj�,-8��t��/�X�������:<S��В�ZNQwA�"��/��CdQL�rDr>��7�mV��w�A�ُ��y�8�`�9�y?v��ZmѢu���gi��K�:P�u��T'��7�C�Y8�% ����4@��o��<+A�����ϓ2�0Z�_��9��=��HO au.Gxc܁W�[;0���Rȭ�C⾸*��cs(O괹�W���N�l�Y%��Ƈ�H��Z.4�T�ڨ��x!�� �j�c`�~�� ��-�,�%p.9���mwA�/�%om���u!��)W�
�������"��~ߜ:�Og�MX�cѤ������+�]�2�L/��#�1��,?��<ޝ~�t����{������)t���rN��cK�j��Z)����VQL'�wa�I������ �A��0���za��`��*+/��z���5;�1C� �� ���W�M��?��G�`�ʌKk׉Ҩd��O�Auw��)�Ue�wV->+�Nʮd@�4&PV[���2�:�7���L�0�~���lm�*ļ��
'�
vV�B�D+��S-\D�Rrd
��<���5�ɼ��!�z۾J���^�ͣ�G�@*e�T�TEj��D�-T�d	�?�E^�"l�*�7��|yO;���>���ߵ���~��7��y��j&��X!n���g���"��Qh�`��h�il����y�����-@)���0����`�
������y�-�?�j:X_��d�D�
+��AoN��#َC�g\��9�}�zDJ;py��p��7^�s_tyⴏ�N�o��_��8Y�W�w�eϬ��vy�
oo�J)�Q���h���������3��}4tSEo����N���ӕp��)T��V ��%)�՞t-����=6/�rB?��X:˗)G�s�'�H�/�<羰����L��n0lXy�[j��́�� �0V�:�o�R�]	U/~I�X��Ga�e��W�z���^�Ч�_V�6��N��#۰0ԃ�I� �a��oD�������G.�}ϖ�����ƻ
�sҔ|�+sT��aZ JkR ���&>D��"%�V0�AL��5q4��-�e-*����:��f1��ߣ�cB�0ڜSc'�n5����Q?N�k��h��QL������G���� ,H�G�S�9솩�P3�d�K������?>�#fa@��edL���]\�����O��^c]���_\I�؜~�ٮ߮T�'����A��!�}z�����Ј��k5˦w�B7`��\�jr5��:I��Oj�	�B�)�G�(Y���־��N9���%r�;��¿~�ˇ��	@���3skΛ��g����n�!>G)#"2���W�׶�ڝ�+hs�c���^I���NoΖ�yHp���c �
$l:�J����KZ�{�n0�B�Q� �/��u͆D	%����Wk�0٥��5o{-�����H �2��_�=:��7���)�d��3Ɗ���3�"�^`�\Ǳ�W���ҧSUM�	�x��(���f�Ш( 6�E>���p٬]�B
*����7���w�CÝ�̛�&󋅿>���E��CD#:6��$�RzEs�|�')/�[	D�S+�v��{�< ZD���"Y���-�z��L"��#�^gA����6C� T�O�-x�V,*%��o̘�S�T��}.���I#��o~i���r�-A���2������)y��@~�����-ǜ�{w!_eY�Q�m�1?�uweݜ��W����<�r���a�Ȉ>��������N㏇吇 r5�:��f�̵r`�o��qd^?�o���ǤI�m����}`�	��8n�>��o�d�m8���MT�zG+v�����謑35U�̀ĉ�w�����au?���%�4�7��/�S[�P��2Z�!Wʜ�gU�kB����:�U��;=����y�6P��ポ���*��V�k�?�t�( �a��m���z���Z	PƆ|cY+'?�ڲ�!�� ������d��ϸ��2���@@�.(�㽙�3��{�L��[����_o����w��>��($Ba����+z�V��aH�o���N��l�x�u4'�z����ݍ��������`�>҄k�pO�`�S��o�\(Oiʩ#>>�6p��������Q�wx��7$�L�1����B���k."��*)("��ة�Ж��B�ئ�p�ZL�r�R7����5�\=r�LI�9�~�C5+������W��쮒�Lm�L5���m�S�P�Z�M/��<И�6(5x�uHR:�����%_SkGw�n�I,K�`���!�t��5O�"�5\8�@!�-��w�b$/t��,>�nĭ��QC��)#z R�c!!nU��)ր�|7�I���d]uz�ۺ��� ȴv�����y�(�8���#����QΙI���GΚ�c_��cM݊��i�ٝ�+K=�;}�|C)A^y�wz�E��2�����-Xqo{����0�u�P�J�;W�i���ؒ�Y�Z` �S[ K55�,����d�*�((�p1��6G5M�	�OO�[��7����R��x�W�P��/�!�/�}}�.Ұ���8X'Z�=[�\��͔ȂK�MH�v���{�|{�y�����	m,��;����,�����J��o(�R�IdD}��Ϙ��ߍ6 A���7�B�Y��6Z��'�T��b�������W-�l7�/6y�	%}���]g�;�o#���nW�P����K���ԣ��v�rL�\�.W�/[�y捈d�m��3�9��az�P\eH�#ք�����c����+:�7�m����9T���1���gN���1[�tL+�b�OAJ𮷾��iG�S�I=��Bʗv��s��1|�!�ڣ>qm��2�l�8��緙�V{HW~),ދ���x:S1!�r��akz5O��5E�`$��drL3j��aX@��_US2=!l�ȁV@naJ4Kʀ�
���k��a���KE�v��P������#��C���sڋ
h��NQO@K�VE�럯Uf��L�r�E������um�1��A��t^���K�&pJou��y�Q�ηL&�e�#��yϘ��6�F Ml=���ࣕo�^yA���2��p�F=��\)�2��>L*��&K��W�e^�t�P�J���R�LX�E�H�\�\J�w-}�� }Wޝ�ˌ�{�FR%�1k2K�x�u+����GI�|Tt!�9$��汘��MHA�}pj�����Y�qDAz ��r�FZ��)�WT3�8+��)��+�� �w�TLs�����o�&��z�1���&QA�=��3�)���F���?}�Iר*vTt"΄��1�QwT�L��cc��0�r{�ĭl�x��R��ޮ[�ģA�S;A��@)�䜥z�+�l����h��;�5ᘘ��_J:�;��b�������@�^�w��x�[\�F)@Z��sN��1�ڑU�'Y*^��'�d�o���]ʼ�MH�e,F�s,��`�w&\�r���e����1cx�w[�30��cx����Q����1����²Rq��'��Ȓo$Bf���uذiQ0
�&aḽQg���m�cd�/Ӡ��]��Ҍ����u�ͱ���<n��D*���|�rֆ2�R��<�G�@I��t�t����<�-�@�?¹7�&����u���H��8�j���-���a�6[�c�rD��冴�fm^_� �Z��u�zۭ�;��8@��I�F��ˮYTؤ�_���Pq˩�{S*`3_9�2kR�Ē(�\���v��hҀ�
��WQ_�9��e��9��v����'�]Lu�4��O���Auz'��7��;2K��AU�M������+*M3�1�9��k��%�2h�em�ߋ�äP�"�1�ùj.�~b�9���#K�B9˔��%�fxİبV�gR�`�\0|#r@;�t/d
�1��d����I��KhA�e{J��GFC�{�r4�bL��QC�i8�%��甜N���j����ֵ���i;���� I>����kVj6��;���n3�y6o�p�[����PDٛ������F��/6W��b9[�oc�4H�.K�lT�Y�2��7@����\���֤�kxWb�t)&{�j���d�߳iX�V�"0�K[���F(_~>o�CZL:
���x��c*ok��N����q���̔e��lc�I��G����н4X���(��.�A��̩�D/3���x���M�f2�uޘ�̢?#$��R���@�,�P��)������j&(��ˇD�s��W�P�H8�a��"����a�v&��^5�:Ɨ���n����1,5Y��<�iF��5�G �P�qeO7�w[�~�rmL�Lt/�#?�	���������?�zL�5���� 5U��. ����Z��ʵ�;�����GeBGu��;�K��������}3FD]�Wf����1;�<I��LB�C�\I�ȋ�d)lU��JU�U�;Z;Σ)�3YN'�`���Q}���ވ�>��!縪�J��'[Xҵ�V�N�.�N����٭_%��<�vJG�Eh�����߳�?�}�����w��u��lĢf�Ē�q�f�徤�GD�6�i�L���B�4~�+@�b�;G�O��׆��w֜��Ͼ��h7�P��e���}�E�]�gz/�^�gƏ����[u�z��h�j�z7'#�X�����sϑȺ�q4�
���hq�P�gg�B��`�1�P`J�s0��Cy1P��\>�yV�s��h��*��#k�B����T�,q��l����!����� ?��o�s�ڍQ:���;\��N{�(�+Tn�����1��N��c[)�4M��&�a�<����&!0��듺ʮ�-�ӯz���Ґ1��c��a۾�[�;)~�;� ���'�Z�r�	�0�p�;�؍�YcA�ą���9, j%�L�AF�xk��]��Nv��a�♷�#�lC�����;��VWCG52���YER�g�����A(�n8 @���B��R��w�9;?��#;����2AY��;�F�%f�c�n��f#y��N��}��
!>�ѐ�����r청�v���ܟ@$"��5~n�\[���حp|��S-�U�v���W�kJ���PK��KP�s��'�`?^�"��B3�*�h�^avH�6h�ސ�>�j��.#�.��y��~K\g�1E&��t|�Y��De?w���o��R�|�]��-!�o(n�oN�4^�X^J�I�	�t}�h0�q�$���� '���2��� \�j��R�T,V�+�ݟ���V��γ�P�JD���U��ֹ�)�(�ڹ�LhI@���r����ȅ�;�����#�	��:�sS�,
���b7F[M�{���]e�!g��	��tt,�.	�m�κ?Q�,��]+�s>p��6w "����"=�����ō����M~��C�y:�A��jŝY���\[T�:OVp�����s���&����K��RA(e'3ݯ(��n��!O�1=����Ջ>�	#��M;��_�a���-�)�Zz���G4�m�	���TME���e-ЦZ߭rm���V������̜"�X� $66O��5?ߐ�!M�F݅&a�\��w�#WѹXpb���1�JLuJ
�)2��fKx%90ڌ�ei�ع3��3m�R�(b�!��S��?�Xr����r��[��v3�����	���9�o�:��T��̽iW�T/������?�l��zc����}���!D���Q��KZ��B�ȗ5
Gz�a|�,Y�LHB�z��rh]��<��e�@�!����&^�2���2����?�Cy����(t/d}?�/�jA��.i�^0���{���C�R]GH�3��wM d���	�a�B6.���� 2�s=<ʅ;r��9w�+z��J(�W�$rM��&�Lq��*N&eZh�*�q8�PT���	*ɾ��"���4Id�	��B$��u��]>�)�!V�\,̚�J�Z�ת@���s�ݽY����fu��g Ɣ�5�G9��T����1�vg��ٰ��|�ϫ��9�@���ogM*d�E�s>B>��x���r/�?���k]�ޛ���VO��NK�Nf'W?)�~v�NR�/4����8C����]��Jn��KA8��-w��^���.K�IH�fǑ��?���{��8��TZ������5e�Yεm�䣢�U�#��1(���i���\�>��(�����U6�{����2^#) c��6�{�5�
'�\>���m�����1q']b��tc���[i�D��yZ6�z9 Z�S��K�j��Ͳ�9��L��mӐ}Cv96�k��y*.B�<Us�oŠsB_����׉�|z�Zq	L��[�|��}f���4.���Ѷ�۷�x迲?�X'��D�[���"�uQ�w�f�F�5��"dQ�ʉ9�sm�K��8�|=we�|&�dM���g ��vĞ�.�-�&�G�^�KA�k�"�<iP�_MG&�O�0���>�%���cO��b�6b�&�J���o��h�����KT���<�|G���*"������>:/f�9�9��U�:?���M4C�
�[8Q�ג��æ�9]hE�
�j�]@:uGe#�nA\��ص#A(?m��K���]�9G�P;M}v��+8����{f/�����i���ON\lY��s�O�< `�Q�<�u�e8d8pV�,r�`�w�km�l�G�ο���.���{�bx�an�5_߮O����<`W���R�h^�S����ż�2" 7�ҽ���~4qݿ{�4yo��[���m�te/|��B��T�Vt��]`UVn*Y�ύ�V��f�W�R]���l;_v��d8�L#^�p;Ӗ��֙)�ߤ�Q$�=�p����� ؔiY��5���������`\�Ñu�f���_�k���c�2���K��,!%�N�-��<O�,�J�V���>`�*���5~w(gV��������!� 8����H����ݑ����XV�ȕ"� 1�2#��9��2��Ֆ�,*d�_&�����Z�w� Um�7�pYՄ�)��2���a>!ف�$TlhQu
�c�2�N��t�z T+6
5,w���pPe��T�A�}h$y�j�~���#�#��6i�6W�*�a�&ᅹ"��(����HjmJ1�-n���7�G/޽�T�'"Mí���m�5�BZT���K��i�7U��h�"!�Ͻ�G���C�z�-IZ`d)7sk=_��b�@3^��k����Cv�e��7�s���*Ԏ�/1�t&��
�ѵw�rcm�ʥ_���^����S�饘�O���MViA�)~ܤM����<w�B�G ��yxX����b+�r��DwJ~A/����[d �k4��t�{�e���Z�xP�;��qX��,��'E��]�:{�=�*_[�R�(�J�m�{����"a���>g��K=߷^Ŋ�1&��B@�U����H	\y�^�|!	��2��%Hq6�G����^}/��mn�ݚ�9F�1�$6��Ұv�&���X#e7�ADo30����xk߮;��	�/:���&P��?p�� ��4���KZ`H5dID�u�'�Æ��&�'@E]�SW��x9�	l>�!ʲ�G�
d �˓MFK-��moIqaF����Eg�S�V�<0�T�t#p'I���h��
�O�icSU1�m��42v���b]؆b��	���;`aB���a
����a-���HT�z'�xB&3��vz�
N^��C'^��p'���{Z����y�)�ҍ|'��N%.ڧ�%�dҦ���v
?��j���T?Q<���hz�{�{`�&��`�Wv��S,)��eq��(����np#J]����60U;��2���k]���s��9�k�^��ؖ�
;ӯ�ְ�t���G�x�NV��=Ύ�Ō��mb>���H��#ƈ�I��$#/8h�Q��}�?	܎nC<
)[�I�v<m�ܯ�[pj}埃(�mcM � �I��k ��+�r��z�zlo yWY�*�	�?UI2�/� ��  s��c+�ϲ���T��|����,m�e	�B�-�>kY��]*th\
�"��H�X�2v{�.jQ(΂��X�9(XI�lw6������=��OG��TA�U{��2�������7i]�;���b8�UH��S.�W�]�^�gkG~�a�m��k�{�΋��V��_�!�F�H��r��H��!�Kv�S�C�buSB;�'QR*n��W�����3�%�4^�gH*B���k�8#��DۢAU1in=_��ς1�e�'@Xֈ��_���D B[f�us*XYY#&�6������Z6!G��Cu�mW�%�,&6$E����G�U}�5��S��u�b�B����7|�IfnX�\�X�qX�c���
�@��@a��H�f�G�n�g�`U(����\׷)�S~+i�G�+i1eh���F}gJ�1�&kk�x)N��C?C��$s� YI����!�ԑ/�x��e<��o_��0�l��e����g�]3$�Uܜ��1鈉2�mFR��u��"6������!>~B��#c.
�0>i��S�qRU�#������ے��2�z���!i�/|��Y�B3x��?l9�����=�~Z)j��}�B�x������^@;�V@�����{EEw��r��f���f!z���+�¦�U=��]K0���b1�5��p�������08מ �*�� 	���U�KܔK� 6�x�ս��+Ĭ�9�tg���`L8�
��F!���p�P�W����a��F��u��L5v��h�N������jvϋ����w�y=�lK3:&�$�y�;DǚgT	j&o�k�?3�\p�ލ�d!�q�u4�%�X�����n�A�`>}�6�1%���B�=�Izw���_�7��j"�����ƕ<7N��Q��!АW�$���(�`s��'>^܌�K���B(�3g|�u���7�x��45���2�v�md9;|��
�����k��6]��d{:g�%#��ؿu6��#"G����|4���ge����s*��@A�Ww.m��@}�G0�Y�&s�?����:��+���8�&�{�jq5�3g�+q,���8��H��ݓ����.:�m2R��Й'�)?�Z( �9 a/ W���x��&�U�x�V�xU����h���4����jq]�b��5"<��y
�=ԛ�G��$�2h���0��&��V=�k�b��� �O�X�#���"�N�� y!����w[L*�	Ri�G˛��(������W 0��>�bХ�Խ��"��x�u�%l�����ЅV��և��<�e�yty�=[�C|��'1�kS��Xf�s���ŕpq���?Qs]H Oѩ�6�A����`�3���`F�CL�*����c
-ge���)�I��&����~c��@g�|�����9���ٔ��Q���D���A�#s�q<ύ���������)ww+2���r���]�����o/G:��/�<1�-`��jg���?��ʉ�A3~RG�m�q� ����dD���U����r���\��i=��i�3�����Ь�t3�,g�uI/B�W6��dD�A6%���tA�P7��\��N��hd��>��3��~]����2M#�:��Ԕ>f��Qy)~B��#��Ѝ1؍ȴ� ΫFJ!� m��\�����#xj�����r΁9�X�޲F��Q�-A�ҫ�!D�ѱTe{2i�۔��*8*d�+�ՌF�Q!̔��q�H��J2�v9�S����^YĢ�Zg���ŋ���dc�7�E_U��۽z'���
8�֜_ٱ�sE����O!���ưy��pwC�j^�9�uگ.�:�`X�)���Ӡ�U5Q�d6�P�rؔ���ZȶJC"luT&y��T�k�k����x�{o-<�*�i���u
���v|�CR�M3�>�(�ݭ�jh�`�3ѿ�W�����@]����2���y����-{U#��/I��;��C��	~�k9�5����Q�(�M۸�d�V���h,���j��6�$,��U�����cs:��m��
�����l!T�i���ƾqV�:e��1��K�f;w	�O�欇@sD]��Wӕ�������f�jB�m}M�V�J�7�J@��H-IO��R�QR5;�}��b#��]iq�:�7�t˛c��J�WbmNQ��`����{Ŵ
��&rr��L�b�h|�>�3H�
�5���ѫ��1�\ry��-���u�V,V�g��"kd|��&��ܷy�9�� 	G<�MN��!'�7s-�.2��_\>Gy�E��Ѝ��g��!f�ދB��O�
�o�Ka��4�e6u���$��V*d���.)��w�q���:ӄ,��,�R�g&�E�܎J��ۂ�D�ln��>��3s�q���[5s�y4A��H�p}�X�*��c-��ɥ�2뮴����^>�B-��Y�]�l<��H9}+fo�Q)�ӄy�q%�x���Fbu��+j��,�S�i�Am��@�3C��C$�8�n�{yOm(	H�MZq�삺��w�E����%�ߙ�� ����������@���oe����/�fB6"��6�F���A9�� ��_-T�AC��pcܟ��NM Jƥ�N]#��6�G�^�P
볂&e�Ҝè�5Q�R���a4��ɍ�q�ħ���%'���Uހ��_�'E<�'0&]8�)�����I��I����6�MMd��`�~���^�����au؎�YWbrR��#���������P�iv�Gu���r�z�R�
�.��S��e�%;��;�)1XWW����s�M�����f�Ft ͩ�'Z�^��J RS�w�p��e�]��yzq'mD'��v��ZQ�(��(S=)������F�{L����������%gM�b;7��]��@�Ն�b�c�p�]6opM�Z2�9�3�����p�>-$��[Q~j�y�w�8������)�@�@�?�=D�7_�}d�0�0��â�ʞEM�8��I>���������:1�X�C+����S�_����0�v�B�-6�ln�C��%Q.~�]l���Z��}���1и��9z�V],
�Ù�K{�#�x�R��%��K�>vrT,0��gG^�+����CXg�S
�5S>%��+T^-`la&�2�+4"ƀ��܏ƺ6�4���)����U��ѡ�N�D�F")P����ke�]�	{���"�Lƴ|r�sÀ���i.�����x��0k���1e ��)�����7�=?��ٕY�/�Lܺ��V����<��3֦��U�����>7A�/h�bQ�솓�
\�ON�`���x�7y�Of���ǉJ�'��bDN��$��&��m��/߮y�H�{��+8��A�R�^4\���ӗ�F�޽e���P�|�|)��`����rxӞ�`;�Gv�N�_�}+9�p���&��\��0��'9�G��I_%���J�E�p��
xr0	/�F��C��u��:j�
�D$��v�5�A��vn�?d!�2(�Z��f�Ƙ[��#̜^�� ~�o�X��� ���������T�0Ӯ�rg�E^J8A�ɬT��������\��2�c�Ί0��6=��8\����
u����n�*�N)���GX&�햫��"������x���۲��ـ��ޟ�TZeS�r�>O��1iwMcM,B���$E��_H�,��0�F�Ƌ���9ˑ�)գ��?�O^�O�ȷ���Y�H��\c�Y��
�g6.ؕ_2_EA���s�2V>G#{���^�.6-�4�z�4�ij�_Ȧ���(����S���7�,@*�3%�TӀtR�	C"g\��HTJGFT_�xS�v��L"�l�jV�T�3�}:ؚb�۪8b6p�����x�U��n{ZT����ٓ>�2�9WQ��.Iy���u�<\~�W�? + �~G����k_�V	��0�FĢ�Ȏ-�pƏ�uv��09���ӏt�����92K�S�s!��@1N���t��wz����*Q4b��k�d�1�7�HH��?��P����a���W��=N�OB,3�=���}��;�j��7N�a@
\i���[�b6C�+����g`����'��1}��S����KTy`���.`�XW11�N��=���� ���_�KT�4B�K����ܱ1��kb-�D\Mn,���zx��\	����Wlq;ظ�����ҝ�;�ўP�)W��k�K�W�%f��^\��h1�py��T�:l��s���zʂ��)��;R�9�Ry�� PQ߉lc���N����_��B<t��ܳR��j�2�IiE`vo2uI[��p4��<�
�}sI6v�G��k�JƋ����5]�V0E> ��ut&�S���rw�R�b���i:Y�$��Y�VFکh~��S�M��{�V~�Q�"����]|��8�J�}]{iPJ-E����nF,#�?�ݱ��0��h�3�t��Gt��*�-c~"1�F���@�qg���3�v	����־���s��a�2CD�Y�p�M<g���9K1P�Ө�8I��0����S��rN�[Ck���q1���2���?�O�
FX�>��.*�c2�g���c�"y|3�",�V+E�q�Ծ�ϱC�WZ�|-�d�d(R�Ҿ���R�e'��R������n���­e��C.+�:������NP:�n6�r�+.zM��x�hg��J7][*J��K��������G�IS�	�����j���5�}L����a�&*��TR*�?���˿8p�T� kP�wD��(�{��Dx�w��ľ+ۀ̪�@A�Z�H7YH�ޙ-&%�m�:��;�D�V(^x" ��|
;�����%:yocBS���I+v�2�i^�����v��Z�� �$Ր���yD������b�E]b���xu�}�/A�����N2W�Oo�\vր�Q���(p�|H�n�)=���㷉jxCoe���j��N���s�)�0nta��������g���UM���X�G$�RJ��!r~�̺2�jw�*+}=O�G�cȫ
�Jz�"|(8(����8'#��SOɈ!�t��Biם���Pcp=�Z�sa�V����~� ɝe p��c�$�+Y���|��VG������V� �|c�Y:�S���^pf���[�O#���'��y�|��`yj�V����T�l�{�XdL��ԠBƒ�H�F�?EB2���֯�vКo�	��䦠!`�c�\E ��LW�$�;Z�9��$�𿒒���m��
�d��t�?�I��mq���[���D��4���B�P>u�ÎP9��l4�F@8�ޔ�h
_0<�|�੒�u��x讀Wh@1$o-ȿ�F���Y��:
5�M�sa���P�[�F�C.��v�Q��Y"ũ շ��9(��r:��s�?`?zкs�Ё�(joxy֑�6���)#��/:����@�����ԺK���?��3}R���ȀKί���8���JN\ס��o�Ax闒.��6W�p��f� %��M��Q�l�\��*�Z���=kVz���kG6o�X�H*U��,��UL"��q8O��?��Qs�;J-|Z�[�1��g�F�郾��M$~��p�{Y[�Ÿ>l�Q��d���J�:�C"��=�<ZS�F�I�XtO�����vu��5�(�*>�aCB�������|+�e]��w��ݗ߁�)��Rga�@S���WrV-{ӥLɁ������dAf�?:��͓۽vK�敀���|b,��x-�҈s�ڨ�)��Zil��c�T���^_P?��@���骋��!I�ɼ�<���#�K��Y�D�˽�
k/\��8+�����/�=
�"�U#0�-�]R�X:2����1�N1��\R���)�L�J���^w��lS�����/�E�h	��S'Q�@�Xd)��p�[r�`�Jv:�Z�� ��b�+B_���"9����o�Y��
o�ګ]���C޲����$���MQĳNJ^t�u#)_kR��E�".H��kU��L���@�0T5>��.�S�2uf�f?n(�,��*��j���Ș:��'�������{F@p�l5�AH�J�nhP���k���=[ے^{2��J���ek����_߬ߴ����u��G~@��լ�Iq1j�C�� Ѓ���X�;,�q�ջ�:���c����HF�K����7c�]�[��8ʡq��3N�v6�3\�ŋ|ɧO�
�@��{�X��k����u��F'{�8���&�O��v���@�)`�B��Z'����'L�Ja֘������z#z<��
,6ȐD�3�NK=�ٴr[�/��b�i���9��?��\��2m�Ȳ`v��b�� �[�7PX�
�XhjO�;ծB�b�A���4���Ϙ���Dc�^+��=�L�����HW5qD{Y^YE`����+ �X�L��Fvj'Yb�e�=qZ,�?�������}˃��}���:��5��$�'��R�7�Jc=�aWY̓:vt�;���^��U�.~5�":��.9SPs�O���v�Jq(U]��7��o�����f�b:c� k��X��k1p�C�_��2.:e�-��Fs�ma�QM*�T}��3P`��?~_Y��,;�A�r�5ӟWw�wEI�%���$U�2�Ʒ��������uT9�=����n=ʉ<N��ZSa�Kr�譆�n�Q>`�����"�s��-t#F��\��)w#&����J��	�Q��Φ�a�TQr�!�OJ�ؙ�rǒ░G`��ٽ�f0��w�$l�'ACgb�y�;7q*���3(#%��-3��ţ��T��<x��xv�i�GG����K�R����q�4����/���2\� ��p�)�������K��*r����
>C�\�r�ɾP ���UTb�쨠���ɁMh����3+��D����%�,�Ѱ�M����2�⊐�z(}S�L�i~�<�7�c�3�&po��o���+�C�jp9�סp.�2�
�=�#0���l�H@Qn{� �N4��eJD]d��b�&��o_�����H����Ä�	?yP�/.pw]�!p8�1���h��� ��` Y�Bo�Q>�q��,w:���/��̄��_m�P+�/
�]G3BL�#��p�uÏ�׷iyd�<qm�"][����z�/ RvE�����wy������W�����ﵐ�pR��G0ϱ�%��>��F�� ��1C"�M���9T�X�r�&����e�v��tf5z�˱sP�Y�%����}�}-Ɉ.�;!���B3]�Si�pl(Q}�C%�e����k0�Ny�o����@� i��B"���+0�'.���o
�E�cb1d��r񋬫1x<�t�(��b��Cn�w��@�ڟ]�zZ�ϞG(W\��X��5�gl����WX��dա�Iyn�j����r?�ŋ��FZ�y��v���9}�ca�������w����~,;x�.�M�v,)*�SP�81kߧ�4W�|V�b� �������-摨�y�4�ɽ�;kyD?gO�ƂZ-T������Ls���Ӗ�L�@���!}6{w��,X��O��l�d��v�~-��D>��a���>ޖ~d3Z�����~�����]wì�i>��$�Sw)�p�ۻ@~"�[eRǰ�N�
F��wa܊t�Vx��(�|�#�N�˛p7�t�����"�s�=���τ�=��p�1ګ�#�#ʑ�p�I�e�W��YƘJ'q�V����,���y���0�a����,Y�խ|��`[�_��*�0�p�����ft�܂+���y.B*h��H�n�a�;��+��іuJ����ʻU��~�R�Ι>���&yd���wtp]/0;[�*ZE���.v�����F�bv��9�<����|]���c1q�mw`�3_7v��W�2b}
��ߗN,^��KY���
~K0�4n���g!T��Z�)1 ���r'Xh�\��?��M"Ԡ��ȟ�ӈv�UP��ӡ`��$����a'��P"����?�#��.:U�<���c�;�ꔵ�s���uF�/�qp�J)L��)��T$��д
5�?l(_T��W7�cpt}����''2�^�h����S��~@���&����6�����l��X��x�f+LoB��lp�PfC�+'o�֭���Ȫ�eÏ�Yfo!�w�8cg}�G�8��Y�i�kF7F��Մ��yT��U��u7��&�
����n��=$~>)�6k�OBz��W�
0�T���X2�qO�d��#�j�7��4�WǊ�d>*�^D�d۾����ḄO#B�nR��@`��DĿ��+`�8��4�X�?Ft3��λ��i8iH���;
8���qíL-�,�i�q�m6�:*��op\�5VN5!��տ�2�$zY���;U��-�l>T�o6�Ecd�;�S!�c9���o�S�I�-��(!!�}� j>��@*��~�B��t�H��a����ԊA�_��50�Rm+H@sq�U���K밝��\I�����k��v�Ǎ���l�>���8SC�����⠮�+FtQ������$�AR�},�vh�<IY9��zc�fҀ񨙊�k����N��W��R�ٲ��t�jӱWc����P��L~��-!}O[!� ��nx{y�2V�=ފ蹎2! ��!�����D�֪�H�E����V�ۈ��b�����l[������P��JqЂ��D�;[җV@��ƈ��9�?�����N h�P���ۖi"�a�Xjr��V�O0g���K�t�x�t��:�-@O��m�!V�ZFXJ�t�]�8��t�1�-6"p�: �����D\nAg�^��FŇ�M2R9�R�"*K��٤?.��ZumҞ�L�(@��ߒY�gj��(Ÿ�>wB4`�T��u��1��C>_s'G�ތh�k[h��GV��S���o�t7^��$��������[�#���Vo]%y���ޓ��� C��k�Pb�c�q��)���rC�
�i�� ���=��U����!�}�
.�;��  ���$$2e k?u5UgeL`j)�sIk7"�C�b#�M���CҚ+k��@�<�:���(��x>hzˆ��T!���LE�M�f�.�eʏ8fn�bor�>�~�ɺ)e��D�#�GN���ː62K���Q��2���q���o���
�W�.�$׮@��o0�ۋ��)�,��s��x� 
�E�n[O���ͤ�����j����EeۏS�C$�є�*G�ptO���<�޾���@�Z�e�Y�К#�l|�2�̼�6%�{�qD:�^�����4��|Z���M�q���h�sO�2����vE���>d?��W���%#?I:r���p�o|.C� �u�<�\O�mZ7Z�򱦵!���۩�Q�O%|�/��̯�Z@?����IJ�&9ٶ��*�J��	'�����_�'��*#���L��%������5�+�x�	���rTv�6�L�#Wx:���]�����Q�?RfZWR�)E�%/_����)K������7Z�OU�O	���0+���3v�(���H��SS��i�$�vª�h�c��0��Zp1�/��DT�Fu��Y
^�c*�^���de�7{hyA~S�L*zb���<��R�����Up�ziٹ�C�,Z��(3����]w͖�ͼ�R�be������x0T�u�������a�R��[�bQF��ƅQ��ڻ�3��"�] ��s��\��3p���u���P;����Bf3l���{gޠ����n�����.��vQ�g�R����ko�UW+Ze(����k���^�j��0Rb].�I�t��m���d=�a����������O�ƝA��h�u����zD�,��#e��b�d�	K��k�%���h�����C�3{d�غ�a�	�*�v"S��������.��Q�i�z	h�~��W��PLIu����3�ڽ��d/����^�5�nh!��y�Q�	��p׺�����8 �Q�Q�,d��tqɰ�[����v�q�K���A%����$� ��.��hZ�n?s��:����c��\���i��a�˄&^�1{�i0G�:x8e�V�>�QA^7��(��$�	8 F���Q�$��:"8�Pbυ�a�U�*2���Z��$�$��� *s�
��ɍl��`q�Do��1ɦ����(����U���m�6����:�;�����å̚s�A��1�S�F�$G�(l�`G�T�]!V��-��F��)�c�yg�U��n�жڑH�%���q<��/-�7O�Ԉ��s�n:�?B6Y�Ra�麳���i���˝�{lƉ���sk��F��7r��l�H(�b ɳ��sw5[N�P֪���q�#f�P�%^�.ZM3�ܰ&���߫�eދ����U���d������d9:z��s�-!���4\��$q����V��%�����!"NI�g��Y����n,"�S
����"�C緱(��s��_���B��	1"]��&�w��[���J'rJ��T�V�6P#:���g�ַ��{�D�P���BI	�w�sY�����B�%��&̯��=�
���r��?�{���J.�a�/s�1�?�����x16/���# ��E�z��=��h>ᆅ
KM��#���s���wV������.����#�i��\vt��̘��8ƞ%�C��q����ɜX�Ƌ��x��� ���������k�l�D\هkκ5��'�UΕ?t(z������`�
�{�����:0�#���� ���Ժ��S�Z�ԪmCC�q<�|�6A�+ �gja� �XU��QM�i��>�:>2H*T�1a)/F̡W�/[?��rY�?�@�0࿙��DA�[���?�*(�/�.�~���G9Bx_ͮԑ�!�۟)�3?� *tD^El5�ff���~�}Ą�5^uc4�n�槛GvTVY�{z�����g%Tj����՟�[M�{��_
Z�?&���������f�UP6nS����=aG��UK�tMs��;\6��|��{w[f�SK�WXT�qr�aO� �+��~$~�)a���zX&/����IJ���&9�͐���קפ��Z96��nEm� h���4��?�V��?�҃Ӹ�A�&������P�q�i��\h{Ͷs�d���Q���os��?#Ε/�v61�.�������P�e�Th����=՘������?E�L�ߛ)�%�
�N�,���+�el:���7��3��>���Z~J.xD[b�H��m�m���<x"�Z�i����Nm��ڹK�O��@��_CV�IBҿO'�:�8�p�t$��'�w8;1w�NHM�,;I���	2��d��f����w�VǇ:4\������~U}ZB8T�aS�O����TtF��8P7�s�gH��V��Ha|��W��r� ��GI��6�Z�C17����Q�qn�Nt�ǽ�?�v&��Wk�o~i#Zܪ�8��	֔�[ii��VU��&CX�~��~
k)9��J�m F�^F�e��?��vA�����p��º�9v��aCOI�!���\���\�vʠ��u>����t��֪�ra,�FԴ
ἰX���_�vf��r�
\�/?	�2�m]�
BQ�����;���2a֓����<.���)��I �Ŭ����Ƒ��2#�d�z��N�V�7�!u��~PA����t���3ۋqi�aS�_1���q�,/���Fi�m=~3��_��ހ"Ѐ](+�,I�q�G~b�K��vbm6g8���w��h[-�H�]�{v���_��q����IR���"3��W3U�%�|P�n�8O�5���&��aޢ�&�-W��ȫ��3T�cW[	JCn�I
b�q^>��s��Pu��#�&u>���Ӑ�g��FP��B��]4�Tʨ�j`�dP��ް��u����Y�	'��?���,CQBA�w������u���Ɩ�t��k�2�v6�3͖���Ǥ�<ւs�r��my�>>sRK9��8]ҧ�۔ɭįT����w;A�>�zf8��B��u!�ƕ!d�ޜn��c����v~K�(ƒIzYp&��Aʌ��7��њ7>Z�/1��b���)��{br�������DN��C��?�d����T�%���>��z9?�ޔ��ٌ��7I�� _��|�i��z^�J�h�q�(L�NB�}��d��֙�+���D>��<���gҔկc��0�����ն-�{����%g���e�>3?s�&6��>d�Q���U����Ϗ�r��h�u�Ë���v��e[�����0�6s�7XIy%(�7�m'K�=���;@/^x����9;��L��w��ď���Ħh/�#DY����RⲢU�{z��0�͙X̆Yy��X���I�D���ǵ���g��*�Ȗ���	�J������%��N��$����s$C��!}"�Z��K|��J�T�#��dӰ�x�u�k�\s>�@�8ß��^1z1�+k/���~�%!'ak�ł������Z�D�J��8�ƓL2��E[�+���i��s�ٟk8:=�'��˖���Ռ�V	7�^����$=��L�Ԥ	`2$clq��C|����
T�%T>U��TD�> 
�w���GP�7#o2�B�;�p�Po� !�O�=��\"v:�fuN�z(���%S6�6Й�k?���F�2�	I�}��ö�g��O�C$���g��	���
�����am^�麮C��2�Y�:��p+����??��m=�Z�� @��i
ƹ���]�چzW,���K���ŝ<hRu�e��5�f�M�I�m�7W%/t��l#��ͳ����|/&/Na���$m������B)�|"��I��c	��.��4Q�zq�f�
�b���G��d��?
0������"$i�D��4w��%h#ʍ�A�.`��H�i��jc�a�D��;TX�MF�؄cA�:�o$m��ob���c�^�4��t_L��CR���O�N�v6���t��Ud��.r��ƿ��F�x�x� ����[��x8�R���t��C�d�֝��Eu	Vݹ��qJ5�ӎ�t�4�ɴ�������9��ڏ��4'<Wc���[׻�}|R~�9qu8 ��ae�jm-�}��z��a��t ���JN/�[�l��D>������.|H3H���X� eR�&7�H�WR�
�XuCiB0�����c���^nS������?���$���Qz�p�TGCsO��C�S�m�	)ܺ�A]h��PvNO��ߩo��)����	V��F����+\V��x0�:}����>�bydZ���g�"�w.����02�R�G �	��5��E��k���$p��C �%���zS����s������H���w��{����(�k3�n]@;L57kC����O�1ZDS(�J�;�p��"�'��>L�\H*�b[+D7�?�/z���[q�|��-�c�����&��=4諷��a/����Ze��B i�p^�jlΊ�yw. 1��r\�v�bZ	a����K���Ӻ�М�O��δ�Ģ��F%�M�i��ے$qqc�/�����C�ZG�|J��\\�h�,&hO�uwc��e|�2@ȇ,���l!��!�o��l`ۭJ��t n��3�����Cl�A\��V4K oZ�$��flI6̝͌_<�0k��α�u5�ʵ�Q��gF[k�F0���t��Й�_�z"h��Tp�9{��F��Y�B#�X骦�K`���j���杂��=�ϡ�7�4ŝ�J(gw	�mx���nQ2�:���=�=�/��]���9]���#v �R���c�);��V4�� �H|�0�{a�Am�7h.P[Bax��`:����߈(zjD��(�8�?�s ��q������f�>�
y&�ɭ-:����5w�%���kՖ��w��iw	b���+N��|��M6 ���_@��x��+�'wd�k���b�%�a���W΋_^:8n�S����"�G	�zt�'��Z��'��Wh�rI�0�Qk�DV?�k�[�=f}�Gb�ʟ����Dt=o�O5!߽�����m�ܢ���]/�s=_��a�z��+{[�~qzu��(C�O(C#��Xs;�}��E��R�{q.o3�Qe���8��6�V�u�Eǖ���8���XC�ఈ�`���+l�Y L��Q9�e1��`N>薑��0��F��3���P�`��t��%HӰ�h�JA_勤&��)1�'k�|����#5�{H6���~�|v��?�w'�^��R��0�x�R�k�tUX2p�aԤe�eq��kL�ʲi���H��͉B�(�V�������h)�2ģ��E����gq�� ��1FH���0�@���waG�Õ��DڊF���5��m6��B��TÓ��H�Dx���bB`��
�f<�ú2�e+�$X��]�γ���U�,]�n�F5]'�N�����p�c۶�lOb �ݳa`,wYYv�T,-A�5{�S�tw�I���X/k�մ��v����֤��q�^�:ƒWR�n�I��Qӿ���]�x}n��^A�IN�v��Z$2����E�"�{�p)��2�t�Wo�F��M���y6mdp�|e@H�+���@}9��������5�tz���<�d��r#���h��@u���:Y�E���l�����⪃H C,𼲧�,�#�&��TΖ���>ju
2[��i�=�tѢ<g��/=\�@��]i���)��X�{��\����n+(�T����W����*���L�]�<����{yu�h�,C�B�F?n��5��s�6��D �J�y�99���̯�'�P�IOZ�4���;�����&�b��"`_�ر&u�?my�V�l>�֘p��Z��^��v�d t�MB���u�:G��V{���x��j܄/@�x� �l0���.c����|��i:�x[�0�`�d������UE�HV/�����UO<��K!����U���OK.�f5�Ͽ�f��9=~�O��Jb�`C8��m_��L�JV���py��T\kƜ���:O���td�����v0 ټ�����s 3�6��F���B�z�G�+��M�/S�q�Y��"�ӻ�Z�Ô̳�CN��7����@o��B���u��Bg�k��$�t{������P��S�U��u�<��z��.9<%�/3Q�Inp_BpҌLVN0��t��$3n���,��Q�қ��Cq#�~G]�wa�I*|2v��,��Vu���C��c��^·��0c�o�*w���uɩ��ְv�q:I������U-����K����',\!���ygZwϰF��8�;�W�1������;�b����[�r\�Q
�<U%\y��[�v��b"�����\�.��5��}�R��r��1���
��j�"��{2����eq��8d�����^�qp�Rω����e���ۆ_����U�v2�6��3�ǽ#V'd�j�f�:�0K98&K?��k*l���K�mvXl�HR��:��ϧ �IeG� �6���Q^�^�V�N���^}:��.w�B���ܤ�.,�dp22X���.P���,R�:�v!��9^��|��z<� �����8*[�+\^}D�+"��)������]Wc0��[	�<���cAӰc����� ���雵� �кn5��볂qL4����(���$�K8c3����6�����׫��~��%
�lY����Ӊt��z�!�vume�P��4�����}\�����?yY�s�B^{'�ڐ"!��ʁ�]NFi�ƾ�rŝg7��������6�W>t 0��������WE-8gs2Ԕ�?��ag���L�q�箅B��,�g	���d�
Foq1�A�$�eO#���Q���H������f��H'*/�hކ�D���⿤��z$9����Kw��!b~l�'^1f�֨������G��AZ�`��ê�����Ho����R��	ʲ����i�?����$���Vy>���f�������J��о*�z>�X=N6���I�y��F���R밸vˤ��)�w4�R�q��P{���IXYi���]���wG��xj"�A�	S�ؼWעe뿒$yY��3�j��p��Ͼ�ĕ���k("�p��PO��F.<'�W
���\��E�3�F���]��4��A@=R���3��*���0��#�<��E�R��^X\��䤰�]��3<(�rḇa��9Ƞ7��S(0��nG� 9k��XƆo_q4F����K�d�J�6#=MbY �2NI.f%X�cb������9Utm���5��h�� ?|����9xJ= ׌0})�M�׻�띡++4�d%ryٜ��(�7�g��<QC�� HwJ�K�zG�
|-�[>A�t�O��T�R\AB(�N�5�NF0$��1��k;fe�r������+�I�˙��z�T)Bk�g������{����G.�����T���%e���흒#�~
;9#m`n������bkv�-M�^��;��cB���2+��0�n4��o�,.m��u��+ԅc�ô�R@[h���������.��sz�V��C� �W�p�ء�'Ox��ֈ������me�1�����cˢi&�4�8�V\EJ����ry �K+A7�Ót��F:���"�`qTe�UP�V)� ���?5<[�h���9z����o3�D6���tuay��;�)��0�u�1Cş�%�,W6�^�/`
�Cz�4/�]E��|k��&d��ݿ~ߤHV6$c	h���&,�B�$ϩ��τ�JU�i/_�E�S9��O̳Sx>�N$�������N3�jw��^� �~ �ߤ�0�o"�[�֙B	Pl�5u�X�̡BV�v�
K���:�	Є �����Al�N>��V˸�������+@K�s2��?�>�=�?��vi3�@B�t=����|pq@�v���C��a��3!+��@� uJ��r��4g���e5�)>�J��}�c<���E������H��q]��ddX����?$�o��NS'���8�,B{���>Q$6�&J�� I�ࠞ�~yu4��x����\����&0�t(�c�v0
�!�/����zt�8�60��N��Y�;�ѽ>g��mpVV�5�u\�1W&^N!��xz���dv��8Q�вvL�V�8��|���[:ǔ�N).�b"���S}U��'pi�+��"�����`��k^���´Т�C���}�:^�'���x�AE�F�/,��8�(��� @ɷ���
}�1���{���z슫4��}�vL6KE8�UC;Q9�"�)p ���g�~�����R�v
'��&�3�]<�n�>�tzx��ߎ��<uĝh�A�f�[#������j�f&B�<��朔�7E5w��m��H�M���v_���N.i�]��/��J�~3̮��"��T�1Zfܮ�I�"g=�������R��v�A!K�[J���B*+�]���V-�"]U?��'�/�I�Äy\Aģū^D�����y�P�np*Ƞ���cڱ[JP�d�v��}^�!�g΄�=��<=�S��{�$��p	�,�&�E�ܟ��}��3��kSTxX�u�� z��Q(Nq�O"��db3uBns��E�}��:���R/��e=�i*�W��j,x(���m�頹ܤΔ%����Kw� �%9�FS��d��hb��	��2�4�b
����q7d�JM,B�sv&Ut+���[���rY��]�aH5��'E�p�_ea�����G�*� �2`�S���;�#����0h�  �u�?���Rcѡ;r�����C�yS�o;hL�ڏ6�*[����+v�u 30o�v����{��[�1�\�i�����&|�۶�BP���zT�T������S����s�[_�=x�++�;��p�-�/�B���(�t�1��[����X�8*��rg����d@����4���؁��j�	k���H]�(kˁ{��m�`���R�"���z�5d ̥*}�t�@�9:��]�xS*�Y�m#�Ȯ�:-�8�Gl�:�u��cL���m�i��Ҍr�~�>�4T� ��P�o��P���h�Sbg��bnc�N��;U�R��S��ظY��h������ȝKq:I�hW���q�m�0�#v�A)4Q�|w������^�j��2���e_f/��)���[�����7g��u���0��΀�38��y�`�k[�Uu�21��%_���r�^Πx�a����1ċD ��H,~��t�o���b����͔]l[T�m�bX�ް�B��+�{E��r�Uv����𬾹Tl��.���������;8
閅�y2G,;�U�^�ީ�]y.5d�D��	��џs��EՎ�1ֳ��D��
��'��Ě���
kM'
��*0��
Dĥ�2Jݫq\�	� ��6���KhץnfY�X��Z4<��US%���x@�':���k�H\"�%8#�|-��ԁ��Xڥ�:���j��tHE�D]�B܆�H-L�KF�g�i�9�r�V���߾�~1����>!�(����%d�=�j�ť����*�,�1-�l���ˀQ@e�=+bG$=(����"&�t>A��ͮ�d�$��k�n����\)�����֊֞$����FT�mYϳ.�-�����d8&�4P���|g)�0nJ/�,%��*��hwC�� !�p�WN��H\'�几QG��C0˵��LE����<�]���pI����5xy�GEڧ/B�Q��wQ%����S�2�(�F�]��H�b�a���Z������ ZY�=��a��_��M$L�$G%8�m|76
R��Ε�ڀ�Z� �L��l�zӵޮ7���V�j��vf�CCm���7�fa����_d��@D�$���u�+!b�Q�jՆ� ��\|�\����Ǎ�n;��{{��P��%�6�1���I�M4�����b%+Zy�K�E��U��s�"`!��⎊[�Ō��8ٵ,K]+h��>�ZR�L���y@G�T&�
������Aq����~L��_��{ҰT�t]����M��2Bd��[��k�q6���b6��4�3� ]jF�zIq��kcy�����3�>�#���V��s�#���n�rK$2QI n�c�V�>/�,ՐJ�j<���Q��-�3���vں:�O���D��u���=�O#�<9ȧ���$��3�]i�1.�]���)a|��8�_Xq�N���rq7I+{��2F:��/
kX�\�D�-��� l�����f�j�/P�ӱ������î�<��uI��J��uJ��;�alq�n��b�.��K���)�m��'K��
m�p�߱\wx��N�t�(���T�'�j�0 �<S�>��ޖc1Tɵ��Y>���]���1�J��"�\V���EF(�+Uq���qA��A~��F�9�����J��'#�����1vp1�Z���Y=@r�7VK�^�z�e�ij�n���*��
�T9!m0z�7f1�ZLGW�� �/�������*	X�&�fgӸ<Eή����jߎ�;D׃�:�A��jx�� Fք>���.{Tb��ֵ7�>���!����b�a��TD�
\GDs�K���* 
8���l���Bm�n\����q>lް�ڴ���3��77p���Hؤ�	����N�	GWeL�+�v�cUZ=�<�/)�!�6�^V��9 Ju|�:IY�q=���n�y��s�_GF�n�-[��K<}�/<����j
>DG���@�TN��U��եV��u=Џ��X֪������4�oҫ��[����E�AX�&r�h���w�j�+�`̥��{l���p��1��Y�6!\�5z"��d̘Z)=���֌�
8��[s�Uܰy&�l��tc��E�^�΢�N23=ռ660t��`w�Mw���
��p/����X�a���A�Wy, ���&��=Ȇ�}�V��
ƛE� �,�:���[:�Y�Ơ�VK�fy)P1^_�p}{pPR���)#m
�b]�(G!y�k<�A�W7hØ�rT։�8yQ��H�A��ָvʟ2̊��Ӛ��m��b��M}U�h̙5�@��3���7RԐ����_�W��]�D���{�=x���Wa�=���`ߐ5y�T=�n�a_�h�ƳG[`���!��D^%Ź�}�Dy�%"���6(���YO����l��-v�t�v��2��|�t}_���w.���H�԰��i������bb�-\��n6=����.I�E���/��v�s7��?ad!`"~R���u�d�d�J�T8�_=�mwGQ����=%@5zD鋽ݪ'����Z��_Oc����_���K����l�i�J���oVo�q |X�+ `L��L�I���"�)�S@���N'��;�z�ܻ?���|�l[T�k;��|ό7*�IU�����kx����2��I<am b��}+��a(�X�c��u맩�iED�n�-�x$��bv��������bko�z�g5 F�wFku��=�#_4�D=�N�'���B�)�&>���U' ZHbdM��s�V&�B�[vX�D���#�S�I�x?m�6B-N��	;��R׻�ɾ�X&ț�D�&�}D����^JU�`{�|N6�6��P�埯R�"+ih<�ʚ�8��L�&�����1����|F_��V�p�W%����Q� ���:=���.�ژ��ٯ�'���HnO���+�<_�?z�!5k���z��j?D(Z���\]�����cT}����H��r��;<u���@��`ZLzMk9�Om�����p��3���қ8�6#$̧�f	M8=�8󣄙�i�<"i����$����ʑ���r��0N���'F%B�%Q�ݺ:�����X���F���ݸ_���W����q�s=
'3�T� �ứ��^�V��3������n�Ą�u���w��x d��_�Tn�Nm`���xF��`ƹ�U�U�9����e2y`��=��./�&���-�i�*Ta،��7֚��"+��4Ir��K�43�댮,��oU[U�џ�r5�3�,�I�vͮ��^��ʹfg��@���q���r��;5Wk��n�i�2X�(I������{[w ��
z j��y���տ��q�K��jF��fE�Ҏ<��Ԏw���P��d�P���z��,�p̜ �����޻��n3q�]�����s��1���><��I��]�	��ǧ9J炪*��f�u\'6=r�O.�L�4��)I� ���8���h�f��7�&����Q~�e�p���$�d{餄�F�/��a��ƥ��:]�:��W�J���"���g�D�̫�W��+ɣ"�8~z\���yw�!J���b	�[��iGbȵ��=P�v��ma���}��T���+��) Tr�@]R�8F��o a<�V:aH���ގ��x>p[���Q	k�9���gV)�U�{�>iR$��JU 
G��T#�a�y[Τ��~�0z5&���� Ə�bS����O�r��>����qDۯ�#9e(a�+qu�e>R�(�Z f9��X�d����yl�?�ֺ%]'�k/�
��WTU��r��2>�P�Z�7N@}\���o��o?�8�c�ӧ�Ҽ��<E��
+�+]YWԬR��������پ\�3HkV孎=��?f4��{d���/��آ`O�4��{��T��5���4��H�z �]Y6�@���eI�W��Σ�R]b}6�t<����Ŷ��X���yk��@��W���3	ZȾu�w�[�����GS46�q �����[$rq�;�k]B��cF����6��U��c�F�i���T�_U��y�8��~��1y�P+��6F��؂�˦����W����B-B��	���q� ���WL�o�P�nY���^����0�%k�KLa�������u=r1�\�~l�����@K�qNN�����ba/��5���Y�燻u!�׃m��c�����c��_�m�.�n�__ܶ�7 D|e=T��'�ݱ�daJi��_���a������,�_?�d��T��`.���a�Hz�}E�ȤK6B{�K
y��٦���9�S�2#?���7h�\�v�^��B!�}_��Ɵh��S�Ţ���q"���7� �	<��R�O�T�\�߈b�)��Z��sM]d�C�R�wų_��p(�H&S���r�h���|?1oA��̍����F򗛚�󿆹��1��T9�������	�0 #i6t^X	��k|dx��������dl��g���#�g#?�J:��-�A�kW8���u)!H���ߪ���w�H��m,���	�h;R�~���X�Q����,Y����7j�G��cJEĹ�CD��K`z�ܝnD��~{�@��it�U�P��Fe�������ۃJ�ә��~K�Wg�ix^VI�ԯ��J,\Uah��P.�6�*U��^�;��g�Mfv+��
�_���x��s�5�qLY�Uԏ�-����^����H�w�7���F*]0|��J��$�hb=|BW`}w	�lX����A�i���>^[��α�4�J=[���&c���U$�Q@x��؁�B���ITԢ.4Wa.^LBgz��J���>*S������2TXw�J!܃��;@Y�I�\l���*9
�+��_��w�TcQ�Yɰ�2�3��H�t�_#��->�.3B���P�^7W�?ߤ�iJ-���AKu��,r�!����At8�(�3�?�S�0�� ��h\p��p�����z�A z����1��M	�fפ���m�p3G!���/�[u@[��t	�dDC�@J�gRu~����Q�l����0�.�mW�L勅(M��w�wA��k���:F�^�E4z`�D�z�D��%�5����(+�A�Dq�n����ԩ��Ź$��W��%>��1R>���U� >����'"���h5�~�C�E��;E���9ԩs��H�köQ!063H�
�F
�tk3h���L�j�CH��$�������O�Ǎ�=�B�ʚ�I/�{?!10�D�	�~����� �i��V͂������%��?C�v�m /��A����ű�h�F��.C[<&DU#��P�u{�c�"�M,+��e����j�G��Bf*~����/L\�U�>�b��_l��i��C��;�[�GxE��b�D)p�y����"�X�3o�6f������Tr�/�U,���u�Km|�*|�פ��ƣ�ռ䭒�7ߺ�-�pt.Q��Ig�����!���W�р�V ��T�s����b��s��������dV.��lN�r=�Ҏm~����/�ψRG�  S���.�����%bhN�:;De9X���%M2���(%]�_�|h��g��B̼�	�������6G�Yb�܉9#4���1�t���;��y�-�d5�Pn�����ӭ-�����h�	�\�#<&�<H̉E�N��v�3�hkQ�O߇�-J�ʾ}L�&r5��Y�����������0������J`�[*/�r]�
��v���M�ʣNٽ��*A14��I�S�2��3���x���R$�`����;F��1��jqx�������dֵ��F�w���yt��b2=]�V�~`���7C��ja�U�ȼ���.�6�:$G�#E\���v��x�Ch���_d�)�p��J���l�Ml@�����7]؎Y1��췗����Df)c��k�]�v�D �U�δ��ct�悳>#x�r�eD������.!��2ͬ�Kh��A܎�͝�I%�P[�d�[��Vc����/5AÞ�:_;٘�2�r=�[��ynV�A�v����7.�Qi�c��38��_�m��'}gC��3��`�;*�J���L[t�P�-���L�T� ��=�$2�W5��H�e3uq烦��*m��"9�3���tO5"�c��fn�<9}�T�!4�0�hK;ǲ���Y6�ZG!ktO������֋oW�ڒ�oa���SET��	1�m����+�ݾ0̍P ;�`{�qٹ�ϓ[��H]�I�ś��k#W�<~���a�2���+���T����m��e�=h&w�u<	
���Ot��J�?�G�u�/��V�E;]�ʭ;:<�J�VĭhMz���i��B�8��Ѳ���ģ�I��;�B3q�Q��ƞ�� ��zu�}�hk���'U�ԅfC�(1��k֦0�G^�5!�<g�[�A��M,�l2�}���
����@E�������q�H�'�a2��T�]a���`��9������ŉ�����!|�U�Ȧ��tm"��8� ��
U%�m�'��R�~�ђ��Y��ڰn�07�����Mzn{L��*ı(�`�r�ǡ�~x��Է�����+s�U�B
&P����кځ���*B�?��8�[�-O�����ıh�ѪL[O�퍽�yV�W���Bv���^��ܣ��@��W��7ż]Y�B�'ˀ��o���d��)i]Ҫd�?�L�5�� 7����;W{d��'��Rf�\X�K���`\��F�L<x�f:�{e*�>�-�u[~�����ևj�ȉi��R�����.Qѻ�\h�8Rln ��+5�6�� ��s�lW�QR��*����W�o�za�����v���F�#�$��z.�~D<f�[�ևGFiy��YX6i~�|�s�S�m7"�zH���X_����k�X��Ef=C��P�©LP�N��Map�^<4A�[�����D;�>eRW�W��%�xݔ��:�o������^����{q2�&�̟E�&� ����1D�H�����,u���!KV�@O��/��<�c+�o,�Z�V���ST�6���{�aO!D�x_XQ9��?�}���ֹ�.(��8h?�S�!�.���a�{�QOC[���8��n��cCg�����/.��n<�-�b�9DU$>�|�,Q�$��.H�T�[��B�N��$����H~���\�%��S4�I��2.���T�5w�P8-R��t7���[9B�Ɋ����=4�2)J�Uh]~�?1�8������q6�/�&�{R�>oEQ��G�4|�P~:a�b,=��=��ͧA�*w"���8����7�@zr)r�U����r�P@�R,���"��:��9��M�|�2w��(_?���(�9���?9��tI�9����X��˟�̸�����/�"�N���j�)��~��!k�Dڠ�$�~�����(��jǦ`S�uBuAe�g+������<`��\�h���V����Ys�
�l�.?^7�L�Wn}��߀|��V��NSqk-�����r������>ϔ��έH�T��g�~=���R�콖�s��~���͎�j�~�x+��^�T"�_��C������,�0��' X�,ZM�-R[�У���B�����vM�F34_N QAaM�=�I�Z�-��eV#��p�X���\7T6w�fg����j��7�
���[W�%��k@K��P&���=���u7��Bt�260Q�0#��2��,1���`05�Z�u2��q�ɂx�YT�C�Yqe�$�; �<�6����_r�-��(��.6�Z�"O���]��>h�X��ʔ�=�%��x9��ANeK���x����S��qs�x��E�β�F#1w�|��T��~��D�1�Y��#�+b�פض�f?D.:q��a�ј��ҕl���/iIc���}-~g	TB�H4&lRZ��G�Vi7�Ϩqcb��<@푗<��p.�6�f�N�/�����g���|�FB�#��,����J��״Y���{����d���e1PF݁m'%�î
���7�$��}AE��#
� ,P�Z<=׀���[�G�ӝ�+�c7�X-�����?�d0>�)��v�N�0i�Cٔ$��My���б/C�M���p�g���S�Y�ma�	�����f�V��Y��R[�\�����2�f����Blac�eY�����!i�i+�<��T��J�`����yf��Ps��)<
��wBG=�6xe�������/�[)�Cb��(9ʀ!-�Y� �*Lå�BW�K@��.����#s}zk��;r�)��ӟZG��_2������]Oj��r�Θ�Ŷ��Z���"s�̫k�N$z�6��u����8I��~-��q�4ݳ$=��?H�O���ט����-�r=SvNZ�����?�[5b�b=�4���ÈV=�P��&ŷ4�
2֢�7�����#�u	�`q����]�{�2�"��8�����SV J���s�(�>
8������`�|�3���ʗ1������,���̑n/h)����Z�� d��Щ�H����]3"�l�-��1x!�gV�x��9̎g���,��2��1zۑ 	���xhƞcC�߲?}�҂R奲#�"���ҍ��ņ��G���2�8mR��;��V����̣mZ�|Ͻ=���P�����y�P!�<`"������	 BU�v7gkT��R�}�#ݠ�$��⎸�(��:�q-�]X��p��qfLM,j|L�9��i���gL��8���������v6Y[��=ZQ�|i�>I��%V�U�R�=��
H.�_cqyEr�e9Q(7�/�U���CW8D�U՞�ʟ.��1���֘1�\dX	fD��a\%�Yb��U�F�;àSـ���ߒ_7&A�
dz��!��=^&m��D�%�ݸL�����zH�Ŧ�d�_��D؁�-��5^���
��3-/zZn]�P�_tE?�)8����b��R��a�h}��i:�0�r�����X����s��� ���\�,��8uD�$�0�S�ACE��I�`V	۶�3���߰�����an�֙vmh����3�+p�ڄs��ڶ��蛟�S��z��w.b�ӣ���N��xϨ�^��r��i�A�����?2�i��m�5�YY���h�ϋ��S�G� q[h�����rYYj᪎�q?��t�cn�תl3-,S({��q��7�5���� �K�����`��ꙔSz�PPŎ���z�(�|��>��}56�%��赌���߂���2 T�,˃�T5ח0��5���v�攝Â��C�j���N(�)*=�$���~��]�
�M�ac)}�C����(^��Q���>���x�ȍ+C|fFיp���,V��/c �<�d����ƪ��̏rc�k/�7.S�h5�hՌ��/(�o0z��!����ྨ��\��\����BZS���k��;l3��"n�)��v�#Nc�B���7�0O���S?��ՅtRa�m�Gĭ�N1��
�IY����!��ۿ���d��&�imV�R۫������ܜ�Y�2-{�A�p����7�.p&������nѢ�N)�؇۱oM!)��|�ig�4u�����SA�+ΓǱ�ֿ�n��W(y�m�U�y)����g�-`��eAg�ߣ-����T���f9X�4�O�cz������Ue�
q4/�DXw7�� I�{��P�a�I��#r47�R ���͔�U?�V��L��X�i4VÆM��A��pbu�b��p��+M�cw���Q#[�|�x}d�E��b�_�|<
��#N�Gc��,я������^Vd�E�C�f�M���LÐP�w7��$�Q0 h����T+&Q�Qz��4}`��j���zƎ꣦����8����w_��:��ظ��y�q�IIp�6rYb�n���&�� P����!���nLS.Ӌ0�9�χF�&o�ޕG� 1!H�#[���*����76A!w{�&@6�C�W������/e�7������o�	�b��#���c}��ͳ����]� p�n�V��L$w��6<��]���O֒λ2mg��!2i�f���h��\z`��jY^ٷ��㚫�jܙ*���Ky�hh��,Q>���K�"g>�C�D2��R6-.h��g��d3�lx�)n�	@Eyro>nF����S\���)��?$�O��)۠�K��P�1�pȥ�@�� V��~�a�J���]�F�ߍ]zP�2j"�{�bZ��o��r���z���%��8V.5���e�jx��n��>�d`�4(���Iö��$	m�����������Ϣ�fk ��S�	Н�U����@J�z��h4�J�BKz��e�5�]$�0�6Q'Y��r	��0�W!�E�G�m����5�{�(YL������(o�	����� ^�z�N#>��g�c[<N
�7��oⳘCOT��+���1�i(���1M�7��ᙶ�B�'������3�r�Qr�:�[�!��װ��*�oY���|�K��9�,n>Gǹ}�5�v�z�)�ev�/�?s��d&L���T�Vd�c�{�W�l8����C�2J T�����
L�(3�j���vzF'��}�Z׳t���8�9�_)Ƿ',�͟���U�H�^�S�}�aN2{9�2s���I��@L���c%����Z��g��?�-�!�ژ�B����L���� =��L�^�N+�^Y�\�t�0���	P��%,�a�hB�z��z���S�Q6	�=J
^�F'�5'�a���L�|J~����s$�1�	��lE��u�P��t�"�獿��������ւ��W�,�5��4���Sa���Zr9������D?�I�:5Ï_�$��P���ź�řή�}Y�Ťlo���������+U��Nh��\n��z	�:�f;ق�;��*�)��M����D>����{�^�|���J��^g��o��O���Y����+*5@2�w�h�������.^���SՓMf��~k�L��yo�(]��6ũpU�?Nlb��gh:܌Y�ؓ��G�!�ů?�'�������]-:�e�U���M����+�S�=\�
Ȃ�y1�hn�:�����8y�m7��naf�����WlH��g�3�F�~���ԋ6A���:�2���bG`��R[�Y�J��2H����>� �����eZ�x������ְ���hi[���1.>����I7|I"bP|�&��5ND�MNmůN�e]�.~E���
��T�+���e]��cC�3ir����>��%�T���t���qL(�ѥ�^olU�*ŹŃ�RG�K�v��(!�s����Z��6}%jm��7�x�1K�a+J��4��(���H
u��"�o�,����èew��V���HU��9�Cø����nq|A�(�ܓv��bX����n�2��C�ĎSĀ{���8Mv�^&?]i�}qN�岄A0�O��p���c�1�ܡt�Ń�h�G??��>ǰ�[��5WK-;���"?�J%P������`�ɢ7��������!O.���q��?r�e�D�{A��´]1z��ӎ�P�e�z��C,-�6�����=��c�=�N?|Ra�4n��p���"��Yq�%�Ї|M�tϳj����%ɔ����Y���(Ȝ�ص��ڛ��J��cv�����:���/hr�F2��)(^�}�!n����O��$�m�9���iF�%�r�[{_��:q.|��F���C�K��]y�`�Es�b���@�\R��:�-���C����mW���6��LANA���B�2� ���tߧ��6�3
���C�N¸ˀҙ8��?*jg�|�Vҙ%	@T,�ɥM�쑉W)n�J6جE�h0�ze����7�&h�$iyF��0���X/�>����|_��������tq)�C�{�|w���5�{���B)�������yȁ�М�h����j��Q]�BF�a����-`�b�� ���c
|"��#D�G;#h��jJ��k/`U��h��=�W�o5��H�/�һ6Ӂp����E=��%E���|Bw'�p���e���|\gU{%`O�� ��3�2��բ�)�fC��W��o"S.9G:L.[K�>�"gw��T㫛�ވ��@x�aD,�/�9��5Z �}�i���>��%�����m ��t��]u$��:&] ��F��3�'R�&r�oW��d�&��&�eL;���5��������su6��������4��>Y{C����M�SS�м�������4ʆ�ֳtө`^��p����wѹ �Ѵ�̿9�L��z֥�b�z��V�[��DvYY�	3hs�Փ���sT���ZQ����WR�����j�Y�Qս�i�$�����a����%9t���ן���yu��.��']�s��t��y�K���o����>G�*x!Ou*��*/8rj�,3Fx�,(����hX�K<w!�����'P�'�����Sd��:�Hze����'�������p��u@*Oyl+R������k`͵��R���닚P'D�y�Q��g9�Au��{²�����0�Lq'j�N*'���XN>�)�h)/,��"����ӣ��	a�Mh�+����KZ��|��f�>vv��m�km�<t_����
��b[������,���5��=�P_6��C��2j�/t�<<�1=R��(}Dr�w���}S������$�u�G\��}�ң�L7���e�t��Iͨ37�f��&�5lıň���ާ-�p���P��9ޢ��2����������� v_l�S	�tE���\5�u'U�򳋈���P���K��
�B�GQ�s�,���0��nU-�H�yy��'�ZqY�'H�i�����Cg��T�>'X�����/�%M�8%�5�_y�t����(lh>��Ak��U��7�Z��hy�O`���z��gPO����k����\Qϒ���ذw�F���!�d��\bT6T.��"���[��[:�7�#��B�x^F��I�K��/�@�����0���z���x�Lm%��"�����Iό�v�6os�~���o��u�,d���}�2f4�s��{���[�?DH�"��T���OA�l�~�XG��r���#O��{s��q�V�!��|�c�2�%�G��<��2;��(����B�h@&Z��𱣨޹�7�DSN*7>���{�ΩB����D����Ɣ C:�;�G����][��_�>���U��*�<fT��sPdBc@Zᝎ��:������V�O= ��z���-2�TҾ�~
��|��	ȨiGV{����@�I{ڝ9�2p}bŌo���-{�8׳ ͌�
t���~��}7=dn� ��*�=X�DW�"f�s�jb*�:9�oM����z��2��c4�/p����|�#��yS���@`h)��y�=�49_�U��'@(��-W��6��<�
S��JW�7AP�q���k��]�}���HY�!��'`~�`�A��k�8!��]��wD�s�R����!m���<�+��C'��_�{�,|��կ�Q!�DC�����iO|ׁ�r7��5o1?~�%�;��� (�*�air�Q��K����7p�o������1���DG�e֝�ھ>�"Ê�E�C]�)&�ܝ�C)���bp�qZם�gr:���!D��^�P��̺��f��+�*�QN�"�i�֡L��(�1ʍd D���S����S�����A���I��sX$P.X}|���;&'9
�;��E�YC�S�'�n�*����c0G�O7a��%i�Y�'�X����_:0�d(��b���s�P/a��~?�c���w����"Е?����m�a���i�yD~;�����c~���� 0[P�{���U%�׏�"��X�>����n�Hz�=�Q���q`�s%��%�ia��ok4Wi"��?��#ӵ���K� ������I:�N�!*m+�������P�5A�4yf�M����}��g�<,B٨�L=I��t$���G�s�N�!Vh\�����]��~���+M��÷�tDa������s�L���e�峆9�X�i≮�D5�(J�i,�N��)G��z�i����k��:L%}���辍��h
��چqĿ�B�AT�#ID��>GQi���m_7哮����Gs�hw������3X������G������� ѹ.N׸�ge%�S���F+g� ;�w,ˈC|��];o>��R:����R�K�hf$���5�Ym"qz�Da0ou�������Eлh^��{�gY�gV�}	�g�@�ɟN���x_:R�=������V:��]a�H��z�L�a�ff�i+���3m��ϠW�� �z�^)�����7LI��oݤ߄B����.K�,�C���$�
༆f�cN&�a�������ŧ4�`Τ�����G>z�[�X�P̿�d�6�7�����O �"�d2��I�C��p0C����q�R�S�i(K'�r�:��������"�Y���D��8�A1���$��s5��EC�XX7�h}Q�RI���2��D�7�>�3Q��q��u��Go�\����)�&(]Q���p"�5�כ~��˟*]��1�iSVU-�͂�/W�D�"��b�8o3ī�L�#��Z�8�Mt�0r/@����d�u��5Z��fu���J.�Lr��dʧji�#�o�	V`\�_���~5&,��W.���]P�_c� �u�I�!D�ٜ�8�K� (,<0)�2��}�<�iA='�yq̔����9B�Ix?��0��T6�wb�4+b�;�]��g��%�!���bǌ�&����S�J�r����ߙ�#ޭO��(syf���~=~2]����G�o�0ʢ`��q�+��~c��^�W�ky���c��C�V�M���F��N?�T�k�FU�S�H2"|�?���J��a(�V�� ��'�u��+W�m�8���\w�N�#���2�H(�u<�a�]l	�L�u�a���H�����Eφ���|�Ś�L2[�{W�$S�S<��[��(�����M
�X��{�	�GM>�kX�����	�k���l�l�!��R��6v���.����H$��ƆP)�NԵ=J��T�x�
�缭��W�����yQ�����d+��V� dS�"Q��~2q����I �4V�`r�3 E�?E�i���}�L�?�UɾK�k=b������g3�M��E�����@���K9C.�V4��P%���� @[rF����h'����E�tV�I���c�����)zUD�����/�`��)�@��zS��a�4< 2�@�L��n��v�׋m�c̆8]���Vt����3♉{���FQ����*&LJR��1kqj�V��^zg�«ͣt��O�U�4-��,��|�z�L�i��A�M��k����ޮ{�i�
�_y�f+҅����å7�{5_�R�5V#��o�ڔ�5e�T�XR��~��2���_r5C�>b�l7�B����F�����*{�:�1"c� �0ܯ��t�4�*���z�L{���~�@�*w�����ȿj�����p��ޮXX��j�xXPmp{p������0
)���e�R��+ӮkY��+@�����e��%FB��s~�-�D��*}�:���RY��5H�k�VT/ { ǐn�B̈́_qy�\%|���n ���.q�9>懏��e���O@~S�d�p詸�t6�Ͳ�	�IJ�Dė;9_=��s�C{N˫�=��̈́�"z�t��t��������B���e"����F��~�G��3c`��n�8Llܱ8J��	�B�אG;=IT�멟��a��V���ח�6_;��ǭ%~����;� !�g��'�kl5��s`�zٖU蔁$�z���@bＭ��YY:�Bp@����6����2:�(֥��ns퍏���r$TeϜ��H�۫&��|�j?a���=Wuek���J �A84���m�
��M��Vh ��N"���~/����H�&�3��fU�/rp;��#��!�N4f��m1��G�tl���}4x�K�oħp��Tmtؿ���x�ǚ�8G׬D�v-=-q �vdtҚ��&{Z�r������V��] �j�J��~�ͺ���^j�"�T�"{��,�`u�c z7��Y�9t���u������I�����$S��i�L¿x��9�����Qһ=��3��5`&��mBkw�aA�a/s��QΚ�����s&L�e��*�2����(I<���n-�3�*&G�c��Qk��&�^D��6�I��w,e�̦�P��+N�3{��;��\������ɰc:=8���r9@A)4v�H^)��Z^Z��.�<T\�}NM��z�����C����n�`ރݫ�ttx�E��Ezg�wާ�} m)���!�L���	˚	�C�1`ɂ�@��뵺�a��&�x�t`_ëNL�"0#_턆�p��A���Yej9_��0OU��<���R�����B!\!;��V5R=��(�*X�u �tm(�Ɛ7�A�#QW���Q��'����E�k4�O)��*z�N�%O�j��2S�+�₧f��q �:�b�K�Y�ȋ�ۘ���	��?�h��4����u���C�3G��,�ʼ��\
R�s�|�ۛx�ɿ72$_1˸+�N���릔1��]G����cs_�k�ѕ�d2���Y��MnίeE|40�U)�
מ����H:�ZG��<�K��rI_w!<>$��J#9�b�����3��F$ȑ/%#�`|Υ��G3P{Qz;�
T$+���L`k�T xKv�`:�xnq2�Pp��k��C��k-��[i���Ji�m��y�k x�i|q
���>R��nd�z絛�2ulӛ~/u`�9�(/�9��P��^�h��Q�bc��m�w#�#
g߅��{
��/�1B��	�t0m<t�W9l��§���Ȫ0Ze�����[�˗�e�6��W5Y"���lJM '� ��y�	p`����Sb��N:�!�y�^Oc�gD>�JZ!|ئ*͉J������,���VG{��4��o�8����?���>����r��
��%��fKJ�XB۝?��0���|�AS�?Uc9�j������}�6��\�βZ���va�Ƈ�ฎ|�z��<��5!���p�`2#T��Fǝ�P�ɳ�� ��!���G��\�Փԙ����ږ�~O� 3�`����_��[IV+�R���s=z3�����v��ZcM��j�ں�kĮ�=}�s�f�i����E|{"5$Y�܌���z�
ъǸ�{������S��=b��|=�8|U��U�@BY��H��-�'�Efpd�RU�ϐ����}io��@Vi�g�e��QTX�ù0oz&̓�����@��Ȯ�(���k���צ*��cb�8��p�ǠT�{Yr���pj��Tp�ߤ��4�3�zc������+�I�{�u`ُ@WwY>tc��Ѧ�N����?��)I4Z�c-A�ц���c�N�/#������C�OeZ&�Q�YI�p�j�\�ߡ�r�=1<O�ZZ��g�E��S{ת C����p�u����A����G��@"� �fl�Ý�4r�ʗb�.ė�MQDF�[{�w��z�袨�c"A��U(�eRil5�V�u:Ѻ׹�d`[g$˥��)�]�(n�/���}���}I]ݧ�)�o�F�J�g9��{D�r±��:Y:�0o��
U�d���S?zV{㩓�	�A�W;Q:�`(/���K���d����I#���Ҧ�jMe�=�u�V�Qws�Ə���J�сo���>�i!'V��y<�O��q ǰ8��m):�Էۢ�䋈�72
5'���LW���SF$�W��� �N���Ta򅓛�ﺠ8'����6>������*6ou�CJ�$,%�l���9�zqe��p>�°�����^�A����͵	��oܘy{����RJ1�pe�0���2k�O;_��3��;.���ra��,*/[?:�zI��L���n���vV�qtP#�����=��Z���I�Z}�!�<��h�w5��Vz�~���Oa!28R�-�i�,�޵cw6p�jX�Ma���JN��t�i��5�n�[�#҃*I�up��sk���ƣ��+�t,�kwyss�Ч���X�c~�u�E��~��
Ե�׿�;��Rqv+��̩ȩ�h�ƀ*5K���)8%��-�R>uT��
�c���)KK�R�pA6�Q�jKNx\�ߋ�d�^49��l��/��4��#}����q�_�:+�Uy��g1�o�V�\"9aUE(R��0��*T��r�fX�y�|�#O"�k,��o�V<�Z���j!#B�"V��.�G�� 
�@�a�	c�kCq�T���	oGL��}nf����\GR �H�$I�z�*	��p���XX�J]�3�g-�q6���
��4��A)�ыCeJ��C^�n�r<ٗx��ek���$�v�c�6�����6��8��ّ�N`�ن��?"��	 X�uְx<�ր�Q]
3`8�Q6j��35�IG�j)J��k��7�����}���-�{�<�<��A*�Q��jY�pHM�6�R:W�ݽ�� ����fM��Rҹ�������
d�֡����tP�Y���o�FN��Uj�0b��cH#�MƖ�n �����=Wh��#����@V�����xo���'�G�K���c�n���6{�F��������diL	��s��:�0�e~��.ً|X�����LĨ�?���kͶl������a�l�	b. �����sj���-��Ќn��ld�#���aUR`�/�/].���l���l�����h[���!@3��y��6��[*�S�v���}l�;=8�����EW��z�hy���x!T���C��V	�ɷ�N�G�~;����äO�D ��<^\c�����B�����/��œb%�$/P�O�3@�����U��J�+2�tw�̅^��8�&���4L���֠d.���f9U���b��Y��:k.���p�w"��o8�W�33ue-�W��|b�PfN�>�1���q���x�s�xfMiϊ��6	�ML	O0���(�lu1x���8@��\2:�Φ���L,�w�������q�0u�)a�2IN���vې<5<7z���5��"ZT�E&�L�	����Y��'��gC�D��At�tm��ҧx8�=��Fͯ���VT�5/��`imp0Z�u��n\,d��%zW��:3H�Nu	f�9`�G$zB��!?��IY���n�'e�:~%Hq��r�Hx��\��5�r��ł�*�\��Hi���y��EL(��'�_g��\ά$���4/���?,�T7L� �&�h:�cˋzc���OiD��=S_r�~�"+%ҧ�2�KJ�!)0���چ)uOq܅��x��%����9J���߆�*��R�n��`���=:@c��� �Fћ��>?�;�v��� ����"��Q��G/����8@�g���d����^!<(�n��ç�)R���HS��=�A�]��� :�K��"W�Aa�w���{�c?�~�Ƿ%_���Lj	r�~��cNo�(�b����k6+�!]�3qG���v�B@������Ȑܔ{����_s��3Yan��;�+�_h�M�iկnI���s��u�-)�˳�ɼ����Fk��
ZӾD)��1E�@�^�47��;nٻ���V-4�����K^j�嫜}a��p��������d��eAE�D(�_8�$w��m�*�&υ\(�Fၲ;�M52�Ǆmfr~(n.��ZVQ~�4K�����:8}<D�C~��޹@�u�,�ã{��S�Ԁ5j�Xum�J��0� p��ҁ�k����J[���P�H�������~R��f������2�(��1����P`b�:MHz�X5�絔��6�?ci+$�(=�O_k��1�~*Pf�������X�_����?���&�͇/�'pܥ*�fPq�_y�t�+%A���?��uS#��V�H�5ZZ�>���φ�a�y�5k ���mf�tUQQK�5`����u���:�-�N�I��AVs�'k���@:��^�>`��ͩ���_�������ycd�3&c��@��x���m�wH9���������t��/D�9C:��~���~D�v�EE��pÜ�d�
�G��z�Yg�Ź}�f�`Q(���!����5`8."Z�h�eS��L��r�[���nX��9�/�Q��i���,�K�tT�}�Be�'ԭ�'�*c�ۛV��R�zBV�R�ݾVA�s�)�Ǵ+mtA3͛�h��4��є��~Z_(m����[�� �q�P?_�f�cg��]B{6�2Q|)�� |&�b��������[Cn?I�ĨkI�"�>��x�?���j�3�`�9�E0�:��V�F	pak���\" .��ͽ��'!��3���p�ӌ�j`钀���ҋ�n�?I���;���������V�ŪFC]�v)�+��=���.�2aQB����:ѽ��c߼�~_�S-�Q�|��Z�cK��(��I×�/*J�����Q��qn��Xj���-��/��?���I�t��w�'�V���~����2_�CY�B<7
�}za:㣩U��M�:)�u'����/偾�@�y�pb�t2Ɩ���]Y�(����MQ��[��4�H����<�9�Gy��Ƣ�ֵ	� u��H���>RBG@lq�BN�F��瓹�J�:jw����1�ؐWV3?	��#�WG2��=��(Q�r���̭RԨ��& �'�I�;��4�9Ń�4�r>e� }�,PP�=i�#�����XE��������3H����YhC��w��7k��'¤����=+|2�Wk��y.��i��A-��y-:�Cu-��/�u�B�b�VtNv�`�]q?N��Y�Z�AX �Ч7n�з�w�����g:o���b�y�b�!�nM|�x�4ˋr����r�U�1�б���q���(�@��D�5��9/��M���ޭ�G���QhW5���ںNSlˠ \�Cw�jF�ԣ%�����5������(��E�~��5�E�;�ż�&�f�@Y6��G�`��Є<T �}�D����8����d��dh �8�$���*�q�<Qo64�Ԏ��NT�y.��H�R�L�����6�!�_�#�k��ƀ��╸�!�ם�L�%*V�>�"6t�$�T�4��y��k��hz<m���cT�{��r����m�L�a|%FX�k`*��.�!��w��л�4(�G7s�=��G�o}�S�*�A�d�j��a���Y����6'��@L��F1wVb�B=����'�JXE�?���ㅜ�����X.b�_�}nW���=���sw�wmKN�^xV��wF����ؠ� "��4w�,��1��C��s�R�A�]������u�ϭP�՛��{O���9H������sܬ�mp*J�SCPI�kJݹF��Z��J�ki�������}����t�Jh� �K$B"��b���j�s�{-gtB_r�P��v��[W����ǩi"�o�T�iw���{�֘����Ҧt�
�.ƈg%͍Msa�a��;kG�Cj\��K:	�J��5,���ū��՜��N�t�?]_֙+�yw�D�S�]��滶]u(�<�S�ɪ���d�G�[��Վ�RX�b�k��\�!�BWlL�z���l .im��&Ѧ��\
�j/	\��k.=�K���H�clľ0��Ζ���${C[Jb��k 53l:c@��	�u��s�m����}���S(>�HD"P7o\
�����T\�C�`E0��OVQ�0M�zi$�k��wW�����z�NԺ��*�u(�V���L�O%ZԂ�O����ɥ��0�I��g�4W�g��� zϤ|�8^�b[�<�j�H���>2p	oS�b�!V3u���>���M��.8B1���_����C�\g�9)��yFnx���D!��_x��������bmTx;�ʁi�Xw;�X������7�`�P���y�����7W�`��%j�q���p��wEm ��@��V��S�k���+sl����}.D�j$�JAX%'7.�t�>y�u3��]�5T���XF�Oj7Q �+'�����3US�j���78�0C6����0�(f����0��o�ي�E1<��t[JS��GT��?��b��jD��$���2�&� ��w\��-z钎]�Y�ֵiJmF+8�y�Q�������#���D�U>,j�I}���6QыY$A� ���U�pd�?�R�ܗF�`��~Q����k}/W^4���r�!6�Ur�ݱm�|���+C���s~r6xԓV�vIz9X>xB�҄(���L�0[��d���������/�+���*�����y)����5�z��}h�T2�| ���|��ܚ���������v�kgo\AF*����b#�RG�ߒl��Z� GCz���˹yuC=�D������6��5����l�zmYJ�e���UBwۀ�ag�^?XN0klem�����o/J�^���7I�['���`������S���#��B�(\̕�.i-�cY�i���d��,.�+�n�ɪ��̔ ���\�N�C5� ���Ý���Y�-Qi�ax�t"���WB���l~�J~2�P��\���Nt�4�/Ϊȉ)\˰􁾌u���;C�Y���ǳ�&���7��D��3����fT�x�>?�����i�*'p���*D�ҍ���N�]m�TT�������}{� �vF���͞���$�[ъ�C��:���ukT�p��:5~d�ʯ�9����)t�o����i���h�v?	����K�6�E����]@��~R=o�����U8�~�c	���A���Z�`��?2��vD
��G��1�0���۲<��!��	�GNA;I��K��M0�$�?�`Gu�ۤı���E��Q^�ݴ�z_���`���΁o��2��}f�|d�\ed�u+Y���l�Z�DJ�N���Ւ��,Zo�m'��V�U=kP"�m4�3�!^�P�%���E�36�_�����d�ף 9�t���.T渄�ѷ!�������`�@��Sf5>QF^�<F〺�P�)z�M�gI�BH5��J#����d��y��=>x��)��j��n�i�M�V��j
	�Д��(h���c(
 ���j�7o�>�w��i`�����O"�a�}�Rb�s0g���˼��ʏ�$ID��f5(�3c"_��Ԏ�g���� ���^a�r�V�#��v4
␖�澳C�jd~���!��[B�G��n�L�L��&�j��.�$�l�+Ȝ�вs0�\�������wB馛;C=���+��"�od���5;��*G��7w�6W��\]�|�~�W
��~�GkuL*�G���}tr�]T��xo��/�����Vx!"�Qui"��龟o��w�チN�q���17AE���*��:KC�vm#�u���%�$k���w�/�bŔ(U#�2�(��$8u}��B;����,�{��&���]�m(@+�6;ߍo�8�5�De�� �� 0��!շ�<�L'9%�W@C'�}���m��9���s���h}`�- ������K���c��%�E�`��q^ߐ�	O�2�m��렧+�x���m�b{ޛ��8"�T:I�v�Ӄ��+r�`믡l�3�+e� �D�oXI4�Cf�^榘ջR4~��K��;����j,��"�MR�nC�{�n��9���quhM��o��.GK�e*��7����n�����2ƅo�
' 	fS����%^���$<׿�^�}�\��\$F�H�H⦡�4ގ�>:@�y��z4�h��>� JE�Wq���'��0x -BO ��4A|�%��؆�+��C_ʆ�W��ȉ�`�:���-\��o���y�+�}��(F.+G��zt%�AoD��̞�ZS܍��B�k��� Q�݀T�D�O᥺+yj��$�Z���\�Ic���^�1���1�oe�ڵ��nl&������GSN#������yəe����+7Ԣ�������	\��#�|U�@�)5�q�Ҡ����|��/�Ío�0�!w�F����9�rXc���x��)�o �Kq^b���s����� \�=ڄ�hm��y����v��!ֽ*m��*h������Y��!/���Y�[+3tcK�������J\Ī�t9X��gy�N�?* 6��^��iQ��ȖD��{]z�����w����Ɉ�5 ϓM����ʝr��XV��T�d����&�?6��u,甝���1�)��Cֵ1 ��8�H���a��w�<*r�Z毈9�gC9�1{L�y��z��H���o�ac�,�g��w�?z@E���ߢ��3,�|��F�^������va�?�>i�0m�|��5���hIW�>?�x�-s��V�(����v}C?�HiNZ�.�'BWǂ�ܼ������[�e��_sp����[T�v).
���<�q��N2|;�I�s��b���46���/����q&�e6[+|��V�;�yHԇ��
L��G��\�~fK��(8�&]��#I�R�J,�y�/BZ���h{f ���OZ-3~��b�w	��'&�C��=�	F�qb�L�Cv���{�E�J��}i*�{��(�;�����ۻ�h���� ����׵����T�� �M���fOV��UF��@�v�.\��� �uP�ě3�����80.��hDJ�*V]�}U�����s�o؟� X@+�A�"|��l����=֫4���M��O�<�S��j�8���j,��ޥ�_��[�o[�1č�g鴆�
�o�T���Y���*rL�>�3@�IF�1y}��;���u��U�j���DqHOɊTf7�6���6���i��=����C�Aec�J�%���V�C$N��ZZ˜�	a��)'���sd=C��˜X�c�-N�(�vȄ%�Y�k��PˉmJ%�~��������/�~��ji�>:P�QW�kx�i,��Vǜ��c	gH����J��J�0�y��7�zK
(X}4ϋ0$z|x���8����ۑS��,e( �ܙ�dK49��s���G�cK|���q�;���
23^Dh�yѦҳ)K�8�=����-��tƄ������Q���[���F�0�ȏ�
�����n"�1��lE 8�tI}�3O�)I��I�ę�Hy!������������M�{F���*�.�;���4J�K��d���»�ޖ�L����q[��1s�Y�-�,Kȶ��)�.O�e^�Z9~���J����q������\��t��h��K8p2P5/76�V��ߤez��}���<�B_Po�f�rЈ��!xMI��C����H������i@Ȯޠ�ʒn�v���)ʛf�b*֮��hڲ��ٷ������c�O��8o]sV�]���=�O��Ƣ��5>��t��WR
Ņ�/���s���S[s|V}^�`�j�� �!�Og�/�%��O��(@���pr;����0�ĝ�.��Ft��x��-T󽶁v'"%��-.�b�,W:-��"��|g�Ow�#��38�p��-�1�XXK���@�;�-�:�׬�m��d�x��d=�rS�=�����ǲ!e$������gHY���c�cG�nr�#�lJ�j!2SCqW�5��j��&#*��tfc�|�=K��,��U���S�F���ue���Ӛ�iZZ�j��b�>K{��Ϯ�k��bp|j�`4� �)��Fj$|�G
3�g�@�Bqh�"N�?�O8�����V�y4~����)~���b���UbB��-Ea
@Y�i���X
b�Fݞ�#�D�x�u�+��2��GƢ��,N�TZE���]YH6UL`�ϴ�SW#��>[�y�QS�����b�}�q���P�4 f�cY�!�B�,��Ci\��Mo	��A��t�� /	 ����%�M3ބ2��#:�g�*uZ�Q�����R_0hM�&Up�6�D��1˦P�,a\t�����ղ}���ݠ����G��������tCCQ���(�k��e���\;4&g�Z�q۟k���H�Ъ��&�J�,m�]%0������'�U�L��Ʒ��:�\R߆��c�.4�	�u�v]{���>��rD�9�\~���N����,i����;��X*��ݎ7쪺���/C{mK�¶�9�go��������A�"j5(Y8u��9r�Z�)o-T��Lg�e�v��%V�&�o�T�偸�ѫr�O�owؑ� S2����*���4ȁsKMxؔrG-��9gT�@80R���KFC�ɵ��`ںL�x׻�tH�&2�<5FG�p��f!�aa'�������=�|@����U"v��$O�'hE�������rJ>;֛��h�����p�D��d�e���FD�̂oH>�CU��D�f,�K`Ƌ���Hp�.��:�b)�l^�Zl�0��d廰�
6���v��|*����`Q"vx��`r����6X�粕��#zsو���2,�SȀ�J.���՛�5��:���t��q��\=%/��|0ٟ
���
K�?A�fҾ�i��ؖ�a��՚�+��uNM�&;��c���^���q�����k�b?B"�Q|�T���+
Qn�tv`�ӂ�����H�͢�
L��u��}��U�tf
1�5�u�[��}L���ğl�(����?ò���?����6[���_Qg�i��nR7���+��1�'��:�	~LI�����-MG݃`��� �9P���Q�~Ʌ���-���jiR����j�[S��-�����(YK�ud@�ʆ���a��^\��;q*{~���+����m���!�~ FTMD��vkM!��ҋD��Ҳ��o�_x��U�ë!nf��;xt�ɐ'�~ZC5Y��w��Ӷ� �7@�;7��ǇQ�z̳4�ʄe-3u=N� 8ɇ��3ql��l��N��		�U�>F$� <I�
�! �U_8��&#��:?N`��e�ױ�Փ�������K��\���\��4�GMY9� �-Wa@����V Jt=�/�j¿�i3Ǹ&k��G�ɑ�����Y���b{����j�w~�I0����,�m�8�[ۤ���oB�AM���n���OإS$ Tmt�
__�(�P`�3�ޯZr���eW�j����l��B۸b�E�t��n����[���~/XOS������L�n����Z)�c���Q�
b����Q �b��N��$Xm�-�Ŋz,ozpRQ獙�?Кɼ��i��h���)$k$��ܬ;RX�@����K� ���Xtϧ��ՈU�d#�<%��G��ZX���P�ܣ���_1�7�\V�ʨ���6�'�:���/9�����P�=C�&b͇�9i��9*ɜY~�.DԚ�& ��%/lg�I-���e,�]j����2AO!H:ey�6L6}]m����kty�ܪQ2`IIz,��{q��AW����R�懛PL�xu��E��=0.��3t����S�G�J�Ӗ�M��{�5t����͊�F�L������t�d�!�<8��4�b���R�p0*-�%�:p�&�w�[�6@�)��5�V�[b������Ҝ��Ip��Ze$�����g��7���7I��3���ɥ��T�L�)�w��n�tғX�4����~�9�.�w(���p}�1���"a����8�*��k~#^�p3�ݵͯ�s ���$�g��qJ�9'?��/a��̫ם���j����s�]�`n�B�0Fd�${{Z�ڠ���Zo��nD!�	5���R$&�-�	�4���-iVCa���t�b:��&T���~tJ�)W��K�*���T9�'�R���~��Cdxq�6Pއp}�i�E��uk�O���qS���?��n鿊()��B�Q��0%�Ε�O�?�׾��o���rP�ǉ����C��o8uͯ��0�>�,����WE,���}��#U}�hI��Z�$�h.'�Xr�k��Nc�H$�6Y���3|����(�Aʜ
���@�h��Zl��>dWM�^���+[)�wΩ��9$��U�`�,\�/����
���p���?�����y%�s> ��f��qsH݄'�e�Y���'�3M7i��gT�f��m��N����F�w3#AM��f5N�/��q\���������s�U#��'Q��°}
���ߗʗ��4�B��<[Z:��������=녵ƒ]�d�����2M��q�=�m�Hr�:��SG*#�If6[i�;^��=��|RB��	����.CH�ů��5�׶����5\q~�◡�;6T35�`o�W=��H�Wl��{��@\�;�du��m��Vq��gK [q�y�h0H�zooe*��~5�-=�%�|A(k{3������kUf�a#.>�����O7���B�n感�p}B9|�v�Ս�,��sTN7�p���$�l'�j��*�9{A�GA�u�������`l玶.��Q�P�~�U�D1���u�]S��S��(6e\�WxSSBG��J9_��<����3����T�q��K�2|�q��h�K�F�#u[�/U��a��� +](��)�o\�ő�#7u��:�S��T�N����]=�������@�5�Z�����#獮	�3U��ߒ#A�6ʟ�蓢i���(�z��-��V/#vW��s�y���YD� ;��v�Ͷ53�ݕ���-ޝ��Gq��W�t��a��X�Q�祝Mݺ����Z{�:jk6�@��)���I���eX:.�0�e�W���R��:��`�����*��O|�+ �/��\�'є'�~�֍N����w�0a�f�W�)�bnm@��d�+�M�o���_ܹ�d�����I���<��S��A�7zW$
v����1�p�J�je���0Н��3O��	��Dm�1��w:��O��b����7�E�#�b�=I�@Nl�������9t�a�{SWgjqf��0(SI	���6�"�Ɓ���۹R�0�R�t%�zL2\:s<5����9g&Ӧ�4���� �,�����ڍ��u�e���3�/��̮�+��fh����:.���t
����U'��3h�\m��¤�����؎%��X��k�On��g���A�����[J|����OˎM)�+���wϕ�C���U蓍��8;\�Z,�7�6Z��{��V�O��^��,N�:�Zu����9�)���#*Gvs�ҫ�w�-x�g}h,���堔i��v��O�>_z�㢔���R��^��J�v@}�#C��e`?.��)�'�Ӄo�SRە:	'�e
� �r��zm���od|��iU#j���jw/"@��f�`�8��R����՞D�畋\�|����X�ɱ7@��	:հ������������c��<ˀ�)�n��o2*j�5�37�+|��-̐�,¶������7t���^2bl+��9�w�����?�Dϥ�s[���O�gƟ!��W��m��ۥ_z��YGS8�(�y���RU/�-��]<�C�\��6+{7k�1^�t��Ӫ7�B�MD~���w�%H-��Ӈ�.r���XLๅޔD�̀:�L1	��z�������%��zޱ���	3�*d��wG�^p�%�`}��J�bX�)j�+�����䨹�g�V��h�( �k�{�{u�_��V��#;���Di�/m]�\���3�Γ�h. ���F9ٟ�3x���B��VR�4��.P�p�0�	�	�I���^5a"�Z0(�cH_?��G����<k�ߖ}%�TjR���B��>�Јk�� ��J�.H�_����W/k�1Yü�.��%Q��cs�Rp��|q3���5B�Xr�Hw�?��EUw������/À�&ٮi�]�b�\�Yr��V��'�ڿU�t���d��ط&HI�]L�b,���d��^�I�CK��z[����iBŐ�;�0��m���2m�4mz6D�V׿����ź� ���>�\��,$�Uw��D�'��h�Q@}��*n@��_=TE쇓R^�}�.or�rJi����查̘x���H«ٌ*�#Y�M5���5Z��l��v,ߛ �'�*7�\�4"�vŷ5S���{q�9�a���YmO��b�ޝ�G��$�W_b$U�� ����Z�sW ���6\�
��rOp���e�J��GQ�Q�ov�	wi4=F�햎("���dY���f-��{O%����S��ٴOF�-�8������\V?47��_�s����Q��[,a�j\�y�NHH�Z�q��,��*�+q�h#���ҹ3�ja};/L[����č����J,���]���=mc�^m"�?5�r�\+T�iv�{*	Bc�ӝ��{g8E%4��V�%�ޕ�������?5~'GK��gj������4��&S��S�$ɚ���I��t|�mp�v�k)t�TR �*]�na��y_%cЌ���Z�!]>���"�)K���x}]	�� E��a�d����a�1J����'fM���W��x��u��=� gm��:��4���&�I �NX�ߥ��e�o;��T��#�/��R ��)_y��?�@𶤟�Þq�@Jy��I�:$�U�^��$=?�Y��a�#��O[�i�m�k�m��+����3]*,X�hš���A���
���3t��,I0"�uE>"�v��#��*�����1,3���GlAsG1��:�A�=IC�'v�CKB����Pw��k��;�F
��4���������K�g��9���bҤЕPOp�
�Y��~o��k������g8C�Gt;�S���d�דB.�1�!g�q�����R�=��i=�	�<F51��,6�:k��A<*}U��RS_�O|���(a��{��^���dk��%�K������3�OF��ȗ��׸���-�gK�s3�#[���j�!��cq�&���X2��=�7�Q��8�f��:YD����k3b�\ĢZ�|z򻳭���F+C}��F�W:�C�b�6:�5�h�d��Rj�wQ��⽖Ŧ���L@�ċ�b��#�6�4�rz�J�LN[-�ɇL�ͼ�v b���Y74��A�伲�}o��T�&%�v�����@�j�2*~��Й �j������Լ��b��`��3��5�t��-a�m3�|)
΍4�(k��0��}�`�mB	�����)�����ԧ�e��b���|Q}���'a>p���_|b�puJI� ;z���ӈ��$��	�~�)�)
@����0�G2�J��'��$�v�.0��P�|��]����9�8v�E6�>�\��M����6U)����@�����31�w튍�t�.qf���[�f�}:\i�{o�K#��ʌU�b��,o Iu)*���|}AQ�7�m���O%&���~5�X��F�n.��ϑ��V���e�
���g�w�-�g�DWv��w�S��h�N�7�=��l�f�bSު�w��_%��`.�;f�Cˎ�&�
�Q��AA�@�̋�1�����}�VQ�P��k�@ZU�_]� �������܃K8 �e��Z�۪��564t�Em��v3U&����2?�8�1 X��A����s1�ۮ������C!=��'ja_ �*�,�$�!��>�U�����Ra[��'k��^�,�p-�F�V�4��kl�9,,�a�iS��EĎF�� AV͕�[��]C%6�eͿS���;䑼agA���Q������-U+��������W��yE�A�y���'�]r����	-�O�̥ʺYP�Q�2�z������ڑ�+��\�1@�l�~VD�:>gC���,w�%{�0�#�N�����&e4�N7fJ����>�[�� n�Ppw����(М�3J��pi���ֺ[*�'6b��G�2��){�XS�	�c^Ȯ�q�Ζ�ʎˋ-7#8Urf܌��W�~��<\V4�%��D�GT4_.��8U�$���e"Z%@�nZ���,�,�']���l��(�#�&��g=Ǽ�R���v��%��χ�"*�'"���޺�F�P�|�">�@���EN�������r/�S�a�m�	�Vo!�ى�{Qٜ�YE�� �lo��;�7
H�jc�?�[O� л���1~�7��B�J�m%��C�>c�.Z�..��Կ��n�ah�N3���϶vɋ1.�%��Hߦ��.pŚ�l��d;;�+[�A*b����,�Z�u��{�7ǑҝAr
��PΞCN�ZK�X���i�	����jo��]����G�J�^6 ��c�VV�-�G��ƺ�oX58_�n[����w ��o�o���{W7s�j�{$�+)=7R��K�)Ƣ�N�+�xu��6w,B�s��S��y�1�:��*������=�o^�x=�t1����5(���E�_�M�_J-(5ՙϱb��yf�L4d�\���tq���*�ء3�ɬ�r�w l�Q�xm�R
��;F�-��9�\G�Rě��ұ\~��Y�a�|y%.���>짻��8+r���+�g�kF�Q�\<��#����゠~�R��8Dҫ+4ٲ��N�)�W@�nW���V`��+�����,@���Bz7�I�wz8<�`�^)XR���>�00ʬ+���!�Mq3�Tk.���#�X#������>Y�G�֞
^I�H{��R�p�/5���ڢ7#g'MaZF�)�\jO;�L�O�~PIv^���0)V��C]xY>�ԑ�
��7Ö"{��7L���{��CZhl��u���S[��v�-�O�Iey�}��\٫acM%����R��
����a�;��zw��~ �Ev��42+ۤF�;��Q�h�^\	Q��U���p�$ �}�D�4���LI�`u���T�\�"��15j�{�uk!8T���#{�L>d��06?&���\��ޖn�?����x�5�[NPi�N��W��\�*%:�.ޞ�r������=xG�SF P�<����(���혼�������^�L��@�����i�~�/��q�l�Ȣ�4�P��o����)2U���\I��S��S}��y�O�r$>�|ƍ�K�������ā�6��̹���<�TH���Gz��2��W[t`D�Tw�<�7 N��\u*��9������[둨K�[*�Tr�2��:GVq�	/�p?(��]#
6�ߏ�\bcN-D�_�.�HpqRt���r���zψ`�P������ӮJ��5X�V6譱��	�tR�*�)��Ga?:q�\���y����re���Ju��)T$.kK�c�?���]��H��R'xE����e  ��0��r�Cwo��JÕ}Q
�� �2�}��{Z�߇��>���������.F0S��[X^�"c�˯���W�T��C4omt!�`:�q�l"�rQ�PV��t�/�orMiD�u8�t�y����T��_뙥�v2���S��=<���5�Q�2>h�.���<d��B�(��_H#�T��_"x�Np�.� ����.�)���i���N{�Z`@ꅗ�f|]���{�{^���g��:�H��M�ݵ�����B��2��Oc9l�2,QT��<�;�y����6Hf]�S��\�._d�tYD?�H���	]"E[�^�&���P:m$��b]_����T1NJ�8fƊr�m�`�w���`�4�2��;��A d>c8�9$M�Ì��	���WJɳP��>�:˜���L�ɥ��~ �|�C@��;	X����ԊSp,��:�\�;m$H�6��u~U��<'����N��UF���^y!t�k�>r��ʟ��Mj]���KBH%Q�!nDt-�㺘oa�
��̣��ne%���@��
�Ҟ-��>��c ��1ڑ7�\�*�|���w�}] [�Gz�������*�|.]����/<�9���� �>�xGt\��D!��� q�4=�����xY�OE��wzP���4���Qz�Z�(J*��NM[C�>S-Po��Q�d�+'��ޥ�uPy���ԑj�~�o`�QV��m��Q�GE$�3�@4�:�k�u���%��o�;��ؓ��`���km�(_g���Z~;dA'�>Wq|LJ�[{�!ۣ\�/�C��4�`ѓ0 6��PE!�IA��6�a�?���
Ȃ�.�T��3��k}ȶ	��2��RAP[��܍C��8�%�'��O���)7�Gt�蕢kpڛ���L��-��R�RU���
��2I��1�#M@G���c��w��2��n���Z�"�|�	=���Л��Q_ ��ɻ1�w�����,+�tkN��)����)Ez���s�*�I���o��8St�Cz���v�9ER��".�Z��m# ��X��<�EEUX�\h�rǮ�C�!G��0I��@�pH)e%m���r�̵07�{�#�~��-2G��ɸ�y����@L0$�\��*{_�����6PH�tW�JQ��� �	^v�N����7���f� ����c��C�]F+E��fN���Lm%@��^ʼ�m�3y\g��%N�U�o��*d�h{'C�`y�zf絒���a�2wO>ͮB� v_[�kl(��q|���8ψj��`$�o�,`�x+1�C��Q�LI3@2"����D�^X����z��-��߲z9ۂ��z�n��jŞs'o5���?��R����4]Rl��~�|�C x���ĺfy��v�V�1D��!	E��K:��r��-SckK��z�=L]�w��bC�{����xj�y���w�G��|Y���w��S������1|��,�juك:��\�M������h.XK@;w��0�DK%I���PH �Fy�rt���i��=���I!�� �X�q�%r���^���/s�\�~r�6	Y������D+�g���5-S�C���^���l�.�P.o��q|/-�,g�;��S��ydi�l�yFi ��H���b� tt�Y��͕<�o��<s��w��
�"���d7��ģ��"m\Q�ڧ!��Ƴ�AE�V�D��?>�H����s��\!A	��YЈ���($�[�����:u�����S�C����n�!�^��^��'9͓k{pob��P�<^��&{W)���a[��Y�;ޱ{�A�b��jÓ{�Z��L���M�O�飇~B��/ߑ��O�"~vV8�\W�������"sK�ꘪ�Օ�!t��C�8�%��7<���.<��fC���M���%,r��}�k����L�L2Sc4�ABȔ�Q|i����!��i5�p���b	惉cʢ����#�B��p�.��Jk��j��<�F��U��H��Ϭb*��u`Yt��Y�sa(gvFD���WҠN'�i�?��ʤ�@��O����ӟ���	oY�+L�|�g����q������/�ʡ�w&R ���T�J��*���y����*Jr�H��^�&L��Z���[i&[d�X���#c[���AS�lr���^խoC��� 3����|�w��u�H�~�x���~�VZ�<P��zD�3"��z��̫����f�QC�_qi��(4{E�f��bjh�`�i�g�i\�h��o��N��Y���?7bG5Ŏ'̨հ��߂S@;�PsK]u���&�N�-%O�?0���Y�eLxl�c4H�٥>�ϰ�3����cN�
/+b���n�C,$�?��5�S��͖4T�(hQ}*����,�]�j"�^�fd�����f����H��_�\�C�����ql�K<��a�'RE��|���(ma�I�9�VH
ˮ��=���΀�Zց�J�����|�-e��'�*z�|�xc�iB,Ycy�6h�~X�'l���wa!���.����o:�6u��=m�K,^RU��d6���o���hG���2�Я6����.�P,FO���{��}��K�9�Ɋu0���)�W��H��R��D4[�E��xk24 �ۘ�G:&�@�C2玀���@`��?'�M�y/��ٮ��E}7���-���0���p�����ގ��'��R���d����=�ݣ�I^�i��& mV� '�� ����1{8��bk��u����d+���&F�1�a��/� ����c��"aD��y�on���D���%�xQ�+4�;!�g\�7�������Co�Rxi�\�^��5{xmU��pv=<(�����A�M�.��[��M�"}�ʼt�[�m��EH�F�+^c��H�_�V�9A{}	z��6T��s���&e�:t����2���Ŗ���e|�	�Em�Ơ M~�bՏ��މ$�4�!KG�;r� ��S_Xr~���%d �bX��.T��ʹ��c�����fh{��uc��H�����Tu�Pn�Uw�+�����
�����t�
�w��j����s�\Xp��q��,�mW`qŉ��,}�#Y����ƿ3�����/�Qѳk��7R�N2����%gO����СfwB�������W�<�r&ʇ�Ѿa�eQ�F�==�k�S4�aP������ڹ�@=�Q��� f�xm�e��_h2���iiR��§��<��ģ�(L������f�$M��l�I_o����{ *>j����] B�P�h���
*���& ѱO`�DZ�y��m�Ye%�[%fj=�N_` E���9k���N�%�qD� �
�I�w`�~t4���s�DЦ�uѿ(�N�'h�MA��k+^@���\��uI]�"Oƅ��O�J;r60�V7����I�N���m |鞤��?q��)L��(L�SZ��O`��z�}+y����i<�4�B��g8�]h����b÷<u���Ϊ�I�3�(��Y-�k�7&4��XqM+�E�K�p�k�m���z�?[��]�\�#�_�[&o�h*��SWNr[���*v+�ҡ��Y��ZT �q��\�D�xo�P��Grހ|��.RX�J�Q4@����E��X�oR�^�$�:��]�%�zJ��=�t��y^W~ou����TsA �����=NȳV��ev1G#�51&M�p�kh?�z��,]�G���çG���E�-�^b�Q8&�R4���G�v��9�M�6���M���X�a?;Q�o��ǡm�u��D&XO��=���zj���/wj�]��Ts��E
��[#	xe;����ɻ�T��_TcOa�NO�g�!_��|U�ٲm�9�u
��^ÿ��4`�A���L��~��Ț���j_-����P"��RMjHn�18/ ���őI�8]�e3�w����	�-?���<a��7�s��7۩���;I�M=��9Ur�F�;�����ʮ^���д�Q$�Z���k�OC��dZާxJ��EjMH��T�hZ?np���,i4/�*��"���ySw{c+W'����8�' ѣ�,<��t$>v� fG�szA�;(? ��\�#�)j77�6� �S�
m2�e�P!��;��$A/6q�HKU�
�PO}�d@����e�t06�B���gK`���!�Z�&+-�[������h�"*61�]P�w�>�f�B!=(Z6�	���#32�	����.�}���]4���YM_@
1�7	�7tXsUғћ��0_m`�b�\��h<����<Y���RUf��4�w��(�Ek�\����w*����e��/��x�;�Ʋ�=/�*a�B�.\��F:,�e�pG�	�^�G��O]Z��G�
���-��dI�Mu钚��'򺴊n�{>a?b_�%���S�#��*[��Vx7u4�<a��l����e	,	)G���hu�O��$߇F1��Xر�[ +.Yr�3?�W3�;�,�#Ж
�k�V*�Ȑ�����,���O�i�����<D6� ��Ry]w�?��>i����Ȳ��9��c �Z��װ�c�|i�}p�6��0U�w��g'b�2�	��)������
�+�p� ��b?д��{[FJ�b;�x�N�6.�� �*oȱHcB�mI<�]h�E�l.5s��N��k]u�Ѻ���|o�Wk[M�xs���ZG�~�ؚ}EX�8��	�Xc�e>�A����im�b5NQB)�׸����Џ���i$��M��ӲS�y%�h��$�e���3�X@<��֡T�	�"��,�$1��c��y��R��||3D�?�V�����n��q:<���i	��������/���X.ǚBtpu�>��C�%�!�YV��M��^2�vd�a�{%�]aA�(޺��������MO�+O�n/$w������MH* q����������my���[P_��������;)�O��~��Y�����s,�������A�f��9�����R���k�djA[�b��{���F�L+�`�v���R1Lg�x~?�!��ɲ"�DLǤ=b
��`�s\&�$��ւF��yŝ��Z�e�J���;$���Հ!�M��������/Y�(:�^jo�f�b8���v}���&�d0�u�Sـ%��ZnW�瘇����o�3�����=�4�?Q�)ݩ�
�;UP���N��q�^� ������&����1��N��)�B_՚75o���@����(éA�#�zV4�U�`���k�/���r���� D*���Ԃ
��\*R v�����Mğ��S�;P��t�vg6�T�/����*�*�6ҿ�ر߈��c���(ɾ;0����H99B�S���h���bl�kz�l�A�f%����cɚǪ��|un������x��MkC�?���^7?Ic�}@<3��CH�H]\�1�X����w��So��d��8e.䋷ךtTt��r��~�A��Z�!��a�@p�T!�=i����C��-Uy�&#6����/�
�E�nSӨЖ�гp��l�4K��$B��W�g��b}J���y�%�P��d���f9��d�;�l(k�d� �@���yoB��U��NM�N��N-
ƠhYҚ4x�W���!k�_z�hJS4�'�ix!������vsw#�]t�D@���Q�"&�_{GV6}g<��v�T��+m���&�e���\�hP�xQb=p<y�/�4z�����T����[���V0��q���ſ��y#OE[� �?��8�a�X�D�Fe�[�&��`�B�
g��g,�2�XtX@�����|�H3;��HT��A��A�V��u���=?z�	��*y�#b���:�v���ek�ܘ"�
�vy��ɪ�b�0����?#⹁�e)�;3pU����gڗ����Fu��Y\��>48d�E���9_���? <�a8��([3���1md����7S/�i���n��R��QfY�'�ԕP�T�E��9���{O�ۼ�-ϧS��*e�H��ޞ<���������E���n���e�z��@�=�n�������������˄�֛�*r��d	9U)�0�阰D�dQޟ�v�AvT�;�Ԡ7�E�;�\���bq��z��K�`�j�<J��cJT�n��~v�Ĝ@<�_)�Iץ�b:`r(��.T�+��K�=��(7_��B��a��\�uNK���1��2�;GP�ے+h��ϙ3v�6��
B���+12�N�����%��U"�*W�^����-w��?��4�%��v���2��g�F�u-I����/����=�|�4Aʾ8E�!��.�(�z�9Z�cR� �����wh7�-��L9��A4pa�����W�򦑶��}ol����- ��D����0��[]x���>�;]�7���~$���|�$��A��t���a�:<���"Aԥd����ɮYƩ7�N�S:��߈�N:�}�|����qd}1�Ɵ��q6�id6��72�jsᎹ���
�h�@-�5qab����KG�߀bd<�UW��e٭2gn�O�P���)�M/IKF��Q]߲w���!�<1G�]z�M���.�U������g,�SW
��'�����eஆ&d��\fIUS�7�&v�dj'�;��q��@W>��������xD�DL2��D�y�r��a/"(�
3Dא�|K2.� 	\�WJ���éO8[�Ƽ�^2�����T�#�.Rc;U����I��i~U�87MX�@���kqj?O�or�jBRq�U�Wޭ�?����i�tۻ8A�N'~}�rx���E��OR���18�q�]w��ً�:ٮ�Pg�G�h�nFBu�ȥ~+?��ȸ��:�&b)Rl�e������ ��/E��ՅG�o:�^ƴ�1�I�*�����~���q�Ѳ�2�>�.w�t�i��F�L�V�=X�'B<Efg����oڕx*�����Jw�1
u�Ċj�u�X�=�*	T��@ˍ�׍ٮc ��]�&���Wg�*��_��c������
�z:&�eX%k�-����ʼ�����N#٭q��HS��j��X��,���=*�X��3�܆w�B�n���Oϫ��N�>N^ W�]"�`м�����N��}�*�v���?S@����
�RJs�м�rs���J4���fH��l1���I�?#S���GA����q�m*un�o�TqFTjG�������x{��v�CY�o�'���0Qz<-��`�ӽ-�{�7��{�~KÀ��l�X$��:P@��������2���_q�%�H����E-|���#��i��Ŷ�]ٿ� �x��&���>﯏�9xF�2^�<'�!�?����du?  ��"V|D��;4�N;NY��c�b��H�FSH�-8������_}"n�����+������48����0�����	^�9��w�'M���A7�"�*>���P#To�9/�&�Z�'���з�hV��멨��$俣�G��f_��-@�0�D.�������U�;�r������(G�Q=w��]�̻�B�vh�����<s��|PFx(>w΢Թ;Y�x� ��+��V\.�3��r���W��3��Xy�^!��
��y�Y2��R�4��C����1�-H^:+���xuE���)�36��Li��F���buг�0�y?�Q�nW��H�.��[+?u;S�/�EW� ����""��D2���yճd����ۦ�Z�J��*߅8�@\���W�ַ���KP&V_��MKЅg�{�N�>������PQ��`��HA�@�*��Xn�A0�S��h��8��bG�)k@Z���*6�U-��O+M'�'\��X	���L�"'�'\��AIխg���̈��5�\�r(AI������X���/��{C5��@�K+�{�:S��P����@��4��/�Sj�w��a�W-B	�[P��)w���sB����w�eͮҩ�m�X<�l�&{�"l�4��A��4�Kɽy��r��.�[;�U%����<h�����7�_x[�t��Okݷ*O�:u��4�\�͵�٤#TP��{K����p*E��'��J}Ώ��]����+GZ��+s���ȫ��XGYD;�u���O��Zx��R�aQө��{M��R����߳b4d��,n��
��i8~\}X&����ԣl�W�&��U�L�E��eXk�@�����>"�n��P'0Ė����#@��6�Fq�S���&p������pR�O��|�m�����K�>���0[���@�Ԋy=�:��e��{�խ�u���뷻�B�= �Q2�[�G>�>\��4,�y+
���\�ȑ�m���S%����L���}������@,���m/�\���2�rg�)}����}Cw������}�lxF�>�Q��(�v�T�y+�tEwQ��
�:���3Ί*[������C�����)������#G��k� ��}��Q.|��.5�%�O����8���|�H��>Vrx��;���0"�CibmyD��]�($���7_;�M���@9��G)ҿ�lɻlT�g��t�y�B��l:�\�B�V��"�WTw�V ��ע4�H���w��펩�g����i;+ �6���?�9�4��	iN*u�W�U�Z*(y����6�UIBs�"�H'����ZKA	Q��d&��.�GZ�R(�%t�ٷ�����E!��3cX˰2��{6{D�P�ń�l�}���y�����!:��X7r��Fp[*�A ���W�'`7)����n��U�}W�Kސ��K��v��.�����+�	�3�w܍�G4�[����Qt{�r�uy�3�5ʂB�٢Z��u��N��3�f����V�|�e&;M�`���[e���6�h�(E��N��G��#h��I�\"���ϻ��p2��˭�U��ֽ�-����i#�;��!�z?�꛶����=�7��$��M8 �����u�k�K6�6��qs.Q6���J�0:bÝS6�������!��O`f-����B��%��B�77rᴓ�A��O,j���6�|F
�H,�L$��Z#�Q��w����d��RUf�����K8�a��옮�E�>c(��.'�������~��=��A���ŶT����Us��J��:x�9�U�?PWa�se#fv�R�����&e;h�8n����y����ƾ��WW֟)s�����Ԙ�+l��0���C�5�q�}�!��m���+�vJ��B��0'�4���q-2�����L�Cخ�N�h�+������F�<�+,i��
"�E�3��S�
��~a�,
BE�G��FC�ܐ�܌�z�D唠BI�r����,n�?z�]����Zz4صU�}`�޼��4�{1�y3�e�8Q�r\�����L�H����X>|e�Y�؋���p�y��%- �Z�&����{O<a�c:�nW$��+;_�f�J'��1��gq0.�L�ς�0z�r���������Ia��O���f}
/��d�0��,�$'����0:��$R�zvT�����1K�MxE|uk�#��d��0Hd�F0p$� ��'�u�EhF�(�� Bo����2��e--&h8g/j����e��Yny�(�����N�7�^�V��1�E�l��G-o��W˚���q=(��wS�TM�8��1�'ǫ�'��Qˑ;@V8!�=]͉ªy?�l��+)`���%Lg�	8�r|`���3����/�����$q��@����_�RII�Zߓ�[+�M��]�"��Cڲ���8,s�����*l��`�Ú�_��'s����
�O����_�7Fױ��׹ɥ	e~AK
���{�yQ�,��%�V);<�i:>ݷl�?51&���ٳF�4��e%�=�έR�?c��6�Bg����)G�#4`��'�{bt*�}���y�"_�R;
EӺ�H�k)j\�����\�{��*���B�:u$�62/��v��Q�!��f���d#��d�����0�l� �:(xR�)�}�pR�|��R��<rU.�����^-?��A�p�oQnD�dn�tcݳ���Qy�|{W�ypY|v��F�(m���EA�����2łKV[����,|�������E�0̘N۽�� �`�	`���>�2`w�'�@֠���(3�\&A����?��K35�S���X}w���6u�9Ӄ �[�� )|~��S!l�o�Żl	o
7aƓ|b��Cz�
��W��oX��OUͅ�Z����Fl¢�����,��e��ܴ#L��������
�Q!	o�� ��WM�JWv�{�����8��~HpP�څ�j��jn�1?�]!��B�׺tA��N��Ŧ5-��߻��FYIB��ߏx�9Kò.��M�&�� ��'���9nG�B�_�.<��X�������e�g��pLb�7��<�RJ���?�k�f�#R��L����c��t����3c�eY(��x#��������{���Qz�
�ZR�M��*uRd�V$���]J��%9��2Y�V3�L�\����w���Z�!Ո�F�|]���%%H�]�	�Ƅ��Q�������8o�tn7�\ڼϦTpm�ސElx�p�4�Ҷnha3b|H�^$�r���~�Kn6cA��;���Jze���_FOfE��{^5'�+��6!�1N�8#�)ُg���nk�qn����<�.{�F�]��dۙ�3&p-�c��w�Ɖ�u�E��z&\����t(|C��F�
{n���s#��nH����}�<��_����/Ϟ2t�Ʀ���	�9�
w%��("�Q���#t3�s�j���h��ɘI��)H�`g���Lm�Vف�S�֒�jK���tP5��<@:�a#�>:FZ S�/�N�|���g� �@��4a���y�M�g�v�W?;:M� m����Ʉ�	
��?�D�2EW�e�J.���>`�%�t_iS���;�(H0 �C\�Atlr��F�"�i�)t��t��y�IĝG�3z���׺�g�6��3�W@X8���nж��D��IW�8�l��9��.O��"U0��@/9s�*��ⷧ��]�j)s����������vF����驑�>��KZy���W��]u�G�����b�úDpڵ���k_Li��a�G�̇��el��b5�[l��k����pF9�U���6hyz�@�G�uu��+
�^u��'Jz��lw:/��_nz|��N����3���GA��8)4�pƓg[�Y@�#vߺ�Cms��]�����K�B�Zɇئ[�u����L�c� IŃ=�Y'���׵�=M�&#�Zy@2�*����KTP�p�a��5�3s�I�[+ʐ&���$���h�r���ҵK`���K��R~}�r~��jr;ʃ� g��]J:�a��K �ߏG-�F4�AD<X?ӣ��T��� ���<�}'v[MFڍ��F�#���5�&�v��X���}�	f����إ��9�#�2�#qZ��ig���NQȭ���x=-`>To��Su4���b�
�=`p�!5���p�0"z��>v�;��o��h�đw
�g+U|�t{���䎗�e#����<��F�0��� :���f'�����m���%Dj���S�R{�}� �d��~�DE�y�ǜƁ�ڙe��>�'S���`ݳx��m̬7�u��IX���-̋w����B)|����yC�b�`W������㲚9�?�`��+�;�G(>��ܘ����q�vK�BC?�'���+��nټ�\���z�5L��0��6A�ͨ��}��
LaX�^��{��<Q�,6��%�n�7��E��u7�����}�#*PJ$��q��<Bb{�ߐ������T�8,l��V�Mm�9�٫�sy|	��׻8� d�r�4XL�@ad�0N�u�$�
�x1i��W5j�q;r��ſ�?��VE��.��$�Y4�OIjF��8�U�_~�UpQZ�d�M��W�z�U��vv��C_��9k|v�d}��2_�ç6ާ۾���%%�&D��D�Cv�}�7l��uE��2F�#�H�ٿ��^R���j�X;E�r���m[�ag�blP��)�5 �0Ă�@]�޺�`�89�~��mfb_��1�&"�^��~�F�(h��������Ck�����S�%��a0�����R����>tg��6(��n�m/���s��]��g$ؼ�IC�>;5�9�Rs��
�hX�*l�I2~�qY�'#�[��r�����q��`m��?!�@pᤥ��P�'�5�6��'�y�bkc�=+�d
��2����L4_������X����!�;�-�,ԅ�$xLBg�ªn6�~�;Í7�O~�Yc��U� ��>\ �}���������Av�ތ�Niϴr�$��8N"	:V][���CH��� PE`���.����F^ڸG9'��T�ΫZ
�vg<���"���D9"�95�N�P������۠��:�8�4�t|��o8�V.��;��9��߂�4�7`�	�\6�Wś�V�\�U����AϏrd|��`�d��w�P8}�|HH��7�R�4�λF�%c������O�V�he�ܤ%R�=@Ȗ���_���O�&�%���؉�y��|_pV�:.�C�Y��Q_>��t=z^G�@)BF��C�<
�� A�HMV �M&��"5�v�V�z��ʺ3�m��1
#4? Ő EQ�/gA	�8� ���vk�7i����Aߥ3	�!��J�g����*���t�xWI�%��Z���}�q��&��ܧL����H2��.�<D�G'�~� 	�C�46���?(�_NT��)���x���q������}ݰ>��D"`p��z �R9k,��������_���I���epl �d!�����ha�`-Y�u���K�>�r]�D6L�6#�d��)i�=���f�
ͨ�.����#�r������'����f/(Yb�8A3{�s;2b��t�؋��氤�Ne%$8�؁;��6��?~�'�z2?���Z(�]�떣%�L]��s~��1�V���"D
���NL[b7*������*&��`%:u����-��'���G��~�¿¡nRS�"OQ8���4��N�k���%̞k��*�}����6���Nڒ�A�6*��>3J@�i�����t��.Vu�	�2Dp��������]?��o��*l&x-!3�#�+ۭ
�h�u8��(�xx��Ź���
��J+ q�å�ĭ��ǰ����k�J�.�	�T�챪!��[M2W�b��ǒJc�0��} �ll�w �#���ߴ��_+0{,�a""�������ӫhS���db�.#9ѦO���I��D��P�*��gP��~fW�G� ��m0����o�*����~��<Q���v�	;��2H�l�A&�M�2��0+��&W�P��H´�'�5���t)�.#��w�VZx�������(`Ɩ����eh��ks]4��ۜg�{�׀LZq��U�6u��1�����w�q60^L�=�'��u�k�h`��9M�����iR:�i&.�F�����%�<+ܩ������2t[p�k�>�	��*���i
^�1��r|�BiP�@`,A��Zo��35%�zyIuM^��4��]�4�a����9񫻋���vA�	�0�����DC����y�q���Z��oe쎔�0܌�B���y����\����l�.��WN��=KBm�T��X�VM-Z��J}ʷ�r�G��WF��}_�����S��˝�D�2��k��������uThjT[D���Ұ*��
���X+�02�`?m<I�ĦtY��AY#�8��C�i���d1R����-A�t�G�A�Bq]���ҧ=��V����A\M�)��aZ.}�1!����ά��m�y�ܾNi��B��<���+�R��Q���dU��]s�P�'����~��AWS 0j�8�v�K�0	�������i�/��A����X���3�.����ծFHo�ɀ���L:��ݨ���ϾV"~��*
B���Dwb8�P}+cW@���6�Ωw/���.�\��9ˈ�&w7����R��nQќ�>����� ]��4�Tt_�^��$��ocq��X����m���
`~
pә��ףO�bY�b�/�����������7�wSC/��.��$��ǣl.��
P����%}>j	����1�-��r#wpo����O�c��E�
�_`�;�Й���^Sݛ)dq���(������N���9�<�?����O��ꍂ�,��!TJ݊�Cj$9]��Ip�$bg�Vi�z�Nէ�EБ�y�R������{�bo�*�'��Ye�cA�{�.2�A̧��X���4�s��� ��Vu��s�����:-�i�h�2/�˥�`������9�������#,���5��S	Ë��)ב{����~�u_��qRk6<^�,sA�3J8#�{* b��:�����5�=���vsve]wc�%��9�!?5��?�9�T�� g���/�6y���;�����P�f���jfR­��0Y�ʽ�k�ѡ�t�]�/�:���$�D��A��QJnC�}�+E=�
Z��8�fy�ϰ�]Iv��?�?�Od��t�FO?��Ԓ�G��đ�kz,vPk�p%������?/�պ�Bs�Ye�gJ���N�;�0�ud��#�����3�W��q���"�5q��_��$�x�b���=-V�Sl۾�|�����d}�C�x��Ѩ�8���'�Þ���� Rmj�,�B�?k�_���׃*�ЮF~��X�"�xH��<�x�5Um�i7�c�۹���_���7�o���3����&·��h�w
�t�]}^������O�d�E���8�	yp��4��A�� �`����6�(�i�/ˆ���X���ؾ��}���j�<v��ޑ1�r��p�x8Yk��'%�ޞ�PwߵgB{��Z	��;���%�4�1��j�6r��Иro&�ަ�h��ww��^��`j���v��fq�����7M����E�Z�$M�eH�k�Ċw������c���=��TR�S��EH�ub46�;�2�u
�?r���	z��9�B�Gx�R5c~�kZ'ӣ���0��+.P����g�]a%
V@�����s9���h�t�L��/ϤK��Zжa_P�x+u3;tO�3N̎��{�(aX��U��S�$A��z��U-~&��7��/�]�0,�8����!��F�%!3��թ��ŕ����w�����NzKG�N�YM�M����A�C̽)_ޓ�����DJbC����$)S[zk@	pJ.�rs%D���-��>!1�����A�z�;6�<B�ä  �֓����ry	�q缐�НX˫ ՜\ECN�������Q��dri�2{7�Z����̸玕+�ַj}�¹�4���cq���׼C����Κ�\֫�|h�@����M�����Xδ5�#.r�T�ȝcp1I�j`�th��:x�g���	�M�݉^nz5�P#��ryF�:h��|Z<Y����"��eP֝��w�_m��l�|>T�z�?�[�<0���F1¿!3�g�1E����E0��YǢ{��婘|��X�[6��8�S`���%;�~GH�=��C|w���%��C�-�wP��"Lj哅jX�ۢ� d?�s�S�g�z�3�=Q�j���Bk�.� �ʽ�u�sJ�ª��A�ZI�V�Ft,�l
�J)�v?Z��ݘ�s@8�Z?)b7L�1M��L���eܾOc������o17.<�^MN�`�ؔY1Pm���:cG��N��f�D��-a�p�T�tX��^R%�H\��N��0N�8����s92� ���s�y�F��6X�k��FAA-U��?s2�^;q�L3���R����!���`��;�݈eK/��s<Y�����F�M��H� ����^�mMq|��+�4��ǒ(z<*,Sݐj�ӭ����b:��v�D��T3P.��	e]!��A YJy(�=�	ve=:7а��!�G�]��Bd�,1�Mv(c~����N��M>eq�7��������2�+���^o�, %ڢ�~n	�`������VJ�a��)�J�_���P�Պm�Xq�S�� IΖ���\���M~�hXsn;�<�<��48]|$����A������g嶂$]��;àv�#���^�����M��)�|�������=5������T�V�{���c���p4������Ɲ�W�W�;�U��m� J���Jް�\���cp{�v��<�u���o}.J�+p���p��,]���:cDJ�-0-�5�o��!ᚖ1��!vJ"�����yn�n*�5����Y����`aCR>�����pf���ͥO&ݶ*�0�%�ɛa������c'�]���EP�����C�i����vl`.3u�f�cM��_��7���: hט�R�e�m5��f��Z�wXnf�,�TЍ���o���{��l�m�9d��R7?���k�����|p5��K�ﻩ��Dk]��|%��p�{�%E��|	4�+ƴn6���w[5����7ǧ�b��C����c:��#�z�n�X
�r����Z�/}�Zn8��]��G��g`�AgQ�I6�V�#��T�ԙ��%��V@%]N�e���]Ⱥ�xK�ځ��5X�54EXGX�m�|�	o��~=�l)_����>a�p�f��Z��2D�ia\\opQ�,�iǌk��vv�V�
�'�p w�xzR��$��o2��=���l���1��7e��k����:�@�ٗ����pb��ùvx�U#��֮�����{��]���fJ��������T�Y����f���x(�!����l,�i�f c_���Q�)�	 An�m�]
�, ʳ��;Ux�^w t2��_Nۋ8E&��P�\�P�,:�T���%�Q=�Q�-���s>�~w����(b:nGjE�}V��-��X\��ںbQU��ěl
�BAS��e�DB�b�~;���{F��>q�|[�T)4���ՀA��yX �OM �#cZv��@������L�(S�Ι�㿚l�͊р�e�=�����S1�� V� �9�=F��?�hC������lZ��c���C���[]*7A����4�5'�5�����+�&����`t]?���`���9.�-{�~�M��:�}ZM��k�j�A��.�Sy��v�p��?�Oѿ��y�Q7$���#a��;�b#��GV��x⃂Mk,�Y[.��t�����ѲO��1���kG&욋����ŗ8"l5K��CO&��@zP�0�u�-Y,/B�Z���0l鍦�����˗�V�a>Gڸ�K1��Eף���?/p����X��q�R�	�Pu�qP�D?�2��H�4X��x�l?�T'f������ (e��<�b"f�r�SJ ӄ�%q,klϑ�s��$nM���1E�VF|�/!�R�\���Ϳ�A�r�<��i����+���� ��N-����X���:����vY29a��j��Q*��-�,�@���G��	�1���ُt#�|�DT�ʣGMZ�'�wN���Ʊ�!�b��8�f1q �!1��Qs��Q�͢'p�gF�5�H4mʛ�5O��W,RI��"�G�����xC/v�µC��״��稱*���L����"�#���01��K��Cl�9�����r��;�œ*Ag�n)��d�6�����ĳk��y�;�l*���	�Ư%d#���y :~�����.�)����-�n����8S)p�:\��X�!Q���P�
�%z��)�6h�^�ۓ�-κ�[Y!^d��~���&�1(��>s��u�Q@���SX��D�B�<�*��T.�/�:����3w�'~�@�A1��j��U�g�7�;I�xN��?�s> ��[�7�������/�s~A>���P�r��W��U`aڕ_����Xc���]@��/h�Jg���W�(�V ���qJٿ(�v܌�Q#$z�w�H��0��ڻoM��efՙ�E�c��N�{c���h �F#���R)��X�+I�<�V~�(X'g{:h#n]�u��u��4g��ź��ډ�"@`�a?���KA���Q*w�����0���P»���7V��9�zX�J�|o#m��+M���?�
Y�I�ď̀Et����E2}���^�����ꨄ�|:m�(��\��Da�������&'T[�7He��2:�x� ���%��B<G�H�-�q��2w�P�с�ˎ�u�F���,����A� ��T���9�C�|�A�u&� r q#�q�a�SJ����E�����������}jT�'-�f"��K��'� q�a��,"L����3��gO�q��򘡻f?�!��^,g�8*�>��
	z�%H�+]$��A�� /$�X�V�>�X���R��9���bK��)}����.�d[b���9JZ�5��Ҁ��"*3��8D}KW�z s]1���Ki��m��v4���
T��X����zaw�r/���3�7������r�fV�O:d)�՘0%��W�~R~I�-�W2Fe&�<R!nXA|���jĝ."�Y�ɜ�$8��v�Kgݤ��3�*z҃����!u���G�
��jBM�g?Ȓ�>�(8
je��4m5oc�l����{����	qr� �S6� <���~�*%u�$VKNUW!�1C^|(�dv��wcC�~9��j�䯏ؓWm�o;�)�� 7(�:�!I~`Sx���t��V����p���jo�up���d B�rl.���$�`��L�۵�
����z�s!2l��(�'mod�������oI��6��I�i$�<��$�i��w7�S�;��r�C}ɡ>9�]oW1�R�P@�%��%&�'2	4��mu�����5�\k�~��u����J��~���k9��X	 ���&�B)	`M�c�&������Ň-��9�:2Ɣ���6�p ��ҟ!��6�� ��oY*>5ܥ�3�y�2�G?���&P�����M�BI��)~�Ⱳڔ�V�mA���y���Nͥ����o�.m� �����
��Uz�#�3���UJcΏu!��f{�y(J�H1��I�Xn�z�Lu.V�L8�GU�b��8� ~@�k���8-�������%z�c+���؈z$����$ɖ<�N��>NJ��vs�>0��Kaf�][�i@��<#�Ru�l֥:μ���<T�����2������p�x��iՂ���P��%j66���R�������&#Rxu&�0��QF�G�'+c��Y���Yϧ�Vٿr�F� ��s��OГ[��vQ�����3�<�2h{��v"S2e^�JO��Le_#�	v��:V�@x��^�d�e�3�ww�Z؊bp�[��#���@6�N�g��c�m��jD&�cJ��i�A(=�4 4B-�с�hm�C�t�3e��E�Sѫ�	k��"4��0X&��0N/L�M�J�4��!�_���c��i�p���[�����@�~�zއĴ�����?<
���R��d�&�a�@��-s�C\�� +�0�{	�0	9��������쑙 �?͑�y�5�3�92�aq�j�E/��k_rf1��xT\���E-�i����~5�ߐ(��/1rb?��$�3H��
�`8� j�gMU�V��X�c �����?'�ډq�L�
�.��70%s��,H���S�ا�E���ڿ�ux���&L�-�XI���\�oX�IÎ������f�U���l�,Z��$���1�&�~t�IX�)�" 	��U	p�n���ےxn l;��f�`*?	���Z]���"Ř3���Σ�s�+?�ߔׁ���GC�X���H�N�'h��o}@>I��@v����T�?:/���_t�6����&�b���p�w��(3���rF���\7����cZ�]��yߚrl�������^%���>ꇪ��>\�iW�n<־����-B�����E�GEȘ=)�Y�<����g��<�����A�gp%kh���;�8���������9`&� )�f!� �V)C����>�Q������ق��+���mk���:�fx�H�.h]�u�/�t֘�q`�[�F`_D����?�3�$��ԉ�)���u�>�%ƚ��pdds:^��z��|c"D��x�4��'����
j��5�rl=�He�Yn�RkEQ�O2`/~E�p��F\�6��	��/9�z�@�G�{E�eљ��j���i��{������Rjh��w��9W�EC�*e���AO��v�)_����?�fk�;^���e�H��&�Bk��y�YRй���	gkm�Lq��V�����zHKڈ�ڌ5��~H�K`������(��`�O�������4m#�o՗h�-��,c�jQ�n�7�˦W�Α9)�w��(į0�q,.n�X�t}' ��X�2D���纬<ʼ�`�ޖ>*��*0� ��D#�;���Be)V�pM++��l�Gi-��A"&n.ĥO#��(�T!x�!:���@s�q�.�4O��S�xc��`Wy.N@�'��y�Y�X�M��ޤLՌ8�t���+#�{����n���~�>��B��F�z8^�&������������0�j��f�w�XQv���~��]5&��~�� A�Yۙe_�j��i� vԷ�~&6�jNA�#������Je���I�����Y�gQ� ���A���l&;vV��	(wc]�rj"W8���
��k��]�>q<��o	0���8��Dq�+��v͐9ꈀ���}����l�ϒoc�ʞ;-3���vv���,-��Ԁ�ƂY֘ X}r(�@�|eg��S<;�5�����a'����!��t~NRS��$3�é��2o4����w�!�-O>�|ZWИW�'<p���ؐ�%�X����IW��G0}U��QNĒ�XS����7�c��wڽ��+�<4��}6��l��ߡ�P&�tƧ���B��֑�Zo�\T"��"��鰄t_kkh��XA�����D��䲬��m�j|��B���p�������^��E%$"?�#��聖h��Z��F!�Q��5����(�i$@sk���E	�Z��#�������
8�M/�$zdK��M��Y6���֢���:��%F���,�֦K,3���E69�ſ6És�0���[s��fn�f~�"fS��;��nUև[$כ�R�خ�� 䆫[�9����n�4_}�|��8�T�:�6% i<*xe���s,�Z�����pZ����܌#�YX�����7g�ra�<�������ǀ��d��N�p+���P;,�7�p��/���H,�ʊ�y�@)-�͸M��4^����G�{�N����2�~"!�V)��\+��gh2�5 fy���ɢJ���ibN��W�{FSY1�Ũq��xb���_΍�PG���홓G]������;]ܟ"�cd���,�O�e��ƙ��^�<�W�B��0K�@�I�\6xZ�(Ƣ�ˮ��=Y���� 9�XJ�	E���$qX�	����(_�r�$�s/��^#p�jg�=�������K#y1b�%�����P�z|Rz��~��.�zJTp(����XS߄	�S���B\O3�H	v���B��_�����LF��E�����~�p��ș���ȵ�u��)��L/t ����殶Z�M�p���8a�W���!��}\��6�W%m�r1�ȥ_5dN��I3�}��v�4,�����۪�p[giٰaEw�{�	ФPd��Vxr9S�UJ�� �x����49�E�~S{�mG�9���O:�Mi� ���x�LILk&6��!-�s�3�rj������ȉ�⺙�c�6�Jb������C�����t���Z�o���98�<%d��|�y_I������S�Y�-U���#w>+#Hϟtc�e��]��sF��#܍�7�g�����p��oq0��>��/{�J�c�`�"�oTWh���տ[�\�������i'̸�+�k���h.dx��͋���-��Ug�N$�����X�к�Y<��!�.`��Se��z��7J�]��T��'�8�L��`V���jzk�&�8s��,�MfM�y�$op�\s��GT$G�� ��s����I2�s-WY�l�o&1q���v�p�b͆Iu��g���gJW=�>�Z!
��S)��(���vg��K�^X-}�����Vv W`���%�$�������2.����Z��}Q�dk�ͯ�(k����",څNx E9�w@�y3��뮧V�sֶw����>���R?C��I��(gH��;n�����y��z�x~�0��.�IR�߾[���d�S�Q�i_�h:�>�V�,�a|��q�Vp��ަ�E$?==t���z�̶'��̝��ބ�f�/�.��M�zFݕ�sH�\���	�4�s�U"u$�e�Ӥ~6\\�+U��-�+~�6e�t����VD����aڲd�;K�1]�)�JLz�B+'X֥�*��)��o-ޱ�n��c)�דi�Cϻ��ŝ�3A�FkZ�)�S��`΋Ww�����g�0+!uw���oz���E���Q���lPz!��D�0�b6�j/6�		$y��L�.>�b쐠5X3��3�	��+u�9|�����v��\��S+��u�yt�!W���rF���pt�RU�Y�d+.��Vyp�A�	a��*����Ǳ�b��r��H�vB��`C���}>��b	�nNa ql��Xވ k����{�J:u��UrZ�0O�G���� �ч�&,���AcD��3�8���K��]KmF#}2���G�7}|U�0�,���5�S+1����x��,}E�*�ҡ��yy����gt�#�0��d2�F�9�4�=!�?`C�� �u������BaH��e�A���)࿞0a�_��	���MC�nf�C��a���5��~�����q^��1u�D�r���!��g��w�m=�螦D6Yh#�a��������>�-���K�ϥ.��F��h�MQPupԲ0�����{:ST�_��
���A���T�*�ziNЁ��n�J�M�>*��ń&E���p���mͩ��e��&V<?]�}R�l�������-]"b�@�Z�
2�Tv���1�:t����ф8���]�	h��B�}�/��JD�w.B�h%͵{s���ZՙtZ���7�N��7@hwE*����Y�A,�x4���t��x.�z��4g<p�$</0Ǡ�eZ��i��{����:�772��.؍c��-�Ay���>*�[�9t�ԉOk��U=��k�*��4Ě-ܰ�X���y,�F�D4�4-���Tѯ���U(Y8�H��O����#Vل��x��N�Q��
k���߼Q�*�!��'�YGQ�tN�Z��V�Gz��V�}�1u�Air��Ry�L�����ŪB�Y�.*$MdCS.L�_�ӊj��*�n,\��W���2��da�I(�ќ�B-��ی�J&�K��ȋ�����>��/w�e}��6� <� H��Ҩ�	ur)�|A ��B��a�oV�O �Yv]���Ǽ�G

��+'\����v�y��*R^zzR4�b��x7'.�
Iu;�}j�Pj��>��o4�9��<-�E�H'�vZꅼb�C��8��[�b:�Q!��Z��:%��	�vFe,�j.�ߔ���1�d�	����!Q+YϞ��j!�H;�P�u��A�����uP�T�ZcL��vKU����ez{+�,�/*��g��9���;D�0[N���#li+��/J��������"G��<�#{[��Ù�c�T�2�5�T����H��R�K�Ʌ"{Rk� ����/���%���Ey{����C���b��Q����l��Ft7�S�Pɚ(�����}SW����;��xtb�Y��;$���}�)�9\t�X.RC2��:��N�[)p�*�.x��"�!���i���)ϛr���b��7�#��is@)˳|�k�e.X��R�A��)A��eC���*�y��+�wK�լ���++��*�Q��XK���$��U7��T�/D�댧��ܣ�@A����/��@]�aC�FF��p�W�����~擴Pjv�����!�!0��)��>�|��MG"�����ٕ�@�e�
S�!�W3��P;���i��O���6v{��$��k���9C�M���.g?��0<d:�ʦ��xZ"�0��o�@t�e��W���I�W0�WZi�����eS��p�V��k�f���Pv5Gi߰c�@��'P�J��]y����1�)�2�glI?g�*��&��˲L`���*4�Pκ��y��"0`+����Cm.ң+�Q�l2�ÒR�{};��'��l7F��3�uq�fF�L@�h��`�Uz�=kW�{�O�0j!I���=Z¡~e��q=#�;�^���o�܏�ɕ�*��w��A����<��=��Xї�O��	I�Eٔ�+��7*r>�(�d�ZUO��/�%���1�l�Q�n*����ɉ�j`s�ř�b��*gI�dN~���{d�͆�m�4��܁��I�}��@�q�ݡ�(A���Ԁ/�/����UPO�4O �h	�K��\���k+0��ә��o� �V�!��<)}Eh���_U�]l�͇?M��p�rT��ށ���Y�����3� ���+��'�.��PS=��e�rV|���}�g��G�Zh�m Y6�lJ�TA�i���
�;~r��X����C`�[�W��0�=��c��Q��^�A-$y>�0#��sYUG���Fg�GvB�Y��*{���\���e�����ȏ�И���sG����-J�Γ�Dc���`��Z��N��0�`����sPzC��T����#}� �u��~����҆�-9��[B� XK%+������ #�*�O��p����"�-G��~�毼ۏ��%�A�E~� �} AYo󍚈���څIV�o"=�T� ���>£��@WF8�ç�^0K�e3���Ҋ��G��(�Α͕���υ�T-�ؽ�@�%����+J��|��_�|���^�
��O���;LfW���,�R5-E�:Tp�,ꜱfXPG�i��s,�����{wR�8�5�S4��t,�oX�lj��0�LvPY�x���t�N�`&��\-�sct�M�S`�5�0�}A� �`9�p1
��y9;�b(�EQ�~�$۶c4�n3��wpmoZ�v���VL=}�v`�0v?!�V���gK<�(���N�@�"�/:�Yc�����4���f�����Xu`km���+�����Hx%�ѠB�f��_L6P�8����(��M
���^a���v�/�z����(	����Ý�. zN��z�r�yK�ɀ:��c�3��L9��=��xz��l����"��N�[
�l�/��I�3�����ڀ��~s�^yp�6����mI}��,�����u�2����ߪb��P�q%a<ї-�{�Ƽ?~��|��Oo
���h��=t:Q��	ƨ���C�V��e@X�}�s��3Ӄ>4ß��b=�������#��/.������#TEƝ�|��?R}���QO�t�z �n�ț��ic�v�%s,�w�~S}k�8���U�B�p��Q76���ShZk�<G�`�7M�=l�ID7�l�^�:Yq�P�)������#�*(�E�u4��-�!ޘ��Y!������8������N�&Dmh�B��!�@�%e�a �%�� �۶sa
b��!���C~t7�����v�	�]�Q:-^�u&�j�}������s��i}�O��7�����Hn�2���r�p�Q��z��ռ�Q��}	�5Ņڕ�p�d7�� ۹J9D̱@�B�
��Ft�l.&�%�X��#�ɚ��Sj��z_�q.�AI��/2 �إ����pYO�&�f%)H���HL��Go�ǶGe�[����'�̿;�pV�Glg�0!��9�n	�ņ�z�bu��ٗ�{��+ d7V�Ŀd.6���I����>T�~�<��8��*o#�a)�a{QR9�ɽʏϩp4�*�z�U$l�xv��{WK��B;�b�A��}T]�gpB#s�ynzpGV��|n�
�Xu�8�ir'�CR⿬�-�p�����y�˭�8�LsRE&֎��{�4���$��kДnZ"�ГbH��X�M��ז�j�YT��,����Rԁ�X{xV����70Q���y�i���&�t^E���ͺ�x/C�Q�E�I�ח}»�����ZS��s|�����D�O��{<���m>+�_�?ŭz'�Z����'��ZtTQ�(�n�Z�A�smV,���X�Q+�"3���d�#��*ήҷ�'B1��˾�����VF�uJ�Z�����?h)�LҠQ�"yݒ�H=��XÅ7_̃���s���A'���C>b�$*<L~F\B{����ծ`Ȩ�2��>7҉S��
B1b�3i<�u��k��^�Cg�ҧ�3�#�K�f�E�����}�9�~&�������B,�h>�¥�Q b-sP�ml�1���3�3j����Y��Xp��?Θ�d��ݚƓ=��"߶fpw,�(v�L����IFn?��"!�t���%y�N�ݲ�F�܋��� �.&��߶\i� ��L��m�5ͧB4}t��Uh�ݱ��jz�4��3]����`��>���-k����6�����d׉ʰpq/sd<�	c�����&.$]h!^���'�х_��ʶ��x~�Jѧ7�y�p߄�{҄B��;��^ |O�rD?z��|=&Wl�a�}�{�.�dd���C{&��GL�k��6�&B	�7(1�]@n���D���N��L�Héw�ۗH֡��|$b��Ow.b��Kmo	%�ߴarڌGTK���jzn��ٖ�]�V��[Y�]QE�3S��W|M���|��ґ{������{�+P����|�Q��hN�կ�@�%�l�O1������՝�e�mh�a.�h;�3F�dV�:C�k^g9���9l����R�a��Kfz���+z��H~�����,6����LF@�{h�H߸:ǉ�C��߀�!^|`S���vna:��a�j�+�.#~{*(���K��Z�a�U��:��-`�ח��w �ߢJ��FV� �x�;��u ���3x����A�"��Q�s�Bx����tB�jH;��y9���uE����C�V�W�nLŕ&����������2��?w̕��7rW���E��u��-��΅w�~��:��7F�5�U4�g�����m��d���.!��D�4��T>Y0�'�$G�	G�v�3�n��\���w(ř�A7��F	����;��[�Cr,���B��g���~VQ.t���t��5���sg�~_r�G{[���m�|Պ`�ۭ�}�ɶk�ʐ�6�r�k#��a���>��U�W�7�&����e���Y�YUkΨ-��{��j��!詵'�nD3gt�9	E�zoX����\Dڒ���}q�����!�x�4Yo�67���Z�����;������0N|:�����57i��������q<��ï�&�Tg^��|֔�Rl �I�1���!f]:J��؈ObDM'��h���e���(RS�ۿ/��Jgxs��:Ltj�7T߲8����C����*�9��H�!�� ��/���Ք�t�{1p���ʘT�����`�����aS�I��
H��L����A*�C`Lfx��5:�5����آ@�>��2p��ϖ����b��X6X+Rڧ���j���C�tj�$�7&�7f�� �џX`��I��@B�U�INl*ץ�D
`_��)?�����}�433�EBɎC'R���wx�߅R)��v1�&�p9n`h�A�^S1��5E�E��8D"!���>(�p�*磊�I4S6�K��i4��4{�]y2	�b8BLi B��%�>p�26g?3��'�RU��"<o����E�-�5ww��^��6����҂^��Ib�N�C��&r�m-�|��Y�
L����� Xy��?9'��ϩ��d̢����km���ǣ�^���]��E���Tz�{��;{:ni`�{�=�����v�&�_@��	|�ݲ�^��D"k��&����c�h�]���V�'BDZ��q]	yخ��</+<��S`��
�W
.�#0�?�� ��˖:V̼v�����FNe2�W�7���2���&�����&��b]�ps��ip K���b��.�{r���j�m�f�g�.s�j�	ش{r�+X��i���&쥄E@�x�M䥝1ۼa�'�)�������?�׉&��M��Z(���|�i�7;����	�f�*TB-錄di�"�ʃ����i�q[��S4 ��hmkL,���-T��n����#�3*�1�\��P��\�V@Va�w�U�h���%�){�?���#�yX���Z]Z�4���*jWǏN��	�ջ�1!u����֊9����68v�s�k��)~�ͲIκ(����m>�d��ܘz�Y��� 3�-����<�8��z�E�o�%����j�!��m2v��f���诨��AB�Q�$tOq��g��p�ow�Ԗ%�\��6i"q��X� e
�����*�����[ =`�g--��J���xKUD}~��u�J���wO����`��6*��b+狤ÿ��{h���v�&��v�����Yy�x�=7�ШX[6}�ݣ�1|*cÕ�&��d�`�\����n<A8J��$����-�K6É��^"bP��"�]%�L/:@T
�#	�g�=o~mZ;t�n�ٓ] Y���ߐY��$/�j��3�_"�?5�:[��Y[�"�+�)BN��տ0��JLn`��$I�eM����.Z���%�QY����l����yuXW ��T
��%|u[��?��J�Z���ύ7&�
�YJ/�3+'�ɿt`{�%�v|}&e�{�d�����5NZ�|��
�,q�z��3A�e�UX7F�j0��F���߽��JΆS�GSlL�����=���o�
��%�t�^(�PP� <F��]ԑ��*t?U?�8�T&�8�N��TLf�&��9��4OLB*��:�����#���=������V��y%*�)��m��8F~���n�!|W� ��vmM�@�S������Q67�M�pod�)�Ԧ�~"�t�}��b�����!���2;b�%;�����(�/�6P�}���/[��!ȇ�1i�X2�">�g�g�����ʄ��i!�bm������p(�����8T��ҩ��cLX���'�_��밆�7�lU��n/f���qV���x�6��)�(٨>&-�}a5v��\�d���|�}��$��[��ޢ]���{ �����r����[��~	��R<���NQD�-6�����&A$#���v���8tZ�I�C�Ô�e}O��PQк�A'��ע��%�W�Ε���H���YL���~N�L;�L|���50N^�ϻ�)�P@p>ߙ~�Ű|~�-�~\�-�v�r�B����2
�o�(͓�iq��x�+"�w�Xך�Ss���,!"�����dG[@� ���,|�RuגRiK+cu�+�0I,��~�׉��[�ӑ�U�(F5Xt>�����:��W)��eR�^Ў��4�t�3�ҹ&Dɢ�Rt['A��B�h�N'G]����c���>�[F���wH��0XÜP!����,����reҖ���M��x����v�N4c0���$`����X1���'�0�EwU�)�9A����j����>�J�!A�ND�ϔ3��ƙm`
�E�l~�L�B42~_�h+$*NåB�"5uW�M|��$��ҝ�%zҁ�휚�K�V �j���c��;Tǘ���V��3k=*cP�r�궶�K3�<p$�� �/�AO��}�E��m?��+��CN�1�x�Џ=aGFD��:x���Ex����K��2�H[ܹND�tzC+H�4��􅩀8t�`vЙ���wV�4x�ƣ�RLf��s%�����6Տ���'�kn-��ND�v���rg�+�\G�c��eݲ��׃��ii�N��n�~��_ϪǗ��Q��(�K����q�p���J��{�:>̵
;@�5$3��\�����r�_�}�ݓ��P#(�4߁���HT��B���S9����<��d1{���$v�+G�b���J�x$��nB3f����G8��i�
��nA�s@�1]�-���lE+`��%v�-�d�A���Z�%W뚇�@�,0��<��������-]*�G������go{rğ%�l]�T���v���x�����+�Ԉ��M��^6|��A��,M��FbU�a�%3��8캍�ǥ��%6���s����������V�rEz�ᒛ�����V���zB[$�Y'w�ٳ~�J�E�+{)}bdb�u�NO��������E]H'-�htYT�-�����	��>���c��*��ö=�u��oB�3tK^�Б}��\�i�,.V埙3﨣�#e5���c���6Oۼ��&8<D�A(v�v��К�d��H8���S唗{y����h�A�V��At+�4T�L�)�.�A:��%�\��ԞƖ�j��vlI�'��['�����e�\�=�#�x����^�Ϧ���b�6�к�������vf>2._q��u����a�F�#�ՀCp�_z7��F�����o�u���ǡIhZ�-`&u줟��Mgd�j+�Խ����>n��g�z�����x�U����'%��r�a rv�*�Т�\�6���í��rO9�AĵQE��+��R�Ӎ���p�|L~��I�_)RD�՝��ϲԓ/���-(�I\�:�7Ϯ2z�����[�Q�6�����$��G����M��o���D7���5��^rN#�΁��)g��{��V�⎜��Uެ���U^�@��&�Shy���2�pNB��)������X4�p ?�FK�J��3��jc%�Yk��Sm�/ʜ¦�/�A�ɹ�T�R?AO�n��(�ux�;KP�eա3���;���A��M�Kyo�D��w̷�:�Do�|�S?��6��x�Pq�"Ъ�'g�Y�ܤ��z5+���G��C�Ih���������pBBD;�q>?��Ṑa��&�+G�;9��\\3X�M(�Q��T����F_ |i~�P=�����R砿�#ٹ���T`qs�9�|�!���,wx&f��a���b�����"��\ɕ؏w�BD�k^��eɍӓh�K7=���<�ȝ�<�X�lj?�����B�x�+��+SnƔ��~ȹ+���(�����7�Z���-��{���^��B�,�睵��l�&>�9����<�U��y8�n�FR�{`B�ѝh�
(J%6��dtt���
��)N��[FMB�i���E̥e�G�)fɱ�'�¿5wʣ7c,��<��#
�� 7?�p��o�=��r)od[����ꃧ�#8^�k�S�F���fU��,&��og�ԧ����N��vi�a �|Nl��(�I�y��ZtE�ȍ;.۔�:� ��"�\�k��$�*vçU�����g�#?���V}��O������(�K�ʌd�H�MܯU��OE2Nh;j����)uVK���'`��v	:���NF����'���7�s���BAS�\(�s$v5�M����X�gYuI
��+��\v_�	�d��ȿ��J�G�������8H����U���¥b	�M)� �#�8��u�H[fÿ��}�!�3�8��Ң�u���N�@Oh�x�ι��xk/	3�3�]�2��Q�*��W��Q1�l���{y�[����Ȩ������PX�e�:�2ۜ��n�Y������y s}�W3N�q�'+I\G���q����el�°�T�@��y�-��H��O{�z!�e�V��pYE�������(�������F�1[��gW�� ����i��:�0�{Oa��a�c\��ϵ1.�����	��3�s���+�4���p����i'��6 ⟞��r�����_��O����T����q��1dń[%���"�lZ��>�ub�[~[vD�D���^N�6�4���H�#$v��~�K�b����<��Gh����
rr(�U��7��w|i����#��K�Ôߟ���=�yB�����-K�{���.�\�)S�"�I�2��ᛥ��X3���גz���ߖ���5h�H���jge@��w*t�5h��.X���Q��;�k��u��k`wD_d�BP̔��0:��}�9[}@l|�`���h�z9�s��H�͑�;���MhGf`�w�N��;3cke���F��*d�F �+��'��"6bs^ȩy����FH��nIFQu�T�9��Z����Nϼ�P�\MMt9�B��<|�a��7�UP�:C�yc�u��{Ƙe�`7��ir�+���H4Q�R��h�U� 9b}Ǘ�mØ	n��ʻ��A���p��!�N�;�_�P������@utU�j#�C��5�܊ǄAo���f�^��5�P�7I��B��G����i�v���ڤ� �E$���tXw�n;��ڼ=g�(�MTN��wEZm׀6�i��@
4H�b�:���V�� �������
HT�ms�/�Ɂ6-�`����(�K�J�H����9�)����s�U�����HN�M�^[�������<
٨A!�P r��1��Fs֮o<�N.yE�K�R�j ˖�zLo��������̛О�;�)���)B#�.}���("PQ��q���5�A�#ܩ�ob�N��o�a%�$z���|Y��cntV�#c���T.�j�7�-V��-\K�0�������m	&��;����ڞ������"�v/j���~�~\5��^����䲛DB�A�c���`
�����WZB�[O�����Z�l��'<hQ� ��X���(Ȯ�©,���n p����~����5��Ą��^D�$/�O���M�dDp|���6Y��2ԑѯ?_�8�}�!�?v�d�Y7�9�3�d�LRƔ!����Z�m��Oy]��=r�WS�/�V(�'�-pv�ݽ�U���f$�mL�V����|���)�-�b����� q��d�i_H�H�x�>�=�T�d;����k�����f�p�����rZ���qB��g�ʺ�(���k} ��m��֣ܽ܏�=S�_n��G��%�I]�`�l�:�֩��J�<�_#�Xo7��eL�k�,��'��ĭ��Euu�S�;���ԇa�H�_ �N�[1G���b�'i�bQr`�[�GrM�� �]p�G���m�	N-ME�T>R���?�gy�ف"�O~4�S�X����g����fa�)�^�f5��7$V��É&�$c�-�|���I_�)W���tlU<���~�I�R��+ߌ�[��t�?8�J��э�4�{Q%�ݜ:�O���	�J0I3���N	�UY"��3xɜ�f�V
�߹'���D.$�J�3KF�&�@&B̩t�iD�7�L�.��������r��E^Β�%�N���q� )� ���+x�"~_�ϻ/ք�aL�?߭�p�]�٫���xGh�3���u^s�~������+�����9M�/I`���Fm}�#/>")�M��-z�	�d��d���zc=�'i�C&qR�����:̜J�OX�?5���|˘k(�` ��D^�T7����+��O
���9�*�J�<�'�'rW4�l�5�W=�_�{��r�	�Q�0����<�� "���4�#Ae<Ж��C���w͙K/����7d�5�%"��H^m*eP���9�C�����_���8�=���8=���$z����]�1��j�E�z6̍`�r���wL���U�����N�,s���@��C���s⑉Iϒ�QCn+�V> B��TJ�A�/��mU��^��Eۇ��b4�8�^��xj��5�'cأ89�%���Ȫ�SÚ�Ңw�	8��ۭ�� ���Ǵ������rZk/�iS���P������gsp.5��H$��90�D}�V� i(;��£��g=����٢%�&�|N��ū����"������ˮ���6m�4N��7�Ĉ�)��/в�ĝ��7vQh�縅�q~ο�����.ŉu9��k2y_�G��j��V�h9Y❉:#�+��t�`K4��((ps�,SL萤����i0;Խ4L�w��?z�4ULu�N�~⴫�Q���@y�	zլ| ��i�N����2��W{�k�و�n��<�G��тI��f�ڍ)X�{0�1����9��o���_���k�s$j�;9?uѰ������ҹ�?��r&��oȧ
!��<�1�q ;�W٥hga ��$�̘|���);���5KK�R[/JfV��g�����o���m=7.b��0:|����[-� C��է
� �%���l�+T{��W=��*w��vy�[1�b�'C�5jI���e!��`\!J��{5w��.��b�j����[�ZQ�b����e�N����P���S TGa2m��DV�J`e��zֳ�L�����}n�"��ŷ��f8bJ��cY[;?,'p�t�4��^Ŭ��1�`�G���1�BW�i	���a�i�iע.����� �<z�p?��w�Ff%��m&�/H'H3~�r0�:S��D�C�@�P�@ί�'k�f���	��;N��٬��u> h�L�%C:O�V�]� �ej$	w�X�9�I�Y�	�{����I��a5*�S_�^�@_�Opw�Z`L��~�Z7j]�U�)��<?�!:3�(Н����3h�YN	%q��p��% �ͥ��6],������&�z�L��&�˭-�M_l��q󫍠����XT� 5�[��I����𔖘9N5o�rI09zAq��ِ\Nr��$q���ik��iA�ujɉ���3����Q����;�!�o=e�q��>5`8�;G���V���0�vd���+�*w�i�*W��RE�z��-���4D�<�������B����o���5�2�q��w'[=N����`�7� � ��*T���v�ߦ���݀%��L��ՙ>��Ń��4�c׽�n9��py ����<�Ʊ(uprS���?�!�H����NμzQ]�O�N���������w�O'�K����$6'�w�p�M�lڻ(f�����O����Q�����I����ÀDp�S��#�d�2Ŝ�M��+�Pn���~�E�����l��y�R��8',�T���Չjm(yX�.ZQa��S^�j��s�Q}�]���x�\-�0���E��c�JK�$�]ש_X��h"�*����5�&_d�
{6��,�5)7�%��*dZמB���Ә��ʜ=������L��ٮ�����ѳ�K�v� 35qg"�"U	f=�P�^L��ڔ!L�f�n�P��_���IR5Z�E�r��ކ�x:h�l��1���p�
�x=�����]&w��}՟|��|�����r���Q|��U�ϓe��Y�}���:[.J/�j_.��a�?��V�8�)�u��M	$���L{��FV���̬���$��9珬�ޢ���Fǧ��~��*�R�a�q�nsY�Ŵ��C�Q.��T9���'?�,6z�9���/l���"�����q���E�Y~�H	q�[G",���PQ�*����%I�=$R�����w2K�4R�S��`UA����!��v,�(�y�L�9��ꃚ˯<�7~�@5��W�X�r	������0�j��yppԛ�B��P�Ӱ)iM��p�`�{(@�!�]�׺go��$����f> ��]{V:6��'3+��B�,v��̴�S�?�CڽE�D/��7���߀ۋyB�eؕkU�Jˉ�,����"}���jS���Ԋ R��
��6���-�n ^�Y#��BD���]�����$�Uk��a��V�W�r����$;>���>u?�G"��:-��A\oބ�z�����t[�LӬ)^��ﶍ ͊{gu����O%�\��C� �{s ��"fv��l����#��nG����Ų����d�PϬ�:�q�r�� ��*"%�*�[PP�Uі��1b$�5{G�,�ƞ����0�6�O�2��p�X���Y�?��@�R��,�A��؃y�1��4'Mů� ��y�Y�[�[}?ưQo�`�w&t'M��PRs@qǣ�zޯ����L'�����?+؛~n��I�E�CKJb[�qCs�	0 ��QE�گA@K\�=m�B�Taoh�)���_�����>�rR|�h?��ƞu��l�1����<]j5���	��7�S�|�y�R��#ydA���J��@Om�H����=Ƃ��T*��V��u;[��ؔW!qޣnm��qʸՇ���=CTJ�K�>v���K_i��fW5X�hj4����0U��W����(.���,ޗ
�;�S1,l�T��R6S�[��;���"JF���HV/�I������ˮ�-��s+'=e�+L�C�������W�T&l�Sﭘ�Q���@��/4.�)��Ub��3��A~�9���  x���F�{�*ecjX[?L��~��5�G���4��;wd|�$_ؙ��6_N�8��P�Gù�G[�y�/�/ߵ �S��/
2h���n�AJo�MMk�M����d!r�3��n.��u�	R�vK�CY������s�g��7Q��đLM��sK�|����|d@�/�j��_R�r���.�g���u7{��X�l��b�<*εJ^���^I�W�0�)=��q�cۏ��U�4J�����k��6��%���
r`�_�g� �͜�f��f�7�1P&��q�����űGl+�2�_�t%!��O��*�L�,Oο ��UD �y�֠q�#���&A��g�I!��	o��� �b�x�N�\�/s�ZC3��fQ𻸘�~��&�]y�m��u![�'�ǫz��kʯ�]�G�8�*����:����|�ʙ�"�1�/��E�ʟdʮ*/fct41t`�gp�vy�9f�PIM��T̕����]!�lK)C4~H��g`P��je��B�Nj����u&^�cz�P&�WSa�p�$��U~u��E�*��
ðTe�'�5�d�������wqG��?�ȥ��D@J}���?���������i��K�� E�Qb���غ�qS��u����|�5Q�d��I.����6�vIDo�n�f�qRXY'�c�I���>��*�ʵ��ƅ_��W�f'τ���:'�E!N�HE��
aO��͉��-��Q�Ӏ^��z�s���,� � �>�W̸���E&�^�>'ߞ� ��xἬ���8�W{�9Kapv0�X�䩤��p׫�Ź5%��4y�2�PJ3��o��u	��������!^�m�1������YŊ�YD{��Ҥ�xƄ��^f�%\������>]�x���v���W����?�?�����Eb�Ӽ�M�CC�D�L���d��$�s��r�tξ�*T�J��N:n��ҽ���*k�6�&�d��o�h�Z��#�@��t�g��XїZu� ��e#����w&���j�&�M>�a�ΆD�rΣ�i,�!Ql͘����Krv���Rfm-G���e�
Y�0���M���U�iJ�[�-љlm�j�%H���-��&��GU��AhN��~P|��aB���ͭ�l���pՎBWXf3���,�P8��O����>yQ�R4XQ��/੿��?\��#�������_��o"����Y=rC�=V�<MN���T	�	%w�¬�̹�~g�P�W[#��a$��;�D\��0};������S'�/;��l�i���~��H�`$f��!e�x��Ώm��ĸǿ���5���Z��*k���1�0�0"w�
,r���$����vh�)����4f�gE�`������8�M4X] ��Y�?��H�+kS�S�����.8H BsY����kd6�ؾ���Jl��l�L�ˮ�{m��lGcQ�3w��j��XV/�*�.+]m��9��d�0l�K��r}9��=q��.F��+	�9+�A� 2���ܜ6��]�w��L��h�����L^�ۊ"I�kv��X�K��`�&�3W���>V����&b*������ϽU|�Q���@�N���|M��ֱ���RH��W�a�Zv�P�^K�<����UH���]�h^z���λ���9���0nr��g�,��R�Јo�K��<u��Xp��>myb@e���=^HA���E'G:�jT�n�����v�VW��؎�-�;b>�)vŢ���~�BL=��P�i�r!]��`Q�5!?Q�����}�<.Z��kE- ��1��;. /���N.���zfP-.�K�D[M��9B>�*�!W��\�P ���Ī���e�^jq��H� ��Y�%0��]L&���?�8@C�*����`I�.�,b��C��>�Kx+�t�L�����E
k�Y�JC�L$���X�#k�Sw�]u�v*&ecηE]�/��Q�́6�2���Z-,�Ӿ2r5En�I�y��pm��`�W��-w:''��NH&Y�`;wM V_\J����w��Q#)�'�q�8�g."�yL
ʹ�Sb�po[vA2#*j#M��o�σ�p GOS@�_vӻ�"|�Zc5����l�8�ɋ�?�Ƣto�E��.dm+�޸Q���	S���ȩ�fv�J�����Kc�6���J�MM��Ӛ�ޣ�D�?�<����v�O�M�FF�m�����un(�&��%�De_�#w"-�!O,� ��r#ش�J�J�&�Є{C�<�g�����"@8�`��Q�w�ɍȘ$���Σup{�PV!%���������>^������t��{�� ��4�'٣'i�����?���]��C?��!����{��QDѐ �b<q��:��>�[�_�`��_����4W(5�w�D�cȺ���n�R6�,�GA"d7��ȳ�qv�n"�p��E ��������u��C�5H`�a�*e0k��cط�� �����������1C�6����;	����^�Zl^�s(�`��'����t<:�ږ�>QBx--ư�a&^F#���o�����_�%؝�{�^!�:����[A����n�G� f�@r�+�"/�n����p~
�'�k��ccN���iX� ��dB�Wg|���~6"�*�,����$q�l�s^�%���s���qO�J�cND�j� ��l^B�	FA��(xl0�dv�r��E�h��{+��x����rI(�<���$de\@�@�M~�MǴNv��(^8Gg�̯��|b���u-'�~K:%>D�i}X�V�H��q��0�C���R�� ,0R�컇�;S�2E����^�J+��="���_p{�C��q ��<�ƺ��#PD��>Ag�&�8N�ٺLK����]����j4�(�Fa\at��n�T���3b��{��?WAf�%�A�@�Ä��V.�a$uΒ`��N�b����+Ԣ��JT�e���hO�s�J���f���!��"En��A�,�s�>�""��~<!u���綵�b���4�|P(ct�M�bM�ň�V��*~tY���B�3������I�	�%��h^�*x�N�9�n]��]���t�����׵���������л�IR�ڦ��;),�?m�є��T����TZ���Ut�t4m�	e3��y�;�1�3Xu�\	Q�{J6�؋fm����q�/;V�J�!^�?U>�=A��3�sR��-=�!���5�jz_��%�!IK��_Wz)��~+]|���-�s���@�pm��$�D�rn���)�G���];4�h����;"���g�KV�� �]��D& ]�$��HP�e~���<g$����l2i�N!�@1xr�|�����mt�βǬ�!�jV|�H�L�u&j r�(��8��ncЮ7�Px#��띖G�+Œi��׿L��L�\����T!�fÙx�[2��æ��.M5��Y�&|��m�p/N'mR� _�*���'��%=��l�T��>�O1.��!�<q�V���vp y�7�X�r�c*L�
�V�DI�s?��ꕽH,N�e��x�;�][�fJ�;Q�Uʮ+�C�
�.,�U:���=����?p;tW��_��H�\1�~��m�.�B�ޤJQT]~�1�;x8}���K�����&U�ᩉ�U��å������s�5�Q��`ꑕE��U�y�p��H+���Y�~� ?+s����,��q�5���n��4��#6��'��w��syì��N�c���f[��.�"u֗(�o�2�_k�,��H�/o撸�B�ټ%�D$�A��]u��ԋ2P��C��a抁ٱv.
�Jt3W<���#��P��;���u�ye�/�`�<�NKGر?"��,�`%��v��+�U�� �=�"O ���(�#Pw���I�!�&U .��ɵcƍ�����E,�y�
�0�(�9�U�}s౤�a��\7sت�q������1\§�w��k���?�r�'�0�T'D�������px�/�n*�%A�&Y�s��ϔQ�������j�X�$�Ⱦ�Jt�'�57ۿ\v}�����.�&��ya��j�Ԁ�!���&PG'ӱMh�������#TGݓ�9�wLGBy�\ ���?��O8�����[zu����삔9-����]#����6u-��P��w oy������G�,��(������[14���8�@�lKj��tC�w��"ڣ�O,�U*yNUVv�v�y���Ň�����@��1~ң/�����+�85Z���ry^)�5�A�P֋+� Qߟ�q5V6�_,!޶�WC�F������La�ZRy�
���(�X���t�}k(��D-X�ӿ�MS�J�_#���4U��2�Ev5\w�M�r�^����롌[BXwa_64sᦙꉴB�#|�R���w������hAϖ5��*ß�3�<�������K�~�ƹ��L8��6�ay�m�[K�#̆;�gU�d�hZKH-�nM9���4��X�� Ji�������ʲ�OJ\c������*̩�i��x��L ��s?�P �Xw'?I�%�S[)Xn��,/�j�E
�4�k�DX�ѭ�M@�<�>�z��(ٳ�l�J�� D�z	�y�3�i���$�9D/*�HT���1x�)�rT�
�26-crRՕ�t����*�_�M/��^|����(��m�g��M�, �q�AX88/�K�N�,�\� kAL�X�z���g�~���!����:|fLI�'#DeA}�Q�SNd?Or�k�m1@��@d�PĄ��\ˋ���zv�s##맵4�^={n&��QO�Y���:�c� �e$[|�_��*��&m;K�=6AP�����g�ȝv�-��(\r ��X���K��rf�]�B���"���+�3�0�d4B���sUQ���ljH��B|ڔ;čȿ#��`����	<~�^DZP�&�E�5�2�Ĥ3fo�'<�� �E{����x�׃�Z a�a����B	�6D�5���V��.!:���ݾ2A��s��ݼ�<YNɐG��$D�
5��y;9��R�|�uwWxt������I���1��p�]�����\2t��]���cޯ-�Y�M�`�G�
6~J���ǜ�Lc�ܗ:���q��#��$�%�UlOt�����d�j'<�G&�Ѹ��Gֵ��R����$Ը^1�VL��š�7<#��j�lY��3pq�UѮI(��o�}�<
��� ��k}�-c��t�W�BZf�ܘ��{�>�;TfM��C��|��-鏧��긐�-s,�_�.�x�[|"_��R���T���D��*Ќ����8�C��
�"�qR�W"=��`�"��q��h�� f�2:J�e�P�XK��P�;C���tk		h(��< ��;��+Ic��� 3ʌ}�8��m��F\�
Ѝ���g�p�*w������M�?
W�<�$ݤi�b8g�{�G��qEs!���C��q��b�"xe;NA		��0�hEXI��,���׋B�i32�1On?c����e�-�E�0
�����<Љ����6|Jw�ȷ�c��ʓ�3��ӳ��m��[<�7RE��� �J�%�R��L�M�,�E���i���UbpmS{��hk[w��[���ru�V@�S�ڄ�$3L{���u����QV��������fY�sifԧ,0_�9IM��d�x��^�1\�w7��j"�z`S��Ӡ��Tb�%V?;��f�ፆ���G���)D��7�+5ţv�[O�%�+>����	�Ur���ގ�eb~\�j���a� b��%�E�t�j�<��߆;�+�!I�Ы�ݰ@Տ��R�N�		پ���ޠ�0��n������V!��]�/�I�:~P��yb��Gih��/�h	�^vXqA��ofr�V�W"�Xϴ$�VX��Z��#��7�T�~FN�Ƿ����?��Ţ��ŋ��吾�T�αZ��۾F>K�R&�T �/$W��{����~x���֎�D�=�0���Bܬ�e1~�8�73��Œ��mn�=[܎ѩ�=O�WΈ�b�b�|��yAeM���0�|��� 
Z@3ԬX\x��υ2�׃n$�ɶ˚�e��]��!;���*7	�{j����}p��K��V�Ek��d��SKxq�ԥ��5SS�2ˈ}Ջղ�H���Z��D�UhdvT/rSߑ}=�޻�(�dq��.ܟ�R<�-���34{�� !m���X gk.�G�LG��%!s�$dZu���j��b�+d�18u'R`"�n�5�Bw��q7&�z�f�����lw��R<g_dl5}-�+R{�l���;z�b9�V��I]�q).�(&�r&����A{;Rb"�dz[�����Pf̶���T�րi�滼���$\[���oI��s1u���X9[�|�'�9mO����!�$BWj�:��x4�á����H�٭�����u"{��:�ҹ(~�HϞ�u=��8��7_�T��<�}�2�S��tT�\�6��Ym�~")?�zj�=mj�ɪbS��ii�$���;������fEo̎r�
x��K8����׍(�n�nj���D������!��90N�&۔�a��7�an��l��(���C'�CY9hϮ���;�*N�*dm��~��Q?&&>xI{���9����RÚj���C��
,`�̀��Cg�_��dt�{̧i�1�&�ӷ�xc�6�
����j!�vC��!
oi;�gDw:r��k����GQ�����J�]s�*�F��mF�Ŵv�7����i����L6�����Ά�Y��B��hY�5�{�l�N�f����<Zb/�c��8��+fp^݄�k�$�'*oA��(�3�Gۻ�\���ff���&ĺ��q�߁��/�]�
/���~��8C�\��^߉��z�x�&�a�&�V6�_S��+�h�,���5�Vڤȷ��l���F�vc��jM�����*��}Ӫ~I��;�X�Mv
�����p��#^r:���iW5ǒ�m�)�C��긫UB��/��7�JӒt�ʻώT�h[��Jo>9<�MV�>Yvx�L�b�戏Y������>:D��`�'�b;3	��,#�>�5[��N�{r~��
���|3u�㑬
�p��\��*��$��7�_���<Bp$�G�(���9��$��3�q&�RéU�DX^��)÷S�T����dY���T���6�Y=�y�'Ӟq[���A0w�w	C4ePRy�����&�Y�=%�1D����7Nn0ݸĜ���.���ԍ�]��Ξ�I~��ݚ�R�Wu�`�N�J���	1�)�3Ő����y�~�PM>���	R�B�Q���Y�=�m/��V�HNoХ]hy�I��!��J�'�O�0;�z!��ζ�Xf���7�^�V>�"��D���-"F�>����i�>R4Ι���f��k�q�{y�ڍ�[�Pr�@�w�n𯞑S���-�s�F�mx�T�s;��"@`̚N�p���畯��cMu�քu�"{�A{��6��^!词�J��O����Vj��%�[�r���w*��?��6���ޒ}�f,�p�+�)￯R�1���&}}����o�k�Uyc,*t�n���-"�]�?qV�i�Q�p�Eq�؅��9ױ�| �e���J��G�#�hVg!���*kF�bZɒ�nχ!�A�{��y���k�%2�P�Q�I�Zey���V۟Y���wR �^���G�p�7��TK�i�o�b�R�xTz�M��|�U���d�rP�B�z9����Կ�3�d/�܅D]�@�Cɢ7=�a��HC�>��.���C�=~��<IE��š��i�B,L/��bÔ�}?��veQ8˅� ZO8_~�/#�ay����+�K��!L���@ƽc��Ee�bJ�\?p��� =mV�O�i��"��"+@}�]�I�]��0��_��4;>ӏd��X����u�"��0����P(��G77�m��_Y��L�Xf5&��Ԗ1����L�P��j�?p��`�[���pψ������-�S����D�yaI��9�R� ΡPb���@�q(��|�o�$l@���ׁ0��ޘV�Ol$j-��P�6^�5m*:y򶂨�O�:2�4��`g�뾎!����h�5^����yG.�a��>���^	,$��I��c��1���@\����yAք��WC$�}3zb�?�-�D}��ė�E� ����LB̤�G~E�ѭV�@43W�FzR��5(��w쐏�v����.�� 0�%��{��q���ú(r#8џQQ����'H���(b��~��2����u�e#��x��7�:���@y�`���hw�N�P�u�i��#WE���������Q�f�s5��8�&��h�>���q�;)��8�sII榞� �,�{�(������cڼtS�#T\�Ŕ>����!��
+.#�qV{ԂK���=� �H��YW��:�x��/��I���LCu^�"%��c ��)ئ 2a��7�k،1�NŧL:�^�X����~�s��k$�������aMa�5��r�Mu0�5g�=�2��~�;�����[�T��K�OacA���t�<����K�Jo�tB�~�9�S��q�K��2�VF<&N�ZA����vU������Փ�4L�A�o�:��T���7�j�67�qz6}��ך֢���X=�k�E������Q�X�(�G#�76?�@��A��ҘY��au��1�2G���Ot��j���u��g~BpJ;k�	�3�@V	�1�Xqq�#��_P�2����5L$�F�?~4�q�$vmtft��5#'`>^"w.���L��I,Gi�9�I�n䀡ʵN�BϨe����ƁaD��O�u<
��%��E��������.�^��~��.ɲ��P�5g9��]I��I������T�@<�4�*o�dW�=|:�z�mψWRUn���5�/S���K�y��{���C�����D�"�zgXd�e�
��һ�C�n�)�Q'���z�;∙�W\��`}��G��O��-ʲ�C��������~�a6��g٭L0Q�"�D�TW�tc�_��j�6��(�q�D`���[J��Z7�۪���ҳR��q��j�je�h{��#L�hT~����gV9��g-���u�O�,�^��b8�b��=-�����zx�,̢��nS�Ŕ�kR?\���� �J�Kf�Z��ǰ�w߳�7��[R޺��CFb�Bu�_X�$&�j��d��w���jU7�tTY�35�@�a�0%;�_E )���[+��s\>V�*b�t�2�x?�ymyKٯ�s	g!�T�t�F��gCW�e?�Y2s��F��r�/]K�M�������_��"ع���M�Q�I����ά�B.�:�	�t�n�"YH�u&.Q�>�,�����?*W�cRk*����Y���T��:�j�G�j��A+�`���$�����V�]H��;"�����b���g��S:{]��<9ԃ
�D���$LP_�}�BT�=̤V�n�S��/�|��ba��~��v0#��V�`�x3�� 1nI�Ɯ�VQwU�����Fqv�<��ކQj�m�M|l����ߋQ.B��s�P��x�������D����{ C�5m��u������C�O�K	^��l�^�^ ��u5�\"��2Ga��m�JgA�!�0���71�f,˭�p���'�D\ǁ!�ѹ�V4P^|�k̷t޽BΦ����y��|�gw�:���:��!�f��ݨ�\�Y�Bl3�����"��Q�Cm)[d�	��~f��*(�\^�*�Ƥ�/-f#t���:]$��/r�Z.>�rv��EӃ�4dAjO�i���^(vN�>��^����G�hW<?OY������ҀD.�M} 
��9��8Ϝ�/�,��}�f�)�u�D�2�QZm�����1�yi؅�X���痥OyŒ�б���t��2&T�١	[�'	�����^��h����ޱ�smx[3�Dcn�����Y��_�Ƈa�
����r!�e��l}:�j���b֏�%o���nW��m�vX�X��
,qg"G�Ǒv�L�7�{���� ����Y� ��c����}P�B�8ݕ&�8�O~���^�@�϶pd������K�O�M������5���d��l�u�� �-x�У_���^K��]3"R<Q~�ןܗGV$�[ۮ p1����ƊSO4LS��d[m�>�Ps1���ŷ��A���/))�$-�pq�����8����\�ݒ���k����B{s(��y�4:������[70:��L�PU��)������X��g]Sb�V��q�Lc�d udʹes	��X��h����ט��x��&8{�*չ�6�vRZ�x�z4��hn&
��C�f'��i1�%2��)�d^��aVs>�<��`���<��ȯ�(��Nts�)V�3}���bu�{}���Z}C�2P$c�%ς��+�v��"qIڲׇX,��e6`gB"�ߴTIPJ���e�ͥ�$2G`?�2g��흀�Agc�J��Զ�xF��"v�@#�d���Z�+ߩ|N��l���Z�᱗����d�DX�և�Wy�:c�g���2c6jͅ\�Nd��v
��oD�j7���A;��4p�.;�]�t^uơ�_���fX��P\9�P�膀5\���Kd2���*Y�N.���]��"��d'���PP��-��f�@g!NJ�cK�b4$��5����������+ك%�>'9�[v�m�=h��c�=��^�����Vǔt�L�Cb.��[+w�C��$��(%7 �e(��W�V�I���V-��MM>��;���e�=N&��WuKĘ�L�j�,��x�0��C}kȷ�k���VgR�����$p��	��*�4�i�4���xș��CV�M�����wb/�X G������S5݈�� N���o��?���2Vil�Ĵ@���L4�o�����B(�Gsc9�?2t:�c�Eԗ�%��J����tV��>�{����e�%Ud��G�k�?ǸԬ%��?0D_�n
a��t��3���,��	p랦�1ղXPl��-��忾�7�h���Y]pC�H��s��_u�8v#a��g�Z8jV�Bè�����b4)�(��H1*�ϕ�[&�!�j�ߏo�PX�!�
�Fqcd��/}��s��9�֭�֯6	7%
�LR�K8I���x�p���>`l3c5�d�J�N��nb(�Ge3l3r����͉	]�
���z ���
� �W��� �|�%ƌq{<�8\E##�u|0Z`K��ݾZ�B3p%��ɞ/��0�a��X6�Y��T/^�B��7�UC�B�xU;��K���6��Z�!ˮ %<��p+"8�$������A�ॣ��ǵ�Y)7Bz�A9�iM�۩<C����璢���G~�|W�冀�jR
-V��irWԐ#6���~w�O����ꄦ�~�&w'H�B{ET{k<����CǺsa�Q���-.�f�&.z�a��C4�Ó?�� "���_[^P�㵩�uW�RY��m]H���CBR9�]�)k��s���I�h�x�H`�eY"�I͹B�.J G���/kо�N���\��_	ܝ�����6DB��ҁ񩇭���
��4�b!-3'U�O��A��hv٤l��}�t���-�Z:�W� +x�� �	��D��A�M�����'��)UȲǠ�HDDw�^ �d�h�q?��k L�AjV�b8��a��zB ��9즙N�Ľ���i�8�����#!�o��7�͑ꊺ,�<��-ۤ!��*�ޝ7��T�g'���I��̵�Ҩ���Z���Y�-Ѭ������]q'�D'�gxe��5���~5|�H�]߷~Y{jxz�P�.a�)��T���D��o���!��ي]t}�j��W�	'T����#���k�SҊȝ���3&3�o��"v���<Ÿ��ޓM��a
����M7V�����{�؆�bI$ɜHR�e��N�~2x.�bb8�6�;n0�%��`���{��'&��K�Q��U3٩�E%�(b~���MW�s�@>�{�z���*V�r�:R&�U�I@��4������$�ӗr�} ӣ�P���ǹ��8�>ֈ���:�5m�%��ͺ�K�d��lR�\���0��1���%���}v�g��VV����A��C �
p��z���:=�T�`��$0�ȡw�An�g�,].��>ږ�lڷ �>i��l�| q�N����P���vJȉ��Xʠ��Q��I*�V�:Ѣ�m��e��n)�6Zp �ή�CAJ8��f�gFY�x�ev�
�D�%��	yv��H�l��x�f��[����7�X�l'o,T�pm���wʨ�+���u}��v�q%��؟2Q���x6�~�Bk�i��N��>�u��˄`�tr������tdJ�_x���DZ��,�uڸ���ԮK�ٻ�!,<'υ��&�D~�KFَ�	�*o�4k�eWvX/x�K�̙�n?c�y_`7Y�Bi��,H+�|p��eCi���`�t��PQ�+9|�&(��E�tiָ�l����BSnl��Q�`�M�}�({��8�cF5���^ﮈt.'ǟ�jd�7���F�H�࿻כr�(?��^C�g�h�<08eKŅcru�i$��w�]y
��p��E�6��{�oj��.�Y�"�{�y$�&��Ů��	bf]�$�6\Zg%*�>O�Dp���	5A��`A�篩�z��ѩO����@=���� ��ma��
��tA�-����	�7�y�g^�zǅqr���������G����Ä�I�i��%��b}Ĵ���gk�4���nn7n�4�zD�)���)�s���!�=��V과p?���q���K���ڧ��Y�)�Ы�Ŷ�Џ�E�#9�;+YQ|�~����5����*O_23�	ǅ͝���%�(���V�~Ն|�P2c�@o�����J5��O�s!�@4ࣸ�^�-��
[���w� �Z�o���W&K��#u��H�~D������<���H�]2�?�_g�L�ϒ6�%��	�,t)4&A�,�Fg$�^ՑܗZ�J�@�;p��2(6t�W?���v]<$r� DZV��T�⒳���3 [cI&F�̚l��z�!?XX�(���8P��/뗩��+�i� �&���+��=M�C������L��բ���o�{3k'?�e+8��B=��31��yrv�\����$ڄ�e���*�Š� R#<��6wJ�P/�q �/2z}�f'�B�x}t�c�P��܃�S��T1VZ��sw��^��Ҁ�%��K1�8^�9Ź��j	!�Q%�?Ѵ���v�T��(y��"+	�H���j6=%��1�Wy����kh�#VKS�T�0�RL�@�����XN��������"f�Bȭ9{��r0s����*�/hR����TL�( uq]�'�9X{�>��V8m�s�q@��Ծ�$��/rzg'熘a�w�]��_k��{d����k�rvzT�]KG��>�Mhr��G��v�ǹ��`�a�ȭ��5�;��m�X��͌^�/�T(/O!R�}~!XIb�"{}��%�K��H��������$�#��mQ�����w�R���֗�-X�������;Q��g��K�� �R߻%3��e���#��KSCP�Ҵ? ��|�ޣ�����hM̏���S�:�Ё��-y}����Q��^=�qN:�281�[��f�nP��j	,<%x��;�����5AvB�`ƣ{��8�r���͊zmPъ�@����E4�O��	�u(A�-�
Ƭ�Q[��~� �)���M�ٖJ�9�LpdN'��i�Ӆ-����]$�JkRu��WU[{�2D�B���1�h��TkQ�|v�^�$��t�b;�*+b�\�_�&}�iJ���]��Thиվd¥����_!��yF�9Lw�="6�B���Zf���E"����NK6,�����j�U���)��?�����6tL_��2�8��$�4(�z/�y�a�b�~��6l�� �x9ˬ�Bk��6ˍ��0I������hl����	�HC�릦����@�k�����(�G0�d�W �&�d�c��(�*��iȆ��=�;C%N�V��:���Kg�넵�R^z3�~���/�MoR���\Y"��c@"{���P�7�K�g����&#�$���c)�X��׳��C]��
>��6���w�,j���v�e�h�!T�Q[�M��v����җ-c�]}$����#�cU��f0����Fy�:�_OުaQ;F��v���4#|��d%�V%ڥx��c
�S��iQ�;�i�"�I�[��#_0���:���P�tC����a�sD��դT��,tj3�f��R��42�c�CܜVr�=��lZ�"���uܽ��`*{�g�M95a+{���&n���G���  ��)�i��a1A�
!}�+�%�Ar��7�)�鏞��B�&WWy����Du���|�1����%Ί�'�c^���\�j9��$��L����.�'��Ri��gK���|6ޑ�'j�B���sl���n�v�5��U�sV�V�����=��aԧ�����
�1[XtRf4�hC�߽��@K:�~Ω�G&��Q��if�{�qC���"�5QQo+j|N��RZ܆|�:yk�ց���ׁ."�q�-��:�M0{υ�3���崆�~0[S`�4x�骲�F�Hw�M�~�Ь��ꮺ��N��db�~�.����X���(�@��/r$�7?�T��II��WB�q!�A9ʁ_��&��0�i���]�B_��,px�>ϔ�C<�`��3]bH(��hMڨ"�,X[�������\D��0��0�����;�ضϝ���zy`s/��KC��EM|�5�`���rq+�l�4�=\�x*��rր���*z��㷂��1'v�|�7�\���B a���Y���3>D�q��N.�fu"%$0�n�%�d72�S�g�Έ�L#�O�UDg�c��#c�m�x�)��n䭗����-���})�,��V�A��ޮ�R8r�=�5���8�%���j+�I�1�N� !�Öc�U���F�z Q������U�Mg�*�|sPh�Os���S�$���)��uN7��m�������ǢN����:���d�~Y�����	��}�w���՘�u:\��XA�Z�e���ӭν�5�K�h�&�ۯ���gd�P�V�E��x�<]W詥��6R�N7�6!�0�&��C��r���������%�S38��i�@��\gk��J�wD�Z��������� ���O�-g�|�D�I�V� �u'�c�~��C����6�>&~��oZVs�X6D["F�(�X����K�%	�sC&7�m�ҘxcY#:m;̂��JF��ԙ6Pt_u@�Uښ�B(ޝG� �b�?����+�a��a8H�[����nc���tԍ� ����%q9ؓ�U��%��h�O'��lJT���.���wyC�U�Ʀ��6���ሱU��d���J� �*�P�����H���NU4xu4q�Y���>����� 5��$�g��Y�8 {4&�]`�?�v�
�2Z���oQE�GH� H3Q�a�V�qQ[��+3k*��O�ˎ�8z��#�!U�ۗ�'9��q�����y]d�ӼS�Rz�I�����y���]�ԜTˑ�fZ_�$���}_���)�u��jZZ���e./֞w���X�ě���{+YX�'q?[�-M�M�o�~����Ԉ���(;?>E*	�gڄ�Ի�Q��v�v�����Pʀ�����5>�=ocs�������ư�O�2�����n�%�Ꜧq/�I���g0=}�F�m��*�B�b�6�o/�6�
���m���30�-
��!0���ƣ�鬒6��7� �⬜�c�17�W��*Y(�E��r���j��;�dZY�6�{�엘iKL�K�X<��ꮢ�B.�^$޳��^S,=X�^��f1���Mf]o��:����)r�&/�?2����),��;MC��������I��YP�~�N�w�ۂb�栁B�\�(�(z���j�?��T~�;�s`"��
`~����:c|ڄ�x�R:���?r�z�у~]o�@sä���3建tH\o�F�q�D�Oh�c�-_I�`�"�p�|� 3(2��Znjvh�뤬�Y�-�U��/t���6�/AG�%Ց������qe���i���;��OI�0[����QUe�y[��,}�-�S�_�R�yT�4�.�+��ٷǯ��"8�Z	)����+��o)�T��ʤo����f���� u�� �zj��#�F�72YT� ��G$N���߉
I���i`��	3vJ�Vz4��徽[�K@�N�r�/{������8��-��l��/5�G�k&�	�Bc)J�5�4�8/�龑�p �I��в�-�M#x�I�:�|V�{]�;�8a���Bj��ό5�!;�*iV'�6D�����^�R���6j�7:����c����xF=e����BGE��gl^��̳�_`|{\v�WɄg@�/�����C�䥼"�L����V�
>��x�$�Ļ���.�M<0Q�m)a9jJ��)&�ZN�NL+�uGJ �i(���[1-(��ό�L��i-�n`��
.���ψ���p��p��Z��U�`Rd.���g��%�⣑���2��9CJ�zUv[&�{z�}�ѭ�����Y�h^ܧ�eWP^�Vkj����3�9jz�������{�.y�֢�pf�_����@(06?�6���p�N}��C��f\h}��?�v��ʮ��k��E֯ ���ZFa�`1'�m��U�m�s��=G򋈖�Q��\�R���_VH������xпG��/��JBY`(���8�G=���}\�q���`���cFR�ɓ�����Zv���d�)��D��ܗ1��4.F�� c5a\JD��tl��;� ǜ���7����`(�X7�ʳ�~�Х��V��� n�����vo��~FQ,����(����T&0oŉ�v�	��9U��N����|]�n	g��s���y;+�a�����Db��Q�S��|�R�����w���(�Pv?F]MW�G~�� � R�2@���e_+ ߦ���|�3mZ�<���� %},���d:���_5�fط�RU�\Hw��/���Y��>e� �b�#�J�-�(%�� ��!a���<�#"W�؟�oo��N6�4�\�5YK����Ӊ���uH�4ѵbԞ�򌵹"]d*�4���c�t���ɞ��2��y�^b\��zzׄ��_ͲC=����D���U[�#�1Hz���dx�~�~�,���N��6U����m���a�2�땒irP��5W^��8ȊM�:v���Lo�F�4~��Q�ڜ����|��,v��`[-�?3SX
�TN�*%�>vO=��N���g��Q�����N�v(W��w��L���7.4k�����b$���1��7��������-j��p]�Xf�E����*=�E8?�_]:J t���j�+�Ȓ��L���M���aJ��t��٣a�_ m	��ʱs�G��^P��$~ub]	�s��.�^]c�Z�q�wB��>�)^��F�����ʌ&X����k�������0'U��|.m+�]�X�!�$A�w����^�L67S�ݰ�8(s�Om����1s�2���<�>�z��N�eKY��?�9��bK�i���`�H���B��E���H�\���٨�o��=��:�p!:h��[�Њ3�q�i&/;�ߊ��E��ǔd\�ޣ}����:���>i����S���B���� buĪ�}﹗��9�,��I��BY+!��)O=*�o�/y��=��D��J'M*�f��v4Y7�������L����A�����.a�?��.� |��/D/k��XV��Կ{�qI�:-�Uò�ͽϐ����1��2�x��T=�7@q�%X'����Gn$�B�O9Yj?�y�l6��Wgbn�$gI��9D�"7�&dt*KB��v6s�(� ��1�jm�ѫ���BV2\���1[�����{�pU\��0���A=%+#e;g�Y�-��v~*T������J{�1+��:����7G3��]N�*
:Ke��(̖Fz�ٝf�-���װ��y��䝚�p�0�J��ȡ��S�RE��ɉ�X� �uV�F"� /���Ȇiòca�q��/���K`�;˶)y�m�J?	T�G�m�b��,���Rա���w�}ix��+"��Fl��]�}�\x��zW�y�F����u�xܺ��O*	.�4\Df��zp3+�r�a=}��0�a���ׇ���?� �p�<n)nF	Ԏ�P��3����;g0b�O���(XoOէQ��=JP�;	vd�X�6���N�d<�Z�fn	Y��aL��5h^��TWX�`�o����J�R}��v?^-=/ISBծi�KQ!8�ˊM����KuhL�$��b�4�暆��:q�V�"p�j3�T�
���MfZ�$o�x���A���'3�[�{|���?�]J옵�d/p��ٯ��/��|o�y5k7��/����`J�
O������߼��K�*s�?Ƣ��Y��\Vز͹�F��n�g>�6zs��X�Σga}2��L �G^2X �Cn7�s#�h`.n�n�%Hʵ_e�Q4���JD�$i,��X�������P�k%L����j�����Wn�BR�G����:�;�M�Wl��(�kd*/�O��g�
��n���bc���:����Lw`�|۝����3d^��8�,�8�L%ס�8���쇔�,unE�����i����NU�Mr��*�,�>E'�}�򝰳ޝ6+QhDWl�љ櫛/?���'[���9K=пU��1�1�ˁSl�C����k�$V�-#؞��x��z����:ؽ�p��D�7�����֣��~�L�ڍ��yr(�!�*��?��-7sw>&óKu�/�y�&�q���s	B���r��;I{�-��T���k-a�'a�M5�"��vcL̔�8�d4��7oX;��\3VZ��rz��b�9nAء:SI! ��^^d�e�)�{�Z���ʧƉ�Eގ��jD�Hqg��-},����*sw[�����%�B�������@��}m]I5�8�{����oX���Ù:��5F��^���8y���q�I�W�ۮr�hX�����Y�r�@�S���(�I^�q��s�h^�����7���swo�7q��&������&�@��|��k6��4���_�O�����<�;y�SG�H�_Y�vK)����"ץ�$h��&�Y��W
:{|��������� ~t�V��]�Ꚋ3�$'}�@�'{G�(��"�!�hQ������+17}3���;`�P�YG�B����|��a0*s�aƯ.o���k{�G����m��0k9��9���+����:A_�p��ȼ���Z!��r�ŭ&�n�(�7��f���f�c�N<U��N!s�C:��XI1E3�ddxE���xV�Y�@�/����t�V��ե>�:s���Xj���X� Ѵ�z�~.I*�x�:#
�� �;�ǯ�[䛣�.T��ر�ƒ�$;�<���|Jz����a�(L�A��!Q(`�Y-����갤��-���F�n䰥)�4���\��Kh����מ�Hѿ	���b�����CK���Ǎ�ͯ�|*W�S�f�&��"�8<�?e�����Wꨃ��I�g[6��Ŕ�/ a��Wέx�nw�u�F-��.�É�y���f�tKN�� ���d
�U�ipă^
��!��{�.C�'��J5`.���5�Iy��Ķ�_r��	B�w���6�� ���Jű{��z���ƒ���F����L���I ��D��|��+	(mgS~�O�*}¤<i�v��d�:@��l>h�G��lZv�2���Q����i9F���OJ�B;(y�w����4�Ju�9������N9���S�_�e�o�uu
/�uń��
�T�#���-��
rv]8,k5��Ƭ� 4��],ʉ����!�m��	�U3�o%a!~#��=��sa���HYC�ܕ�S���x$�&�FЊ㜙�s;��EP�R��mҩ�n�
 P���e)����qr<�gGӻ����9r"/��:�W�q�;�J�����g���P�*t�(��ة�1�LƘ=�K顏����V��2����+������(�l��,G����t���Ce���S�ۜ��&?2���7�)TUЍ�����`�RQ��,���ɪ�y2l��K�+n������:F��P?Hh��"�8
���@����cy�b{G݉�d��wH�M;���pd��^�&���P���s��n����q۩��L�Y�J�XyU5��WxG�"�o�K�֔Z5���x۾˽����~���&�~��pgK�;���쇒+[��	l(Ħ�Y\[7G�^�\v�V͠sH�M��%ߒt��Mnl\���ׅ>�"�dݘD�t@=��Gُ�)��#؃�ЪZ��TacwktS�sVw��ov�S��5��t4�d����<�|�������+{Mمd�	��yΤvI�TI	�e/�H���rբ]5��^(Q�$��4wz4SQ�i�&�����!ʤ��c䂗��N�k�$���I��ұ� q۞q��t('�݉�=����Pk��\^>�gRyڳ{��x1�6rp% �b$�|"7�x��e��ê������m,�D��Ż8Ӎ�`6X�q����BRN�v�DGV�Q^��ba&|��K�,Bj�zc�X�����neB�Ů/ն�bw�a��W,����p�l�(^K2��iC�A��l��|�*f������dd��<�F����C�l�z��ϧ�A�����V1LX$l H�j���ft���-h��{�䩗k�ڗ1�$;Y*��S����m������ՇC���n���x� ���D�Y�x�M�	� ;4S�_�o̓�e w������o��.��tc"��1��2^�+�S���F���=0'�J﷍3ɝ�"�i[ı6� 9�8�,�ܟ��%���O��SۃK:qh�� �*;0��� �YA�x�����/	e��_���%!�=�5�cn���	=3��߱Ym���^��tƣH={����N)�qZ �0?=�*л`PX�59g!�V;��q�/-���  ��o=�����~_aq"���I�`�JJ�j�+��K>5@V{o�1�ɑ]3�{�]��@m����Sr�"J��Hm��Y�/�
��r�И�E�ť��܁eC�,p0'���uFijN�z{Ʃt��Rh��aryB�\52r�h�h;���/�'�Xa����1���؂��L�k���nTH��1� ܲE
oA]Z�h�f��Ao��çTt��V���i��|���{Ef�%�w�`NT@̹qN:�)�������R)���sV�OZ�3 �*��n��W.����z�z�-��B���x�!v���.�O��A��'�;�!ڴ�"P�
��؆�v�e�P\!�`�LvS#N�vU����&fi��_�^G��S@��&����Q��'dP�	�?�>��H�w1��ncKq�t���ר�|q�gm�p�>Z�w�";i'��(sE�zvF9�Db�Ч��b
(H"�M�U��J�T0a�Ş8��_s�N"��Lz�ԝ2~�iۢ�������]���j��eag�@-W������h��"������J�$I�A�Y�o��X�W�h�f��a��k�j�7�	�wL�ܐ��.T3������ ��7W(m�k�
�K�=�U	�?��u/�����pW�jB<���k}^��J�͍kmQ[ք	�b�d	�h|�TD B%d��3B������k& �L@��
�'��٤�vg�w�[�.-g�b�/4��g�C?�5�͒��>��Y�[b�:^�F�D��HF�R�t��zS)�O�Fܐ���Z�ѫ�E�B�y�����"9�|>��F���ݗS[l@S�	1Ÿh@�V��f7@yP���<�T�@���-�L�̮q獫�F�Cd���^�IC��~��E26�*�%���������P�ED4��m9� ~sЌ[M�5l��vQ�M�+)ט��ۥ<�TV�Z���M] �}�am�<�e!�
��O�T�l�Y�7���x%Z�zq����e4�r�[�v'�Rd�^ �"��Eb=��v�(�6�U�H-�9`bhs#���E�ݙZ�K�+�e��Ե}/����+y!.��Ћ͵��w]��ϰS/=�L�/1��D��8u�|CO�G���0�MB�VM?#O��N�W�m�}W�⯧� �ؒLK� ��-Y�	�V#�K���$Mrh3�K���Մ:���A�n�t|h�ܼ)v�r���L���U]����A������*�wm .]�ٓ����E�`-r_��x3�;Ĳ�Œ�p4 ���L�n@(��GH���B����@����2��l���x0���㲗#�N��	L����%Z���=)莪��8�A@n:��w�E��W�K������3N������)�F/z�=<���%��)�d�l��{v/0��?t���@�����)"��g����t�6��m�ze���r <ZG��$�-u�k�Z���߽v ˘o٦y��A��I�[C��XX�>��4U��$�xGXP7�D�\�sy^`I��4���ڦ�K��^M���1o������>Chx�{Ӻ0d�%�e^���=26�C&�8��h[0De���H���$T3�ސ~u�����F�sW���v)��^�����I������B��!�Q�-e�1�R�Z+���o�~��Zb���(��<X/'�Ft��^���yN�d^��e}�m�+��{ݺWj��T8{�4o��Kӥ$l���z��G�a�jZC�ךf��j(����5�oB���줹��4�UlBr/�I���M�a�H��-S[�[�Rs2�kd��#Zq�;s@�F$U�9K�<u
�8/�.�>'d��+��ŕ4�N%6V%�$����H����n�����=u���!�T4�`R@I���q�)�0Y�C��"��#�[x]C��k�[dj��I�c����Q<s��[�;G����0���K��~G�˾G�2�=Ч B{Ȗ��M�/�Xc�-�5����e�k��+��;[`F(�����	�:��N��9)��\p�"&<f3*�hų�6�C�T�[�V6ԍ����SW8 XgRD*J���v�W0� #�$�|�xn��� �0����pF��$��ǩ@��S:<^m6zq�N�U�[��·d����g�q?�W��E����-	��I�N}A��F�v6 .+2���ز%WQ}D6p��-u�G�,u|
��]�-2������^Rt�'���k�!��;�b�Ih��#�m�^ׯ,1oC�N��~�^Hh���՘��ӻ�N\�ʅ��}z.ʾ��c����#��$�2��By6͏�U�)��o 5�`�
0�j�����f�4���Lt��L���{��Vx8@a�~��g��E9���j�M�#0�3ʹIv�0�B��NdBc[�8�d% ���.����������D.��;�kyY��2��w�g��d���&#���n����7oܼ �!���u򄑨�ƣ;�1f;j��؎�.�xN���|����s�iX���I8�������M�i�i�Dg.z�]|�<�k���ôrsJy��� ��-��A�M=|����m���l������ݬ�V��p���:�X�-sX�LND޲�-c㺝S��_��R�5�2������tF-�J�6wj��M&h��،Ô���	[������lLhq[�eE�n՚��,�ز���+;U_|��Rb��uX�V����x|��
���A�mK�^$�^�8��ǻqkf$}"��'ۃy4�	S~��}�E�.����M9��^o��p���=���\�Q
�G"���0���k�IU�0K�4��Ѣ����w�߇�P�D�r,M�!{�}�Z�\�ܽP��b}�f���$��꽡/�����I垢�B<�@)㲋��W:X\��]��f�ul��S� ��]�3k���D'?��b#����Rd:�����+p0�ѩXA9=XJ��B/��!TH1'�|j�B�x(������lI1ϲ�� ��ߞG��oQ+ȋ%%�u�y$��ޥVS&�Ɩ���`��kz;+l�Hڅ/�n��XB��1��'��ͱd��?����O�?F8�)ڊ�[]�M�?��n ����ZR
+�K&2�#;K� ˀ|�,�h�\Ôw_��6����N���4���ʗˁ��e�૟�T"���p��c���e�<Fё�%w0��e���g���p6��*;��
)����If�LnL��
G��_[]�X;�V�訤��E��-z�r^`�6�I��P��N"y����s��9G g�۷�c�/="q�������x���_��{���0�-�o��)7�9��o@�c��s����5�T����-c�F�U�1��ǝ�z��o�S*�-!P]3G��uhgD�I�?���z�/-�F�h�Y����/[��ވL>3����u�T�v,kI&�j���-tTa�Ѻ�l�?�\�	v�&�!�����iZ��4�ZV1��$��2������v0g����[����W������	�Bifm~��ھ���q�;l�d
ꣅ�6R��o��"�Ō���F���<���.<H��Wvo��	/�r��|ͷ�������n%/ņg�A��|R�l�M����a3�cǄ�y���4	� �H�Aՙ���j-��"��:��"��Ӂ��V`�-������r�����JE�S>�iv��ʟ��(�N�h0�Jt�s7Zu
h�� ��f�v����1����v2O�;>5B:E�)��ÈD�� TYU��Ē��7fz�rZ6�/�>{VHib������!�2��<U.���aZBqBoDF$���/�L\�?��wOW� c��d������R2w�WEɅ�V���8�k�u���꒗��w[u~,S��9h��%��L�4��+�<͔Rl<�	�gS��G4R����񍰒�U�w,����O3��V�x�SD����1X$��X���\|�v$b��ң��\�9��l��vr`!����ؚ�׾T�5a�����[�ǁ�*�D����_xJ�\��eF�,z���;c#��76e����A�*@�*��"��1��k�FU��c�a�㸍��8ה����x�+ś�ggPb.�G�C��¦^�F�[�2�����Q���h��O�*d�ɾ�숳?pc��BpH�}znm�2;v�^e1oR���GM�{�SGm��Y8
����UB\�FzB�5�6��VƵ���S��h��ճعo�E�v�0Zy&D�S��jc�����0>�6k�DG�
��dJ�w0,��������\@�9�g+�"�n�РC*So���xw(� ��J˓�F`�b��NZ�d��ƍ[b�dX�R�\�W�Is��r!�n�󳫜����?
]
mH�iݨ�Y�R ��	G���p;���Z<cXO�dC�-�j�~̯�n�?ɵ��]G��ڇKH������Ԓi���
.��7���(�3L�� S�т�ao�u
78?A�a�X
,�'SK?���c:���0dA-�)(X����{�n����u� ��U������P��Q�AWS,��4
t��{_T�՗��	�D��<�\(���وU�"e��C���f��� ��K;~���U�Y�f%�֩��Y���U�ż��=�E,Q�}ގ�e�nE���y٥�%�&p9{��s-%��V�^��� *%�z�b�ٖة=`Vd�Yo�GZ��Qlv������ȼ��򄕂u ��G$X�( �p�I�Ą�޲�5<�4^
�C!��J[$��m��!~�����cW*�d�>�S���˟�8��&Pt�8�'��e��?3'T��i�1�N4O���bc�_`:�����������و�n^4���{X��"G����鸲�X�7Y�eH���zӝ}�Ɽ;Qd�V���Ǐ����=���K����kP��Fkyf�.�����M�C�ך��@��&�2�!.^1Z�J�o�F�v�]��Z	���QE���;�̬�	��NwY��xoW�V�U�H�$m?q�Z,��j>��/�Q;f�g�wEB��5uE#������h�j7�f�\V���K��� ��9E�<����ii"$�=G�ߒ� |)��P�2�[�T@e��9P�<,,�A��6v[�6W��4�������,��}z���\�b �6�R�5�`�I���1�8�H�!�\ce1]<rP�Lz��Yƞ��t��v�T��DN��Nkӯ~��;Cu<{�U��o�J��g�7_,���[� �v���ڝ�V*L#�����A�?}��L�F/fA�/�]�d��$�۬n�F ����tpֈ�P��[��1K�ֲ���uq�n�Ub&������Q� 4'l��� 	"�T�S���ҤM��E0�D,�|��� �p����^��i<do�,Q��@�ё����V�8�5��|����TBָ���\���[d��aV.��XF�u������ͅP��'����M���Hv=G�S
���dyQ}�jJ	d��Qa��_���V��Q����4�?US��6��u'�p�.Uf�-��H��<+��a|p�GA�0-�:�8�H�ND,iT�@]b7�.�k5nR?�!V!s�ք�)��t��x�O"e-S��g+���^�����V��Z1HʁZ7L�/������l�� :#���d��`N�kT�m:Z�[
 Dn2���<�uK+U�P�C	��qM:�8x��M!(�NM�KY9|#�NSX������=���γ�A�����A�|�����l^��jR�I�(X(���.�Mi^��a^z�mTD���O�`���&r��Ӎ�s���fIcJm�h�M�ݟ��b�Ov���҇�A��w��ֳ�C��i�z_���O��y����̘ڞY��k\L��vlX�Wu�m�7U�,�9�囏q��)����W����� �P��%"�� �o+��+�"�!��0�	$7���t{����w��/u����6��PB�ȫQ~����R�]ܰ�.Js`�����{���<���Pw���u�祑�B{���@^��P�[p`�v�˪���-��N询�����ն,џb)�'+~��c`��v1�S�H��G)Z0'۫�=%����?��q�U0���ۗ�lq�Ԟ�D���<Ō%�f��E��f��&�^9Y�T1 ĬSl� w�����+�-�^`^9g���**с�M���o���� ��I�i+��
ZgR>��B:&�O��0t`�&,%�R�$�E�6rJ�����o�)Ag�>f�/K�gV�8����������)y8.r&w�j���G|�d�/�%�ع>��M	���{d�!J���Gx-^Y(➰���(��_�hr�����k9��Q7�X�G�0=M:؂׹KͱfY�ui�[!�HdeBxҐ�-���^մ5�'��R���~���2)�&$�����I���䛘u�nJ@�G�R���Q�X>�FR�y*:0�����K����R�#51�	�հ�F�x��x�"�'�SN�YZ4>���I���z7���	�"G���b������3�5�
E���P���?G�T~�V-���)I�� �"��b��֔���_q�|֯���Y�LS}f��]y�a�Ẋ��\��R�cEUP{�VP���*�Ar���&�N.>,��T�A1�޵?�i����	TG�h�҅[m�1��S�����D�%�����Av�s]��[�_	��^���܄�Ԭ��A���Ӹ%,���fm�ɘ�gH9�c�~T��6)e�;��"3.C��P۪ q��Щ�y_N�^�2Ni٭�O� ���U�{�S���24��O"���[��k�7��5@�dF�b�֙S�'̴n�I�y��@w�A����7"[��f����T�.��H�#�?a�2 �'xmp
���k�T&_E��A`�f�͜[�`c��D�D&���M�&�*�т�>��7���₴t�~��S����Q��i��~=��b;�}'[��f)hZ����I2�ϧ���_9{�E��̴������~@���6��o�zm��!�x֞��$.����b3����S����K�^^_'2�Q�h�r'#�>��悞V��呴k����̿P���q��ɉB"�4 o�M]b��������Iy^��ǯ��ʮ��B���g��+����- �"q��j�B��`h�}�𑡈�x[�L�m������֑��e���UF��\�G眨^ᒊ%ʪ��@p��	����4F��(��1@w�tL=Im�����D0Y�����K(��6�x6jx���>qԟ���0�UpTX@�pZ�Uoa[��|W�����ᵹpN|�m�3�÷���,�ٮ+"�����Du�ģ��l�-�\�h7�{��'��l|>+Q�waYׯ���,B�uxd�*�U�X���}����G��Q�D5OUߠ�7�dfc�FY�&>j�,��)'���7E%���p��g��]'�S�ߋۤ88jG�Н]�81S�]���]ZrP��9�ˈ�3;���-_#'$b�������f���%��t�)Y��2��Mm��w7'Gd0�،n��4p�[
�u�A�	բ�^�B�9��d\��^\�v�b�L|�0Sן����E�t�C��a`��ɉa���m�s�U5�K�r�k���?af�&�k�$�:}���.�i(���qx���?���CA |-�T ����}�5�Cǚ�d�A�͵N�;U���3��Ԁ&B|�6lLP�xI��$b��X�H�P��q*��p��7%�_7,a����Ֆ��Ȫ��VJ�Q��e����WL(���*��fզ�Ό��x�wSc��_��QQ����U��2��D�uɕnB�*��!z�H^��r�4�xi��K&j��	u�F�Ca��ʜ^�O�}�Ba�o7�Uq�a�KF�9�(�7��o	t�Jɼ-qXV�#�{�+i��$�R�ai�S:#���ꨝLh#�����?}���N<^ ����N�p^
h?���/w�a���4.vk�4����4L��}N�F�,�[Kc��W��(�6h!�p�岘u-3��|G�{�Q�[zk'�t]��4]Y`�
�t��]��\=P�	J���K�����H����^�Iw�FB/?������?x��/\���uSyQF���G;Y�$H�k=��w�lD�={>�6Q�yp��im��]k.<���3{(nJD��_nO8�f{& �"�Y���s�#�tak�����wH�z]�j��_�)l
���h��<O���r`��{�o���@��l���e���\���^<����\���_�R���0a	&��$վ�e�QШ�+�޷K�8�h�@b��"��H��?m� ���\��V��u��0uH�-�~>H����	���c�� ��*�W��Ow��'��鉿e5d�=	P����=a@Jq���`2|YR&׃�]8���ݚ���u������v{t����
������#�"�y�8�Xϫ���r�fӫ���J��"�&�h�}�&d(�W�;+rn�ލ� �c��< �m����KĕB�A���?��d�Ÿ�.�yM:*��C*@��/�%8ns�H�N/�����(b�,���J��eu�eo�Æ�B�Rr]�t��+Fe�x��� �� ����WX�~b��e��`1�� �ɶ�M<�ʣ�ӟ��/i��:���ebo����y²�E�v"�^�(3��/��G�@ɐN�w-sE` ��������]0Vs���n�bKw��ps��¹��f��XȐf>y�l�lԙ�*�ю���FА�p����N�tU�53��W��ɍ+x�����@�z�a���Q7��Q%Ї�wX���]�Qa��e�=��a*@ސ@�-��a�xO���6D[=Se_f�?��2E�� �ӑ�<:>7� c�?��=�1��\y�+S"�x�[��Ύ�s��U���Xam3m���Ħ�Ї��9�l�*�󼍋����-N�(��Q8Lv,�u��g��t�X`-����R<<q�m����n{j���(�����G��\�B5��'�>�$��� ���=o�׳���F�+7�E�+5Q�i����@�3�o�Gz�{��|��v�^_Ok�2`��<l����E�Ʈ��K�"��_ߨáB���*���s��z\�w6�]�q(�#n=��	��&%>�[b�Ϙ�<ŞK8�ɠ��1]�Z@z��m����׉_R��ߝ�~�&Mxw�|D��Ҩ��@w�}�B�L����8� ��D�K��9v5�d��w����uh(����飉 !ӵ�����(u�b������([�fEV]�wq9��WD�s�=�����5?����� �Fo`�v�`z��M$'��k��N��$�%E�MgP���!��_��˙��k�9�9���#�C���b�J[S�`�TR5�AO�	|�`�&���t�����s�1������1&-paL��t$-��Lj\�2dr������	d]���\�"��hhC��!�dd\
N�d)�z�q�f4Ē	B�V#�Q�����S� �$Q[o4��K���P�c�=�=����ϋJ�q���9[����%+�Ԫ�|X	Q�|��U��3���ν=-��3��j�S�8ݐ��A����H�ݎ}�I��
����H��G>���ߠ�K�l����r�.&�s�E\�g��t�+�p�a
���p�U�N� .����M��s�+���d�:��.�(��U��oG��x@��(���-�E�-]���v8&O�������b��P��: (���w	����B�i����v�h��*�{6�8\��Ѕ+��O�2��'��k�hi���Q�l��1"�'�e��x�-�B-�ܝ!��^�%��񹱋��i��aTU���.�"<.z����Q�F��ަ�iG���$D�#�DJ��ώ��Y���K*��}4�yuHf�8ӼO�ꘛ4B�+���D�J�@����W��@�	���k&�b�M	�(�|�T���-U���%g�\H[Gy��y1|�T6��ނv�f0�]Rt����%��
�~&>��gG�y���'�U� �g��0zꡩ����6�_���,�`���$�9R��N�i�ySaA�#�Yk�nB���f��|aO,�xd�f/9[
}:h���!u;.b��ymD``�V�=�l�H學��}L��p�|�����8��>i�l�������w�`Y���'�H7�����-���t��9d�����8`�'��p,apB,��C�4�t��� �f!k�Ъ�y*�T�nM�
т��?姻c\ %���ϊ@N��� YNFn������*�$q���b�k��2G���ϣ�p%�L��2r+;��0Z���$x[������r���[|(l+���<ʸ���܊H�p���HLO��6QJ��c>�6WI�'V;�`�������}4s]��z,�z�,*N��o7���i���o�d�/	Ko��r5B�=Q��)\:��X;;���]�����`��X�Arc�f�Voq@T�(��Z���
�4O�O��Ĭ�j��@�g���t/V�nR�P�#���C�3�I�"��{��`z�=���7 ���cT����������B曌�����Mm��5{���oj�
պ�5H�8�A�G�h<F0��=���9��T�0I�K�z8G�<�W+M;��7�=ف`���>�1�.w-]���:]�
,�+uX�/}D�Gߕ��O��a�ejUQFFyK������\m]4e��&c-�T�4�'���\�|�������He�D��~D�#�2��y������u>�sw��-�n}��H�|-LJ����!t/����	a�pA�|��Jx�;ӕQ��$�E��u�L��,�^KG�K5ޠl]2�G�2ѡ�W�]���L�܎�ԝW�S�P�y�+�fSD���`d820L;9��>�g��Xrs�����	ܣ���Ɋ;f΢}�J�Ozq�Aށz� I=�Zy�	��7��݂,���|��p+��I�)���M���4�FzUYG���D�H'�����"��$�7�����Ӹ��У�lyX�?Y=��s��ԓ�D���	�V9O\� �&4x��ne^x�eP��� �^s�MVkzr 7�G� �sV�:�dX�L��@��c1_�79�D���𺱑|8����ǏE���$���D��2㫳��������Ҫ�+(.�`^���Z�q��xf����;��,�01�	��f�TJ�Z����[~Њ��6���|�2	�����ޅA3~����u[f�ļ��)�YMw1�0��<j8�j��|�/E�{K1��E�������=V�u߾n�b�0Ə(ee�S�֣n XH�d�	��� �_"���~?M�00��cY��ܽ	8P\$��\���no����7�O=�
�W+�ou_��r$U���!B�g�.9O�<<p�l�R�h=^�ᓽ��:�iUz����x��G���tTϺ�3hOmi@��w��?A6���&C�t��Z|�O}3��ֈ]��2(TC2����L
ј�"'g����+5;R��ŷ	��\�S�bl���}bD+,����~�{=�C~5�/t P�)�ʭ�տR�*�B��e�S>�;��ϻ�)6�2e�˟��Cm�U����,L��+:�ȿ\`�L����l϶�+�O�N�W}5� 58�Օ^A`X�'�^+M?铋����a7��:1�� M�16"6�*�Ǡ���|t�paL�B��[ �ac�p�;�Z9/}{����.z<ݭ� $����񹌾�DY�&ݱ�-�[����m~`/p%q�`���j�ȱÅAda����S�|=��u>��`��Q�X�Ul½Yv86M�L��iK���؂I2�s�>Daf��"Xiko��;[ Cr
��v�d&�ߢx�u!y��n�'ɠ�
��-+�Z��2pL�#���	�Љqq�F�ݒx�T-s}:F��U��������Դ�O�����:�A2�v�J���rE�����Μ	ǲɔ�@�W�%����,gr�s�8z��JW?(�I����o��0[	f4~:�zs�(?��18���ñ���i�U]ux�3�l!g�|l�-;'�`�U���)-��/�,�ʔu��7����B;��&��d����2e��7'p�z)��E��Jjw���Ztc��݅����2���������4�h������#?�'��I6���i��X��SZؿ&��s��4��`���
t-�K�ŉQ�#���a��<�~Nx>椮襎��k�L�M	t�h����̦0�$AĒ��z�J��^j��ܘvN��lE=3��(d�M�W{����"1;z�-�|y��� �W�7~%?���4�B57%S<�����/���
I��[v��۠[*.��;R娹=!VP¾<�������tM{�1a�4�<Vq�9�d��~w�q UX�7x�a�~��_.�L�A��X���F�S�!G� i�"�٩��m�u�޹�g$��6����X��#,ݻ(%���j�_l���Y|K�đ�,���ɜS�g�o~ϥw*H�"ťV���e�p<��p]��<S�7rh��70��i�^��d�;)�ݓ<	��6е��hR>�Yi{x�r��y��>��ngK�Ջp���@6���iο�_��D`�Đ��a��$�$�$b��)/��"Lԡ��Ʒ����"�<�E:�ָ���E)�R���.� 9 ��u	�,DFcgS��9��S�W�Hc3k���8��=^<t[X����ǯ�����8�'v^�S�k�-��v�}�V�5����9�/��C˂f�o?� �K�R�¬J�l�w漄��$���!�h	���֑M8�T��*"~��殕ZD��s��h�Ul�/��l�J�99�s�M�#���Ѷ����SF�p�w��6Í�=U�hT~�X蹈NO�kS�[_�M�[��7�|�-M�W�>>&�^�h�������Ph�����Y�ETP�O�}�`�A���]@���+����hQZ��������ė�#�֦F��/x��w�ʱs�Ǹ5+`�+Wu�
���D#
/ˁ��Uƫ�A6N$P5rQ���9͜�f�s���]5I��W������xc >��ڣ0����~U�  �b��H�J~y;0�rY��i�
J\X���1��d#��5��$�L0	z����J��26�p�J�QYQ�}IUS�e����l��a9C�9��x��������3e��lh�Q�]�a�K�V�&�Ndq��"�\�hHe��HwF�Q�F�zڔ�!��r�/�9��]`���~̶�<�-�j�X���A@�k)�4�i�t��W����G*i�Q�jq�=���TSu�cˇ������o��..�!@��^�.�nHD!��� b~8��|���*���e����d;h1;�P	o1�N|�O���C�g���S]E�v�~��R�vY�g��Ȝ�&��YWl�eq�OCG����Q@�B��񱀅����Oe/�c8N�����w[CJ�3w��Cw����JitĂ*����j�G�l�j��2�9j��������G�����߅���������z����C#H�X�2��s��m�n�};����M�Q�X�CBg�b&lg�8τs
}ZfQ3��������r�{"2i�!���A0�rڿ��$i�ϒ�-�{xn���JU?��&w*�,���ܯddtm�N*��Ta����1��k,��P�V�Kg3!%٨��� K=��-X�;�G���-w����!�9�,�O��NL����QՎx�O�|�8$�����gM����ѯU�!qm�h6%T�[6���k��(,]��>�~X7�ApRi=M��ޜ��>�Ǆ�L�(�Ά,���M�s'��:Y�ǡ�&*ǀ��Yg�7Ʈ�_w&�q�8kQY�m��b�@5�U����ƃ
�5fc�D^���-�=D������R��@��ع=�i�°�W�L@��g~���	�_�9k���8r���/���jt{���N��!vDF�t �yX �~3ni���:}��\�˽�XB&/[��"e�V���,�wEiO��\ȟ���� ��8_-,0�͏�.�#�7��x���l�̖����s�ө�`SܣXk�p�j�ϝK�mEvo��ƫ��F���ig6��FKSB��Gޒ�.�b��go*�Y���)H�C����K�	��\��Q�����=����*p3܈��s�8�L�}5����/��t	cq�,!��Q��̶_���/ޣ�-���&A$��0��J���V�Y�5�bW��eoS�p2o�C�\2�{y$,�MF����|whCl�`
�0�ȿ�r����������~�։r��y�H�D͸�Ғ���ƨ�wiɊ�Q$�g�
�ұV�*����r/�ߦH6�SU�EB]$�tq^����E�8Ĭ�_��
�r�ހ�����D�#�W�)ݳ�ej��e��e��3���"I�E]� �i��oF������=/Q��K������]��K��q�-�,jQ*�&M��P$c,X��C�f��ɹ�>��\��|�mpA��0	)�n�j��ڽ�9:?.=���Q<]�jJᅢ��{��9/�^����0�̻vcv�r&��7�)��2�
�"��C���m\^�y�fV�w3�ڽ5���	�O�w3�����-�����V���$UJ�B�_�t��+A��|O�~��%~1�Y���~�A�|�k=;�^��w��_�9�ptP�"�WD|HeI&���5��Ǿ�B��+���CmP2�,^��'��,+�Jʏ[� ޙ<6���!)V�p�}/t�WԢ��lZt�-r~̚U~u��lf���ю.=-5���wԍ�(�{��OΊV���^Rtp꫿�7WP]&�)��'q�l��Qr��D+����q*W`��%+�
9D�x@�tc���	9�[{�>Wˑ1������F�W#��>���c�xDMy����H�8�܏Я��hn�	��99���|m�&��ð�0��S��q:���q�u%��?קPz�v��}�XBW�;1R]����:�kZ�����uy1���	ġ:��C��ގ�$�S��T�E?�+���b�(ۏ������j�0m9��
B�P���W���!@���/l��)ׄ�}j�-��V���	AI}��2|��0������a	�vn0˴���Ԃ�E�a�2��8W�)۫��[�L�䱆cG?(��8�	E[RO�2p5���_��R��r�[ȡ�Qk�0�ew�H� >\�5�n#�7_?�5P3K�s]���ib�w���]�M,�#��1u����"$<،����f<fw֔ߵ��Hc��-c���< #��wC�x:pkǑm|�B��%g�Rl��\i���4��kX񪼐J�px��P@*Iy�(1c:~�WlS�����\�РR�팝�S%<Й���>[B�ޫ��O%XIs���[6Xhq�IȤ :����J�[�#e�&��)�k��+WSiy���Jbʧ�OO|9��'�H��o��7~ܱ���E��pNr\�V�4r�m
��z)����w�HU��$���I��4��0�/ށA5r��o\#IS��q
\�3�ү4d[��xDS��e+�!�gZ05Oŏb����@��)�к�M����s^�_�A�c�0�_/B���iQu�2&��08(!�տw7���g
:��^&��P��āYx�ɘ�W!Ӱ�<��Fr�-��X ��b���ԑ�p���t��f�V���5E
�s��yO~8�g��M���p�~8V�4ф�Th���J��RJᇿd����'�{��=���B�7T2"V�"%̤�{if�4)u&*�Ȍ!��.|�JS�� �k�uOf C!x4Bwbk�p��K���N>T��55Y���@>;(�	l��>׫kB�yT�&��ˈgu��=-���zLoZ����W6�_�7ǵO��ck}�Q�ø�5}�V>]_AR/����:��4�:�d�
-��f�6�N��3|d������>�����2�{�n˰�F���O��.�ܨ��a�<��X2�h��P�[��O]��Hq^�uw���ol�pZ߱�∫]��rz���;6�+�Y��JS�ұDF�Dy��vd4�\c��@x"e?��,w$@?��,T�^l�~Z
%5p���vM����a>�&�hgt�8��p���R��U���_�3S�t[�1�����,��~]��R��@3�ƨ�D���+M�<�r��N�CS���UdZpm��v�ب��g~�`e��D#�HIchH�z)C#�\�?����������,Y�-Q�HLC8��f[��AWX�k�JO�?�X=��	�
R2óC�C�b�㕦��a92�ъ�(g��	��B��X�����]���7�,g��~��f�LK��s��O<C���b�#t�w�|�f��D���Ӹca��)�PZ�A������I �����\�`�3�
|O(00���?Ii��Q�	nV�Y�簩Bkp.�d*�y6�6;e9v��_J�j"����sp��i�R;�3H��	J�R��8A/�G_�:��	�}ѽ-޿���ž2%uά�` �if����'ix��Y!�τs' �/q�>vV���Jb�����e
dO�:p�_�k���9����1����ac�Q�a��L���D���V�4�FD�z|�J�-�v��;z(���#��Q�	��C���6���힅z,k:���$�e܃����#���۔ �'΢i�h�i�?���T[�#e���x��M���%���J��p���|(�� ������$03�k8�2t��c�Wd�/�G�S�m�	rV]�1����tO�	��NL����Y�f����LNF���J>�NyBv�x��.�|�.���}\
O�Iyج� �tNt���3L�4M8J���/����'�ƕ��0v��a���8�-qe����+_2M�& �-�_�Hm�[ii��$Q�ȍ��|��	�c@E���C})QY� _�@ĳެ�t�Ĳ'�\��\=2k/�!=��e l�&��
���3�MI̢�u�`���6�P?���&43Z���H���`zX/��\�M�V����������dej�A�<<9ml��Kx��q��[^����(}��&���r��a1�W`K֭!��@Kz�Zc�rҩ���g��է8���=�mk��M�� ��(�g��9�z�A)��p~ Z0���>_��mDpm8!I{�Bu��+�a[ܣ�2.�����q	� _>���>���Zb�"N/��|�t'B���pZp&�M_��-*0�͔TW
s�/�R�������,<���XOV|@��<���5ꦄF��p�����]���[ղu�V��UҳT=F��s^���x䍾�4�CK��6��.;� $i^N�Ut�'L�*؞��Uh] 4�>��kx�n�:@�K������y��>�"�:	�����׎�S�ހ����znC�`��O�?Bf�7��#���S�O�\�GP��"*�>��Ԟ�k�t`Ϣ�l��QDr$�rV�}ٛuP����u� u�ma���眃"��v�=�ڥ���^�`9*��m�����2N��4r�,VY�ט/�#5�#��(�T�!&XL�ιM����x�wzCɩY7���Y�BfP�A�d�~�x�}mx�)�t���#Ҁ+�,R2_� L;��4����޵&�}GC�i�7T��g��\G���ZK�?��;͎�?.�T��'�����E�%��B�/�*���P�Z��$H������6�T��m��Z��Q!�����یK����r?�l��	y�KЦ'7ɿ�І��I�!1KP�V�6���^�!ua������^�Ȉ���[�^����ݞ%�u�t��	R�dj7@�&D�^�3Уy璘!�|	�p������[nY8V4̏���_�:��ޛ�T�ko}�/Ś����7�w�h3R���~N�:�ז�.�D_)��"�8�e��>%ds��� �!��'��[�K�6pfhQ��ǔ��'�����J+W���}�Ņ�O{UilͤX�M8�):�rh��S�M�d��-��FJϞ��ī��j��/���#��F�������F��07�a%���N������0�M���r,�:�:ȨmΞu�sT�XvMa�Yf��Χ]#\C*�Q>��W/PF'���qD�yoP�U^�Ō���ͤ_zF��#��h��P�[��]��Z�F+�A����ޱ\Bi��{SH��[�\bĊ� lhm\�h��l*��m���T���Gω �4PXH^-0ic�L����{����d� )��^�5j)#�c�SxX��N`Q��ǐd�{,\ d���z!�h`�<.Aި�K�ּ�h0��h�z��^2�p}�}ؗh�K���X�x���g�Ֆtq���p�_	���.q��C��@1��c���*�)A�$�j�F�Y7���O��n3��ЋV�o{��mw'����amX�9��+s&��f�M�<?z�HH,�N0�l˗R�ږ�+�{]���ݡ0=��8��m�g��`n�n��b0�s�զ�	�nQ�#HP���-��CJ��>�����~L�X#h��DD�e+��{�lc�a���뺑'���7J��9�o�0��7��C�%Rc�r��v�]�n3L��	&Zs�Ef��!�o�j)�K�f���^�Z8�ͧ<(p(Bk:{श����U����V�F���B�8�]�m� [����#&[BDw���k��$C�g�|�D?����l�\��Q��3Q�4Qd��R�Fֈyʁ�'�+hyW]�����P�\ԓ�ϧU���Ƀ(
�>��I��N[����7��Q2�A�vn�+]!���5H�f�T`��� �­���Y���K���	/��*�A�Rk�"Z�O��� ���}�pY�AK����dV�?�`��R&:��<��X3��3<̀.���*Q3@��SwlS�݅�\v������:� ���s�=Y��r=T�����q��t)&Z?�H�h�E�������;]���0��O����P�G��Q����s��Y`zX�6�/
��wN =|C��ocT�)Bm��B¡Ҏ��f]�+�҈� � �Y^�M2~�c��s�A�T�VT.���=�Ë���OueCJ��+�^�N�'�Od/����G��b��W봤��!�/�ԉ�ds���qvML#��E.>��_k4�l��"��m^\Fmk*Rig܅������� *o���΍�]"�D���HX�)����X�3p�뷈_�-;���{5�vkc~L<g0�;u��=s�G	J�ۖg�'Y?�XB�#��(�w����m�$Q��0���P
ק��Z6�E�����s���"��ҧ��t1W��$/��q1�N*_ ��c�^MF�z�5�'�p��j�*�F~������36	W��)4�������<F�X"5����W%���T�+�q�<��G=�!�S
�6�~+���x� ��'�$I�X4��ǵbL��:�Z�-�TFѣ���mܱS%a��%���V�
�,4��Iڔ�F5� �́u:�c2A�D�퓊��{:����f$�v3{���K�o�'\��z}A�3��DnՌo&�ƹ������|.'���=��?N����\i)�o����Z��*c��Ee$5���a|s�P�?�V#�}�1�G1�ᚑ�>�X*zY����e'�o"�gC]��D0�����g�@2��k�#	��W�3]ďAp����1_�҈$���$��x��a��Z�yy튟��tx��#��{߃���v�� ԅ�*5k�y$-WxG9��_[�����:*�gԌ�����"i��[�z�LJ�*�����ٻܔ�� TK��k��To�㑃���y���k� �Ş����z�ѓ�%�'�c*���GB'w'��z�J�ۈq:���q�O�倬k�ў[Q�0������|���,�A�;����ĳ^�0�@"�˪O>��� Р���]�!P_K9�:�(���'���R ��y��G��߬I�F�hɰ�3�iC0�)��'�MPMJN��ӮL�qQ��B��;���3�N>F_�_+�+�d� 9�݇Ʋ9�s���o�=������]D��Y6����J%j�)2&��'��tZ�
����׽�\���WU�4+�R��O�
%aW�9�(��gptu�!d[tޖ-N^�.(Y���#�V�;,;I=�!'<  �S�����鼵���|�\ 
���(���JM��K���9�W����h{1�ӓ?�M(젂����w5,��'xЭm��β��J�Z�%{�Y��K�Ѥa�n���X������h%��o�&��$y�F�p�G.�[:���y��z�Ajf
6�w|$��l;�eٍ�b��@�A���&�!�,��Wi�1�e�X�y��f�J׶PR������ޖ�KH�< ��w�i w)��Y���令=	�U(�os��K}��Vc�IZU?�V7v���x-~���
��ʮ�}����y��6Qa�z.~��*��>+��B���x���4E�
���-�x�4�S��`�X.��p+0?���@\�Vqٕp9�7u��:�on(ޡ�o���ZB��| c/�{�?o��
z��S�3���D���:����9���Ŋg+kl���bj��^���'� p���*�X�奏�A�?����:7^r�a���j �C1��o+��S�D�ǙQ��ԟ!��_Vz��$i������]�����P�r�zB?��\��%�� �nɋ��e�q�2�6�3�-�� Ux�z�.��7���r�˨?ue0:��z7^
�PàY����]:�M�i��%V�>C3ش�����n`�nR̀4���ȴ7e=�]M��N��y1[G_�;D�Kg��S�V�ڇ�3�&��"�qp<$��%
��hug��Sƶ���fr48��P]qGRyɀ{j�"���۱B�#ʚ�a�ru��-/IHVZ��v��#W�N�\^j�<�J�V�j���%�[�@ԸD�֡�O9�����j��[��d�d���N�FF�r�>����+��q$���cE�/v�`����T��xd�e[ �t��AZ����&|=L�� qk0���?~�K���`���	֊��,����֩��d��k�V�\'�c,���{�� ۙ�� ���^h�_�{�w��7��^Bq0*�Q"vg�ԪƟ�VvKS��M���<��D���Z���v�4:p��QAu������ޭ�	#q��P�41�;���v)5s���]������[*2o�@�SۡWK�z���l�U8N몔�7[�[K����+(�pa9q��^#:Iu��B�;�(G"���ᙲ�3��X#O��,:'/()
1N�=��³8��3vr����/X(�p�����A�N2I��<�'���`H���X����1�)h%�E�(xIG��U��ʌ,r$��6��,�y��; �Y4}�7�+Wo-c���t�y��Q"Bb�zyU�xNօ�\�r���4�X�H^9qE�]�9�+%��Z��^s��Z���� ^r51¡5[d�qP�N�(���Z��;5Pn�����F[��������������Kx�5���bw��������_Χ�,4�<�
Za���{���+�}w,¬ҹ�yeN�;����I��s �B���X!i�S4L�� �K�g�U˃�Z5N�����a����Oo�䓇 ~l]
��T��������d��������R�z1M����^����;�Z@���7W"Ş���~��^4:�c"�Q�3�(��
�z�4�3�>0��H��^�y,bIS:Yy������Hu饆A_Gt�>�����[ͬ����0��[��8�<��60*���zS�˸,�H�`hηmZW2)Jɷ�p��E���0*	L�/����������8e\3����P��W��t}��p�E��g�M�2ss@�*x��a��H�)��E���X4G�Vı4�˛��!�´kr�ӊ��rzӗf/��Y��ux ���a:�N����
,m��M'�
6:����[����_9�n.��ł�%�@�b�]N=3�g��K�^�~� ~���}p��r�ycSY�l����8�j�kϺ�������^��7m�Mk�Q�o�8o��Ɵ�

��$�P�rYP��莼�]e�M����A�q���~-�.p� ���})����bŧg���	ݩC�����(~�g��I�bC���R�0jF��$>�PT�	�^*͚p�� h��G>oI�s�������*��� O��h�|���^n�x'JQ�I�t���t>�F�\���qy����W&�@�#d])P��#a�>��e����&X�,�����+@E	����yEJ��=f�9���5�'�{�m�T$�&Ք�!Yf[��g@L�M����:Юu��Dݎ�]���O~�t�R�
I��Z�׎=�w�4ශ�'+��v�R}��>!�GB�2+�xC�6S|�����ˤ��~�[�Vk9�P<� ����=��Ä��#ԡ���D��gs0 ����';8�Q��yV�'F��^x��B3Qb�P�oA!�i�l��8��	�(+�� ��|:j���k�a�y��c�kKUIp(r��H��G���O#3��>)�{�#�B�x$;�>� �Rv�Lս��8=e�U&�UlWE5$(|Sv0��q>�[�H�6�!���Ax%�����F�&<�������Q�N�D�X�>���6I��M���vNhJ��;{����A�y��2^����u��&�3�cw/��F���_gvkP�����f+%M0�1�iA�����W�;+ۨrmЊ+�P�t�����p��c���l���+~��"j�m�9W~�_@ܔԳ2�����n�:/��l��E�k����ʯ?�Tg�1�x_������$�?�{��`�������~�m����c>x�{�x�.V,����3�"^�P�Y�5�(�C�j��Y����F�K*�se�%wi����ҺJ��ϓ�Kn��Wo����M��]��`~w�#<ߕ�&��$����`<��d�HO��� �f��4��D,�S���ױ�<:�Y>]�9��qV��.P׽�$7�����L(s}�k/#�F�s�8�m�;�(x���Ya�bfm��R�E
^	 ]U�B��=�3;_����* ��d�����fL1��^]h����{�������tQ�Ӂc���p�����ȹ��)t���I��rLd&�\���ι��0�'IUN���ֽ��+���s뼨����AC�@�)~�-W��C�D�>,y(����zcV0�t���g�
d�A߅�!H斔����7�{]nn"�ln�W*y
�;�|M��� o���������
�E��(;"�B28�Mpq�W�������
��D��'cꋼ;��u�K��O��&�g�����}`9�c�W1N������!h�I�B�7Ɖ��$�/�׶g��w���uKB��1,�#3�����Q�<��@�g�ݻ6w��u+M�V���D�O��j���x�f��R��Â�]x2�X�w�w ��H9�z���x�+-�Ryب�D��/�613޶E��$u
�]X&�/����Fڧ��3s*���g��� KaC��.��ӽ-^��a�O|^�*f��G.��o�PLK��Һ��)R�F��}�7q��7_��6|�f��
�E6 �[g���J
.�8�
��+�w�G�[w�=�9��$=f�BDP1H��
���wD¬! ��Rieәbm��z��>�,	�5Y��J�Y�\;�m���z#�Qg�m)�d��h$VBJk�*����	R}�|�9�g���_2˫����"�s/g��ni�_е�W0�(n�v������&����Gq�.�!��~�׬�5�u�i�-f�D�JY8>�{���{[#�6�?�G�6�h%��E0��Hp���.R�Z�s���;�����_<�Wg'���|�b�1P�_�� 
8�TL��s�s�X���VZB�N!`x;R�Ia=��@NoF��E�C��rYUu{=����X�G�IO���Ue��f�>���9O)�QhӇ��ؾޚEqn�(2��<�`�
2�7nO��2
���(�l`ލ��*���י��C#,|��
Z����*�(��m��k��
��S����H53��@�>�f�W�skd�8�XD���o���w2�Z�r�M�=-R"�X9�;�m�Vg]����C��g?C�#��C�8h�tǈ�Ns����P[G?P�|;�TA�P�o/���o���;��ˡ�+X�}��������'$sF��g��/q�d�ǭҐ8��T�-d�cd��5uL t_�E�5m�.{8�d�y���C�8�)� Ϋ�cI�F�I�dal=�.�``=%{���om�*?��J��%[�Y��Qb�Ƃ�7Aʡb�ڹ����) KOB�`�<l��D�{�5���|���N����%�+8�-�.�7��jXs D��
}�ˏ���l�6	L��3֜�<����xHrւs[4T�ڮ�⼦~
�#�*9Z�x٩'��N�ª˥n���-k�p�wo<��}�p~��7,X.zxG� �9=�_�vZ�h��yv�gR�����Kz؋��Yp���6MIͯ��]��?�Mk��Y�����OOi��
�<�.iw��@�J�G�!s�WϿ�,f�e�*:ކ9lHs�Z��ma/c4�|H� �G��N�w����3�|]�"v5�O���hmKm�K�J�Ǒ(�˫�U����v���#�r&f�����<�졵�i���ݱ�j�4j8x�K._�-�J�� n]{Q�,-��P�a"���5��ql�7��w����+D�~ �����O�a��1��~Vi:�~�s�x�6h����0:�4�"�Ł�dgcɹ��K�����V�C�OtۻS�S�����%Si��<���)p�� 	~~��r���s�v���ɢ���������I��>�R�nE������CR�ܪ�w/�ь0��!NP�
ZR�d���%qf`��.-����2%-ơI�s�:ٖnI����s�
L��5��-�E�$�(a�ǣ��0���=��W�����,oʊ�������{N����2��j�R����T��#3��7�r)�5�<|�cN���渉`�VJT��D;轿L~=��p��S�t���i��>�X�ot(��UJz�� R|a`� m"r*� x����ҎD<��_��1v�J�pMf�A�Q�}��=E�}li�o����';^��i���8�1u�on-�	h����6(!4���P��94
'3��_	D��~�!`n���dp=C�_��Em	c�o�52��W(`jc��h�q�����~/;ZL�NA���;���G�,����c<���'�� <B@�3q��Ğ�N�-�96;�(_��ʇ
��I����Z�t�J��JB���Dp��K��W�r��kF��+����tԍP�!��D�"��M��>VYe�kc�vݚ���(@\��d�:����C7}	w�s�����5x[�5E��g��߬D
�㷧f!�]	��O�$�D�n|`�$#���J�<��w��c��V~6�>��^ѿ�R-ٳ�9pO�mg��X�Ko��d��;���0гs��.�n�����C�*�@ƓE��ʋ4;�������JW��?@h�%\ ֩,`·*p��<Su�gL�ﻤ�>�Z�4iཊ��[9�Q+@�R<FVC ����Gc��lgM�Z��/+�_�ǆ�IVjH�T$T!�r3����M�đ�s����m�W���4��D���P�*�2�}r��z��s��_�o�,�y������"� m��oeAp$��o@?F�%�1qa\,�^PZYU�"2R �aw��fe��e���]OZ�Z���}֤�W��g�+�;lwo w��b����i]��2��t�79Ρ�,�iȚ��;=�R�CP%�7Vk�H��?�w�#.�%��mhߐ��q֖�Wl.��M�rF���>�$�Fe�\&ys&����7˒�T	��?���_�odX2"y|o/�[}3Z�[N<2�SɯR�~G�u�z����sȫZ����O]H�6C޽7c��o�(�s�+��l�缱�=�ȯ�ǉ�N��C��=�k�z�r�~|�Z�ni�o �C*Smjѐw��K0����o���A�^r�v���!2��ϐ�+� 0�˧ޗ�����nm��0T����O`�^3�F��Rg����%Ԋ�?U	��>x������I�vukJ�$e_<���)x�RB������O+�����xp��=��|�M�QC@Gׯ�PaX�ş�qP���C�+
k�.�>����WW�T-z��rAx2a�~��k}̀�n�EpW�@�	��?��!
-�,�̩#E!`�*�����E�鵕f�R��G#���q:)C�SӾC��3\���b�Yq�2н��E`s��@9���u��n�/��Y���a�P�`ݯ��>PoG����{>���J{�f�p��(���}~�����������^O�mc:`��o:v,le ����X#f(�S|���!9 ���gE�-M�w���u�I���ܖ{Ps�~�D��Uj5�/�yԕ6~M�d�^Q�D�A2wU��ۮ���E�+Gi���YrPk5E���C6��8z�X'�Ջ�=y�s��fX��4-� �=$�Bo����k��e�:A)��?�3�+�C��٢y��Y���ـ" f3��ee�:~#
��{3�L�fv:�eZ��[�ݝ_љ�j��U���FC�`Dw)�d
1{I��
�l�@�|v�������~�|��Z;"����Ӂ!U���i�]����NR�m�,M����[b�L�4��Q�x���g��t*tǱ��Ԝ��q��X}�7����|LEҊ���U���<+�}*�@l��������o�KZ5a��R����r�~�V���^l�o�:>�����-��D�#��!o����<�3�2�T
�3�|&Q"-u��R8ʘ":z �~���1�� F�S�>��! nD�A�4�~Q�"f,/�K����OIm�Oq���E�����K������ZWR �U!�B�И=��rzt���n�#C�E2V�ދ��!��b)z.��<<ʛ����%v6=i����
����d�	:��k\~���9�+Ar��Y�����l~���Ɵ>�7�
�Ԝ����EL֨�Ea���ի�^ov�������7uo�M�e{@�!��>�9�ߒ�.�d$H�;�8ʪ�P�Ď�QU�!z���Q���F/"���c�_l�[�Yv<��@ˠ,�g�f�>2��R��ϝ^�sP���&�~Ֆ�j/0j��N��Ls���e��F4�Ǌ�����}RJ$��Ns�w-��lc?�KRӹɦ�^�I�x|-a�����PA���됎��"�w�)��|�R�P��m�Xt¡\� ��𬛜8Z�L���y��&d)Y�rI���z�GUɅ��1��HmL�p'��{�e	�p��-�{��.�g�)!?���k��I�Yƻ#����0���5U�����v��>�3�d�S��{��ϣY4Vn��J/dG�<*�����%���h�u���eu�z���Q�c&�BM��qrZ ck���F�V��}2�h�@"�����h*W?����|û5f��zzzա���~��%���	���X�G߂ϟ���P�*����Zs���%`�gE�YD�&1\Z�C�g2ɞ'������w6���;/Q�+FD6\���L�$2`���U���J��'�&�#���E���V��(����������ё��w�Tq�A�4�P(C�T�PG�hۊ�v�T�m���8��1q��_�-�k=.��G��܉���y3!ϊ�NJ�1j7���v;�!ߌ��{i8��~�C^r�I���������񕺥�Å�"J���� <�b�"4�g�s%`t��;s���pH��V �3jjL|�X�������xC�2�)�ܧ�2��>������4�%�ml�߶s���r���Z�G�U��2b�$@?��t��UFx.8Σ��]�R�!#�/�8��/�|���)���T��%�^�����j�W����؎�N�x��.bX�A���}��m-M�,���eO���:�M>qU��8�8� Z j��� (q�*�BrncX>
&�C�(��րd�����k#����r�����ռ��J��Y��ό�&�!-%jiX�9��W)����|�����s+c�|��Q�O�3��Hӵi�^rJ�΄�[p ��O]&b��#�����b��m�	m�/��\�)ң"ΦWc�cz��	��T�@t
:л�*(���(1 �(M�f�Ӓ���# d�bH!��[�}�{��`���+����k�S2a��
��rx�>q�^�*(�lM��~�{^9�9�������6��lk�n�p��F���T�榻����;����+��r����l���ξ��o��_@3�K��N��� �	w�^9[>."h&��2��S	{�ho��1����;̻�'�ʿp�|/M7ݑ����~��)��'^7�\��X��
ԍ}U����g�D��..��
�wUx�{
?| #y�|�f�RD��_��"	,��%(�V�}0F�J�'���uM A ����/��M.�!��HF;~m̭=����{M�V�ݬ��	��f����84� z}>X�ys|34�$�*���1�A5�������`��v+�Di[Vn�Ҫj_L�9z����D/��nc�?h��{��X�V�~^Ȅ�n$���-��>:)�yU�N���(��)P�ߧ�����d�6����ݏ\����e�ڍk���@�����6�9��������>�Iww�%�4����'��>�c����t*�X�qQ7�(_(�=�Wpõ�z���p�u'��(����W�t��_�q�<q�5R9STal�uE�xxϋp�ϻBO8�E�(���PE6_\Т��^nj�/:[�J�����\�ͳq�`7�Z't��w��uq(r��}C� EZa����QIZz���Mh�n'=oH�m��u(銈��"��(^��z����C��Ǫȕu�|l"��U`A�_�G܁��ʝD�Ȓ\ 9�ϲ�&}���}���D�H�k���\��+���g tvSu���i�C��f~��O�y�0qb��#ɀLp���J�x�N��c�cz.���a�2��c%�����B�M�L��;����yh���h�KKY�˴ߤ��`D����%X��h��M�=>i�����T� ���`��ٙC��q�O+O�g�^�����h<(�&��Ԗ�t��.D���Dߊ���.Q�Lrַ)�I��w�j߹���3�
�k=E5?�V{������=�*�9c�s���gߩ!���+k�	�l�Oj才���#�v�b����������ء"��2������Z��'�}$�u�kĻ�^d�?�R�;�LEs�ÒD����q�aĕ�}�3��ڽ��?���*7�С��
.
Ap��_��r9'��z��k쁯}��~�
��W���(��$�V����Q`�?p�ԩǰ����iZ�v!��bl�8,,�	��J1��܈�#��y�P��#��>����(���7��]h���d�rʕW���+/Ɲk��I߽�R�ĈK����%h1�F��(�(�IVc��dI�U��̟!�z'�	׵)��W�6�fmĨ�-M�K4��}�!���/{��G���qg�pہ|�0S>�p�xt�6c�H��ҡ�*�5�#���M���ۧ���i���\�z�E�0q��ȳO����	�������T���%n�$*��%48 �W]?��X�:/�v<:W�B��l f�!�J��w�q?��V���l�Hs��� ���}g�ٚ�')����8[��B���V\�:a��N ��k���3�w-anG@�&���T�������i]�k&� ���&a�\������1��L��j�=�V~��VK�XM�I���܅��'x�èuP�e�%B>�eXU��S����&P5��Iز���w#�b#;��� ��!F�\�g��"����ޟM�
5C���,o�e�F=���~�:�+	W��U�C4�C���Χ�_�$>6q04e (�l�\81�GZ���C�?��
;��Y�gNB������R��Z�b� ��ƢR|�<����Pvt�\�~����'�xC(Y�"�7 X�H�c#�]�T�St�$����ۖ^9�IK�8X��i�����EA��`��{����O:H��XT�6jo��Ux$���"��seo�J{��w�m�N��-����0�T	�����o9��;�k�2 bHw%)�ԇ�j�_�Z�T�R� q��,���Q%P�QN��H���'�J��wЫqox%��S� Υ�H��.�=-y��n�i��p�ޱn�rO	\��W^�-ju0�F���;N�wD�		�R.}/LvY&��@,���6�ݷ_��:KGZ��K��g���H7�����N��K��ET�|:~Jl,r��b&֘Gs�@o�{xN���IpΩF�
?�S
.��L��������G�W��+\`��R�V=$In�n���	KVĲ�Q6�g � >[�l����>J9;�	u�P�O9cP{��k���a���阅�������[����_+B� "I�%uPv�Q\���� �z�ʛ	����8I���:�ۊ��D�B'V����,�\�.��ǂHl�.J���(�?��f�l/Y���Q���d��הXs���p�a��Vg�����M��T��_"m��`���@h0ް)4�
�L��%�Yb�H����j��|?��ܜ4��yX�����P�1�?/���z�E�9d��RƄ�Et�c�H��>�ޯ��BrY�G��ý6�m)Z,�k�X��9/T�>�F��oy�{�j�6�eTӽ��`m-m�;dR�����wfՌ+]��(�{�P��0ʸo�F�^��H��BJ�y6i5�g�2s	�ݑ-�N��$�GϷ�!C�#@��^�.��ʆ��eչ�u'�p�J������:��<������d߉D��}����{�b������JC���b��(��F���C��wu���/2�/S���>;�*X4���Wڠ�A��\jz�<mk�s�}D�p���\�^��3o�M�)��Q�0A�S�5tF�2���^��P�2��6D�CF+�RC��08�U�l�	h���L���@A��ޗ;�DĊ��q���n�:1�M��)�ChH[�fl�����M���y7�O��Y��J�zP�ucI:ѠD�0V@X�~���C��S�syV��QK,�!k?'����k�!6�j{x߯���ק���e�ʘh��1;�d��耚�?�gߥ�5�'�xz���o_|9�>��/��}�y�.���7��|X�Db��x�˕���<�v%X���s�_=l:�ٲ�+y�c�/�t�ө��J?v��P�l�����lA�Y�<����^�,0���Z�p��]�
{r�w��>��8���@cx>o�E�y>�|ٵ�� hhxo�$p��@�
�Ү<<������5����5m̀�f엧$�	�Mp��a�2�ƸW����u�6��^���b[9��a�&��B�_��N��ZpC9��>a9����k��p�0�B�e䧿� ��������#T���.���O� �@�;�D���It�I�r�f�<z���e�}�X���- ���P��z�������/}P�0(�D����bPH�	�O����hB0�&!kB���/�ׅ�di����V3;0,xD���u�����}9�2�)]�|�&�rX|Z\ļ�)t�4��.���u�$���D�N�����ɣ��g����vLuK�j�&��_2;§e)�<�7���9�2}�xc�:/������n��i+~2�Q]�\�/<���r�f\Zv�cZ�^�E�r��w1&.����\qy(��C\[ҥ�����n�f��x[���"�X���Ɂ�)'P��r�\6�E�{\A5�学%�x���-�@��Xmf�
+����&�#p@ j��2�(��8�<W�_EO��0|�:�V�{�p�X!�8:ł������oR�SS��p*\�s�����x���c�yo������N�$K�'B�44���J�JU�4A\ra��w�{~2�u�4\<��B��G}�m�1����d9C�<{r�������Az&�^�n��k�{-���K��_��%��z��M?b����s����
 �Q��5�e^�$ZYp�C�-'ٓ�=���Je�G�gLX�Ej��.�\��X*E���C�:���y�?Qºl����d��*��B��(ǣ��ܻ�Ñ�:�"��MZ����R�HE��֬^0��f"%�G�pWw���(�-Ar����V�3m�	���0��I+��1��=!�'�/3�T�[��"�R� �X-�X��cCdW���gp�)��ՙ��Xc�{�0�h�F#z�N��o��9���CU�,C�q�ȷ�-��=�L���)�_�54 �q����K�!xq�B!��%o�t�NVcR�o&�^,��w얕 �+c+=�Г��r Ԙ~���uZ W�~����>�/^`O7A,��7ߤ����J�㷖O�oR�c�>W��>�H�l��"�H���ڙ&��n���bd�2���͔�	������8����{�/�=�H��^:���V�7a��$��O>qp�*4�������ʽk��g����p�ܞǿ5�N�WT�\����������<�<!�8��B�=Ġ=����Ma���N�ϔ� �N1����$�"�?G���`㑀ؠw&.��x�ѫ��I
����	Ç���rx\�B��A7J�ĳ!Zk{{h Ç��h$����k[mJ'��Mt�#f��[cs�	+�w���vbu�������}��%��W.&��( au��q��ȽM��[~q{��#��>����t�o�$X�����#8e�@��>��{�{�]�����E�k;�?zqC[d�G��^>h�ɤo�o���9}6�N%����>\��6�5G ���k�, U~�h���� �M������`��˰�3���"<�]����n⿎�s�,;�h_?���/��{2�3����t��Ňr&�Y���w�6�ܿ��"E�jz�ީa43HD��o��Ӿi��Q0ҨL����<��x7�z��J-(��7���=?StMjX��Z9���.��hp�6X��B�Z����D�.4<!A���\� n�����td����G�`��)N�%Z�<�!}��^���e(���������|Y�$��n�w�r�M�U���J�'t��my'��疵���w��,̥�ʐeǾ�T�\��^m�Bg
H���/,�����d)�ă�� �<�b���w̸n����*D����ű��c��Е2s��-{��hH�U:�L�m����e���N�w������X�d�jm�/&H�G|N&��+~�*ˎ��8��!�?Ͷ(N���jy��r7�l7����/���HY����ժK@����()X���OLǓ�ĕޝ2�]WE�ט����0��v�E<w��"&H�	+DRf9g��M��8��\t���s�ZM�H� ֑�D�����F7%�0�|É�B|���ė�j��[Z\"����='���� ��3<�Z%���̜>K��;Cų�	j5��%Ё�
��Ϡ�{DƊ;0���ϋ�2���i��d�Z�(��g�����C�	s<-�GS�w�cKǉ}9M�g��B�������
*�P1Lٔ����O��K2�I���W�!ӫ�/�1�"��3����1�
Bc	�������^W����T5I���>�R
�zJ)���_c�� 및IC%vYV����͇#�s�]D�y��q��c������+'{�k2\�s*L�6��Ǘ+6hmUȾz@ ��3�fY�d�u�a�{G�V�i� 
�;9���?�Ӓ�t4�����b9<6�D�fH��)T�`,�h�sV����ob8��9	� �wm܀;EW۹��{�q�+�6���z6�@�@O3��&��e6��eUDo��D|$1��?�FLB��H�#�g�mi���S�0L�Y���7Dŧi]����'�Q��}����T�i��cd��i��{ܹ�����x4{��?С��$�6� ��(�tj̟�g܍�l�C_ް�O�g��|k5��Eq�~F>FnC��U��w� �;�ǃ��&pλ��#��̩�3���#��C�r��܂1���&}�NV�P	˥e��:�a�t���I�%��{ur��Ѳc����/�aA�ە�(����̖��Pc�xyg���$�:�G���W�	ǫ5ǩX^�,Ȧ�̩�o�m=��D�fH�t~��j�"t%��A�D��b�^b^�8��|����U[�@���,X��\�B��;s��}d]�����\bE��w��}vu;T����g�p���$Dd\S���Z㑨�ǖ�ءió�q�"�S�����IQ��j��qm^���Y"�C�ޜ�V���V걳^�	������}�i�5�|����>���| ��2�a��@�?J����AT���`�t7������*��z~LSO�t�6?k�^�[�g�_�a>A\a�$Z�K��Dؤ��j�^n�$�\鷲��jO/#�/�.,CV^@���P����ue��v��
_Dq�������,S� 	��W��N�teY^F���_ʝ͟`���[O����Z����ƫ�x�������/��D�١9��Bn��%;�����A��2�,�=��X�֦f��*�_-���(���n��>�g2���(���Mm,�Ӌ̆9�<y���Y\�٪��� ¨��]�Q�˵�/v��xL29��Jx�!cyA�Or�w�?�6T<Dhm\�2H�_�D���H��K�L-��䱉�E�����u���[��2)zc<1>�I�6Z�Dh�W�ǭ��Ԍ�}:�`'�F{�o���Q }+������٤�%E��.�
���U�ʝ��cv?¼(�9 ��zW��L��-]���m��H�"���.���QbC���!q��N����>a����k�t�@\�`�uV��i�s��Պ@�;rr��R��<R2&G:sz��U훜�4��N��!oj��FxOֻnu�}S\�뗄������F�R���OLGܽ`��[*D*�.�D*V�2��-�׋Y�O�
/�\���Li��SCan�,��;d�X鱎��>�����7paP8(#��+vʧ�%wCB��^�(��l�"�@�'��0�_� �e�2ˏ�T�r�2�wk_��F�#�a�B:�)"�8P}�|$������J������5��)���Dȏ�Y�t2l�$���ACj��>��������ԟ�m_��D��z�Z��n�kZ�c@k3>_Oo}H�{��?9Z%�*�-��h���ro�#�/RX�2�O��g�$��A]����Y9��@�e�B~����f/$��!
��tͶ�j��l�x7��6L�oGO��ߍ��9y�x�H�܏�$��ԬhI��|��\�g蔄���M�8cQx�,.���}LH�{a�^��)�)�W�wdc��u!n��vw��_&U=�.m��3��u^:�@Ϳ�0'�p��b�K��w�W$g�����u��Yo��I��Et��O���!�iþ�T�uKy�Yӻ�����#���>}^A0R��%�W#�7 Qc�3�`���#��N�n��ɽ�דB�E�-I��F܅���ޕX3b��D�]^ ��|R����J�Y�5U<?���\G��&���LZ��ϡ'�\3'm���`��`;͌�e�G�2����W09w�R�R�(p�R=����7�j�x��ed�>A�
��;jW�!���u�z����8d1Fԫ�1J��^��З?������4�[�{��ir�p�bW@K��J?q�X!��x?*]�1�t�jv��|�(�H^
���n��]A=�h���f���g��@����&5�Օ�e�����ǐpbb<E죙+4{�2ׅ I��e���2�a���~�� ����������*K]�~������XٶwZ/;��+r`G�I��Ho���29�V�}Ŭ�z�꾠ӿpٛ��E#�����\�`=ƌ	��:��&�E���L��Xr����ü��x.@k�ª�{�M��m���U��}Ec�B�������W~H����O*�O6�~r�d��C��/D-tL���pR�X �{@2T��6��%����V&����X���Ԕǳ��������+C	�)���������YR�`�_�hڛ�&� �n�U��_a4EnK�q�Z������7��I�:�'�w��ťp�Y�<�L����
2E��F��|���hFL��%�lL����6G1sh��иCz��m[���o�����mn�����$�����FIf�a��j'Q�v����⒟�C[ ���s�@�a��&�����f�BUs�	�y�$���.�2I�%� j�=����-<�H�^g�]���a�7�uDk7I6#��l���� F��!�7�3�cq�9Q��2�s���˿9�CL��X������á��Q��E��)L�̺@=�� -�_��1������ �_�aV��I��)���i#%E�w������`� ����:��|��9l9mZ��a���*���@�v}JRG�S{��z4����gEE����A�K�颤�\�}�L�?"�'�~{0�<�(3���hB�,�j�/��7e�ؠ$�Kc�/Nd�ɱ�d��;�˾X��LA�N���V�Rr���=��0wá����h%��*���TF���2<VS~�G�#���u������a�P�4��R�k�YW�A�Du����V!^�Qm!fB�b���#�'Q�/��$H7c�h��{i�׭-�L5�����#�0�^)�X� I�\��)P���O�ז�u�+?��l%��Iɖ�����+)ZJZ�,QVk����0ؐ�"F<�g�}�9}������C5��oR�~	��V��̭�4r[ʹu}�d��{�L��:㪮J)�7T�@4}da��#�pR̚��ޛɜ=fJ�F3%ɷx��r��Hi�o�� X��ĺ����_0�G],�p�y���J���H:����~]`��q���Taމ2�Z/�؄Ixt}c��$�7{3�Bq�x�i�-��fp�0�9�s�߻�%?�=(C��#�S��g� bT4��PFY�G6H��|��L:?�-�k�S�y`�y+�N���4c�2au��Zs,��Z4��J<߭��SAL����6j�0��Ax�J�sP�U�
����N�#s�A}����x�x'*7
i�a��#���y�����6̕M�� �ߪ���==��R�!��;�UVm� �����n��'�/������=��q�\�蛌�Ȝޝ){Pb?J�G�'�I����@g�,�&\�Z��K t���b�z�v�2vQ�9zR.��/t��}Z ��#�*� ;�0d��*e�*;����(�>�F���ȭ�i��;2�a���s�"��Me����ZA1k�\Hq=A��5�q���B=���{�W���}RT�ٟ)4g2Œ@_q���`���G��u�P$���l�^�[I�{C(j������G�[�?����(�d�D7.u~��g�h,.:�ƅ�H���`o��+�H���(���z1Z��2����=!~�

���𞬮��k��۹ʯ��"�
�EQ����`��2���>�"V�����7���f��>����^g�����Z�iq��]7(��2|x���zǓ����R#���� �H^y@�9�A�w�_��>5)�Riq��{�7�M[p\Kx���j������U��b'Ƙ/,��D�a��"|\����uǇ����gj�<C�����~R���Q�Z����`��g��Mv��O%N*�A��%\,/˱�����0�ܳ;1	�b��J=s��x�8����ˁ��=����Vm|T�ӄ���d�CI�5^�_I=��>�~+}�^��Hd�?_�v���u�#��Y�A5��\'L2h�Ԧ�Fީ�P*�d��W9�����T���d��ZL��nE8���p >`x�o���D�����=�8\/�7� )1���2�U��Y�R���/�s��Am؊��N�c���Z'�./�4-گX��%��1�tPn���xsZ��@˧5��):��Sd��Hb/���X�j܌S�Æ�������9Ϻ�����g#*��Q	�
��V�(G��c�pz6��D�䌀�� |ub=&Mf$�.I�Q&�r+_nN.-��Z�a��ɪ܅�
nu��&ڻ>q2 �?~)+�A�N�HC����h9pG����7w����S�`jI��Y�Q�;ѽ���I�:V��?��v�K�bY��K�G�`i��&@�w���ׁ�Ϲ�x�@�O:�t�젯_E�eJ�ty�]��(�?�����=cpB����ǵ�����<k��IG-Wh����"f��,<*w���d��x��>h=k���ۿ8�K?ZN���H����'���s'��T�D�N��i�y&���5�!|�ȡF��'��FLώ98%��;��S�i��9*�	�#��Z���x��C7ċ��i�W�r<{�����޲�GO�fx�%��&��q	z��'
�c�B���_��n�r+,��t��/��3G$���b��O>h���X�=�>Q
x���{f9"��W7���@�U������j	��o�x�����"0�T#��hn'
����@^���Q0Oc�q�]9�(�I���#G�5P��p��ǆZj|؅]����!�W�5i��@�d)aPظ�l6Oc*0���Kf�0{E�M[Bg`X�/((9�̟�sfXM�ǵ(�h����Qg��j���D �	���j�5�K���1�oS�5$��s�D��24N~[��e�|*�rt|���}SD�}Z�=+@�}-�I�Jp<���à�ȥ�	�:�Q�:ђP���̂ùΠ���b�/( �d�:�1�v�&ȢF�� j�k�*<D����M��'dm ��!i������L����>`v��&�r���]8�|As�e�פ1?�dק��u�`���5�x���A迼Oל��*v��P�	�`g֨���U��,t/��������2��n�`�B�[��:2��>��:�YEr{�pa�%F0�
iM~x�p�]{D
C{m�p�6�-,�H�����j�g[<K�+7pF3Qoo�,F���|�������~ބ{N�~ȣZ�i��VK�ElH�Q��57&!&�<.��ExQ� ��Z�t�uQR��X��`�NBIů�fy����ґ�&\�P;�NZ9.u�|r�] ���N�P�Yu�P�K�]@Ʃ����I���!�~@"�R��P��S�=ħ�\���)�t�Z��@W0�6j�y*��o>�Q�b���=O}M���{#�K��d;�u�+(����Sf��D]7T�z"��-�����3[�k��O��k��sD�C�ÁEy',�י	���+נ�].�>|�,5�M�*��c�2�5oB׋f�.�=D�����|���E�Nz%���-���	�<a�wI�����L�}j�;�V�<�A'��|Om�7@m����2f�)�۶R"7f������>�>��Ԛ��h���
m{J�6�]Z���C���\r�r���^Md�K|ۥ։D��/�7 �V�ru�i�Ѳ4̖���G���T�}�-,�~K�T�w����i��~ۛ�6�#.��wa�B^�#��|I��> ���W�]۽�8�є_40g�ӂ�?)�e�6?#�YO�BYN�T=}V�C5�~9f NN���kU���ַ`CuT�; ��Β<	�;��� ���h�&3<N3�r�~��X6҇碷���`-��S��L�#3���Ws��\�[͈c&K�:i�+�̄B�<��C�ԡ�˱ԟ�
��s8���c�	8`~���b�@�m�lz���c���C)�%.P�`��k�<o��8�4��)�Y��;2����.8|�}Mv?Y��4G����|K���7*\;��c��V�H���9����Vs9Z�z䬸�}��$t��S�� ��O�D���-r�E3롖�K��U�b?�) ��E9$#F~3Dp�~��{s�_Q�)d�� ��5�z�=���ކ�$m�(b��fa0���O��ۊ��T둁"}3U�/L��]%3F&;�gZB��u�rڐ)�t��`�zV;�5�_����w��i]I]�f���O�2%�C� C
xv�5�{ֈ#L���*�Ӌ�=RK<�?��B��q�	<�R��MQ�9-���[� ���ay
 �����P=�u�u[03OR��uߧ[xw��0J&6���L:=�F�Y����E�F�m@4���	�Br���&L¸ �*F���^cݕ��R��qe�����W���c�_������;�!�דu��B`�q�q^ŀ�7>��u���B��U��E��6"T�`ua�ƺ<.2��A�.U�z�å���o<'������H-L�C���?��q͠�<<.Q�ȏ�Q,��ab3�*��.t����!�H�.��ǼL��;��rI��2d,�D�f+����F->EOs���O�0��SL�O���|ii B��!��竢/�A�O�y|mA��� �E3�z��C���Վ�$�!������A��"��3��zŃ��=���6y���q]�4�|�qD����S�[^�W%�L�~qg���,�Y�[H��J� �WU U�Ѩ	bz+S8��3K��;��C��jɁ�^G�
�F��b�������d ���j!a����M�����ԩ�/f���"���a����T�!������\��q���Z:�Û�.�^�s� (׺p�8ǰ����;�j�Y��ȃ8w��G��P�����Y�3`�v
��P�� �uB�Ju�NF0��T��;�6iS�H��&��8wV_��s:�b	���551��T�d�LmJSv������HF�^��誔���vC������,�W���R�4�
��C�77Ԝ��D{Rj���_��v]uN�����-��v7V>��Q���!���
yl�B���h���g�������P?"w@��)$��u��U�&b�byO��2/�a8�����DPN�L)QW��]��tS'�O�*����PhbY51�M�W,�ș��31?yX�9��ARd+R������]M��-���%ׅ�]v���dp��=<�g�?������m�߽�;�o"s�������;^a�� � :�3S���mp�<0�dc?�����*h�}H��L���^�'���ֆGң��`����Qҟ��Bp�����Q\�p2�f0u$J=j��r��<{��Y��w̛n��a�ZKX+-`�j��k+|�5(�:���03�.�O`o��2�n�DJ,QZ���<a8�r4��<L3�x�7�2&;�Z�Y��K�x�㍌���E��5*n�mWfRg8�lmahl?*�l�L+ƚc,;�����s16��*]q`�?����츞&ah^��>���x��C���?ڤҔ�QԵ��8јB�����z�!�r�k��q��yn,ULݡM�7F)�P�� ����d	�?N�Cz�o�'��c��~��I�����S�|$�G=���y�*�>A�1:��:�5���3F%��R������U��-���/o���;���� j�9�8�u����W�)���{K5M�EN+�«�r���;u�U�E'�B�0=��zb��\�^����qf9�I��2��¯�<���㽯b�?0��m�v1pEpr��8��ո8Ռ��lBsA�3�%qT8Clcs����-B��/�_�b�\�}��!ӝ��}���(��"0���,0'�H���|Z�����P@�3��0lk=g)6�W��u�������l,6<��]�S�5~9��يO���D��] �F�S��_Zm�j�~9-z�y�����U':�C5�(XV8>5cA-W�.���5��*��.���_�1�~xZ�aR�B�����%�4�9��T?1'y^B�	�rp�l!�4�@<��Zz��ź{�}P���h��4�s�����&`�5��r�Vrl6�ϝ�ϴ���!����;�����>8�2o���������A=ߖBo��]�.C��!j���$Z�9Qt�P7���.s2��"RKp�Mt���6c{�@@=�%VNw��4v��J��G�`���ʑ�U���^5�ud����R�Ǖ^����Num���a�W �G��|:
	TA�������Q���ty�����N��#pƺ 1,�яз�R�j��1�
o.��G>N�����[�hS�v�Za3|l0�.��2�|$s�ehF�Z��q��nh��ޜAM[��s�1o�����&oz�?�*��0����;r�)�����{����svx�V�+E���S_:u�`4҄���v@X�IzoQ��L�+����;���6YB�J#>����k8�?0��P��������D�w�Ć��ڵp�)}��J
eÇL���x����H^"��e��$t<eNń�TyN��=]�!�k���C\�#�fn�D�x�A��%��0�HSh��O[��fK
�9�J�o6����#@l���_�M�^@q� ���������5%*>؆p���x9iͬ�=,�8��R;�fa#��,<�4åޭo���"1�[
0G"Pn��@x�[�x�����d`�,�+Yr��"�y�V��e���cwS�a������C���H'����(R�$�gG�����	j���'�޴eQd4��a�Ym_�/�~������ii�!��+�1��@e���nz1��l.���54u��	�&���Þ��S�u�U�9�8Ȏ�1؏/�?zN���#�` ]h�)�±=$T�<�s$螻��u��6l+����AJ�ag�Y�܈/���s���7%nQ��*�$�,S���ذ�w��71��~.|���^�Bp���Yk�E���|�ǔ�AZ��tJ}F'���&[��͏@�2��=累��k�̘ݻǣ�mJ�}���~�"zG�4l���m����zt�5��V����FNe���8�յ@��?du�׾~q�"�bxM�._��M�\�~Z��b�חT)ζF�Ȁi?i�f�TJ��𨉙�-1Q߰Jcfd�ڷ<Vh���Cuw���J�?���Q7�32����_���	Gth�L�"OАA@�t���`�W�7`�l����M�U����+C����/�G�����Y[�*�k�e��-�J�9�/���h��@��w�"�|�myӭ"��������"��VA�3��Q`��^���Wh|o#��qPղ� �*��/}(H�ƽL-�B�����Y �ϰ���D�Z/=ӭ���HD�_wm�� ս�.�^X�Ʀ$9h�ؿ��$X�p���C Ed�]�\�}g5 [k�Wl�4˨���;�Ê���QĒ@�W�R]__�Dd�c�D��.�B�S��Z>r6�EM�����_���Ā�w9��
�Ç#5K~W�6�Җ"vw� aA.�_21�PF7s�#mݔs1�����xu��~z�V`!�FR�69�з �"~���+�DI�I=�Bՠ�>�I�7
�鑱�� �7�N���#�(��j����R��A�"$_��G9�~��*��a=U��NI�KcJl�8])p/7�>�:�"L�sU-�tO�$&�K��gRȇ\�0`�7RِvY�F��129�m����4����9��$��B�r�@�)�6�ko���4_��W�s��E�
s��NFV|n ��`�8^dtÜ_�/�l[A(�ݚ�x��,�=��M�_f��3B=�q��q��g؂��&v�$x�%�I7o��Ν�C���Z��2;|F|A����&O���V
�j+Ꭿ�f�'Y�Nx����Y�Du�)7m�\����[���X���@P��q�~u��5j���-��T-�z�	����Q���|~o5;2"�SZ���oN��>���c^ٙ:m/\
�dv7�z�?���N�0Kg����:�%�w�"�z��5ְ�Z��)��a�h%�>�A.�����&z����}�|�����_
���oɭ�Z�r�����n	52x&"�O�x~���`ѳi����3^kA�2���9�D��T0�#�����D�����$�2�F�|�L&u���ޤ�d��̭3}���i�7Z�x�4��壯DJ���V�U��J������=��^r�^/E�:ꪥ|�sEG*"���{]I�\���
��y���p]ƽ��M
�t.�����Mk��*�]�Ya�.kh*�&1x0���!6Lx�%]�W��9
����,��$_@̮����s���gÐw�Su����*�_cq�G*{,�UM�UT��P�12�-��A�\.�%���A-R�}s�.��R_F�1�ٳ�o�r����#��Q�/PK?V�-A�I�À�U���r1[aX*y�Ə�l���\�4���O����O[w�s�hqu�1�Q�t�ݡ�����XS"��p�=�������	��35��b�$�Eʍ%*���m���pq�I�Ӟ���Z����F��}�ĎP�d���)�K&B'�{$?K2�S��;_�w��瓡Ô\t�)=�pi#񵜆����al�<��72�\�)�["����\�����/��Ur�	x���!~���y�Db�)�\`22I�"���;�N�F�k=�04K�nm�����Cd�r�Gբ궽�A�bCe6����j���k!����j�T@|ub���KPa��8���kl�L�#2<>�Ƶ�*��:VM�"(��6�z!=�OS�NX��'�����s�3qPh1��oA�|^��v܋�K�(t�|ʽ�����E�h���͇��`mdR�Ӧ���{Ǉ�y:L���*��n��g�i'X�(-�(�̺w�1��[�kk�t�ܿ�+	�H� 7�����Ɗ����F��ls?�$Se�괼�6!�>!YqU���!�ȭ�&F�uJ�w�����'?�b�݄?�X������K�pAb�g:�����Ҁ��OјY]������'�NBn�m8��b�*F8��}�ę'����U�q�B���d�#���Oj��Hȕ��)�j͉p��"��_�96��tp$��s$?z��q?���q���z����]M�	�%��V�J�>:�fc���3%�uD�}*{�}r��pĂ�lh���f=�Gi�1`R����1�P��yoR�,�k4�n^<ߚ�t">�o��,�F2�8��f[d�8}B�zD��A2��j�k�7������>�́�7��n�����~,V�{��z�O�E���I��yR�u��dM�LRR�-6 ��������I4Ͱܕwf�Y��U0���+�;��Ju;���"���:ٛ�w^��
~����u:��K�-{PK���tt;d ꅮMo�+`i�Q�3����M1��Ƴ�H��,F�Nd�{'�� T� ����i3�{��'�@XS�d3�h�;7��ɰ�< :Э�o���Bb?��Ң�k}#�X°ϵ�,�����S��[�N�$���c;׬#��q4��/�>o�J�Gr�I��M����j��I�	I�?d�8��/��NؕK��]�T�{�D�
����p��iN�]�և� n��+r�27[tY�h�w�(l0��=�ޕ�� ���BT�*��s��B�J b^ƌ�J^rzz���A	+Ѿ��$1�gXn���EU��q�fF�r�kQ��(����+��Z{.l�7��bz���)�=:?B������L2#^`Qh��=�)�,6Yt��`��CnHA�����k�d
I.���(׶��Uc��K�� ʽ��=�w��dN�h��^t2��3Α5��qh���[ ?Oskdh{�ۇ!� 9�����Gq(l��~m�5{^�� �f"�҅J��<���0�F
�T�u�2ks���w��	R�ÓHӒ�s`F��:�l����D�����!�q�������4Ư�%�E�K@̈(��t��e���$�b#K�:�-N���]__��ԾrOP�;�m��A�r�m��~��;r> P�Hx+��U����$_��]|�-W{��&��ο�CH�,��5��{�	\y�.�Xun-�d%�
��tc�m�󬞥�2����R��h�61���8�/ђ�%3h���J2Q�8`DrX���v��ϒ8.����.�����Z]U?^=`��R�]*5���>�ӼE��z���	���S��f���v��B~h V��i0��O�����J{���bv�*+�3^�dx��_�,����˜G��r�t�ޚQr���㐺.��#��=�����SX��|�a>�,S��xCDDs�4y@�)�Pu�5ų|�_���ݷ~�p�`���h7D��ј�u��Ȉٛk{�p�v��P�M�R����\�����=D��������t6����!�	���Bo19�t��1�U��\@��1�U5BE�:~���h�\�Cc��\�Wzz�n��m[���'�L���id���Z�I6���������m���?��y��m��,�C��p<�����n!��m�t�@��pQ%���~�g�r��J*<��l��4Q��x]�WP]����F����襐PWM��D���AJИ�0��4�T��%�Ɏ�����B�
6�����"Bq^*�u�]2dK��r_S4;~\'*c��`�L�fh[�H�(�+���[z	��Դ���ŇV���@b�Ý�z8<_.�>Z�� S�WcGK˪�zn�O�)rt�/$��0u���	�-���~P�&>�iOW��p�D�.�BOP`�:�&��4�r=��5���q�>�#68=yWQ�7��C.H˲~S�F�U"ɪ�"�0���B(J��5�`���(��僧Kyc6B Rqg���Is1�M�H��d_$."h�u6���-5=<��� `��)����S�-���L���%��+Zx8$���v�g�� ���O����r�Sy[�B�4�јM	�
�.]�;�<Z�����zƟ,+�=~�t\�۩Ǖ�ܟ�1��I��������?^���|.E�X����E���Ņ��>���)�6�ibp�^|�k����k���;���(]~��� BL�"n�Dߵ2�T`��$�q�=�)�k�����	���G�<&�ֆC��ƘdSI�܊��*q���V�,�I`mo;x�8kK_�x���C���1ID�Y��ؼ�C����yF�V{�d�EZ%�lp�Ж}sN>��ڴ%�^m'��,��.���N�`������o��,�Zǻ��vC��*�VJ�ч�3@4��Y[/eI��z�inŌ����kA��aw�����N��}�S�L4�>��b�v���F�=�E��Yuzru�S��;n���:�����������VF��)�KL���ok��/�/��\t/p�a�������������CK��n��a�y"��L�p�����P�*X�7��)���X���YBi�)j�i����6���	j]W�C#���?BP�O�k��n�����8	�n��ЮSP�R�2�F���K�`�x*��� >�7�>�w�C晾�S�/�$#���{I�Q����_W'�8��hlu�W�_e;I�@��N&�{K�
��[��zH�z%EO^��%����Eӡ)��j�z�l��V�����T�:��j( �8�����&x����	P�-
�L�4a[Rޑ��$0�mǵ��\#�K`��]Xև��C��E�o[����Z�<7c����c��o�����ٜ���kNK�d���RyP�́1Bi��ւR�$
��Ǧ >���Օ����c.,��ؼ�j��SF�o�x�W�c����5�}�!�D������&�f �J#"��}Ի+a��}@q�x�E�'>��L(��h���ޣea��R��h�f��� �)*pMM'�����)�z�!��]�\��	���K�
h����!����߇ ����ڦ�y(�b�zOs]�ԡ�12�Y�_�Y5��������hGo�x���ok�N�*� ��`\�i�H��:c���%�^uGV�?����_kɯi�3��n��S���-w��f����}�_���P�f]��ʦ��?J��J���h�JB"Ȳ�<Y�!O&ɤ�<$��z�ƙ�� �!]��]���MX�e*K8��
{ �����a�.x�lyEqʒ��
�9A
s9��Ŀ��^T!�P��q72/�3H����!#e����{�&
�&����i���J/Te��(/�m�]a���ɇ��W�<û��wxC</�a�w��:��:S43+�8ߕ�B�^�3C-�ND�����9����o5E�w�w[q�3fd #�%l����0����6D��1�����xo���DO�=u��X�+��O�|EK�珁>>��ܗh���b�6��}�t���dj�%��vJ�*�i�zd)�o�WU��`�5���.KV�y+����p@�谴�x�����'c��"��jX��cE��v��䎒�x�+��t�X#t���|�n-�"0o�|Z��4���O��fU�㘎t�\f���=��H��\��K�F�+&�E�ⳋ4;�zZٖ��o�ULY�9�џB�Q'H|y�Z��	�%"��gTv���PR�x�_ntA��}�|���S�龟mV9=�����tw4��\�}.���m=e�<���o�Xt�|��;5ۡE�5�:�;�,ގ_2c=�{}�?������&\��:��j��.f��'��Q ���J3��F�B���}�����K���/�4�I�[���/�Oۅ~-y��Y��f�M����b�$ ��b��W�����y�Ҫ�^t�~U�v�ڲ��Ȑ��^�K�k�O7��6�ĕ�k]���؃��i�X:��?�E�a�}��+p���=��ƾ��2W���B��A�URg2� "T���\%N?���iф�`��ӋE�!��b֘�iȊz0F���'PS֚(*��ؐ��ƣ�4�D�f���+@��X�H�.@��F�9-O�@����X�G�xu�Z�4(U�_j�2��!���^`��]}�B&�U� ��.�C�7@��ߺ�N{����ՆyP2P��Vtn��!�2n��l�i�k=[���Jy}�U��U���9��XQ��|��Er9<=��w�8��YSS��y�EhG�����Ͼ�<���AQ���-��B�[������#�c�T)nW��H�;rHU	C`�l��E@Q�g� ���?nG*�A_�괆�hk�����)}��[8B^�3�ym����� �}�XiL��-�
�H�+^��`��j��8�j��f��<�v��s�Q�5�뚹Y��RF�����MvB��F�'��f��v�j��}�F6�M ��U3l�L�Ћ�q���OHJ�����t9U ��`&+��!3�/��d߾�_� ��C��0Eϣ^��\�дF��_񬦌�I��gZt��0}`�9�x��>Gc��`��UxY�r�	��ċ (}���t1��!���0�6�+}��Q|pd���` ӌ����i��5�.6�}-��*e�g)��0%���I1?n�iх�W�b���M��	������KOm�1A���٬���E}*�e|�U9���f ���c���/�v
FYK�R]���
�+��-	L�=�p.N1���r�.,�r��O%�g���!�U�� �+�hl"�q+L�K���wd"���T3b�a⇾7�T=4���ݒ��p��������k!�;��d��y|�Y丠�;��%��Oe4���*e��l��"\�H�&���~YZ���źk7`E��e|�B�r
@$b�l�f\�����8��q�(y��<��>�����k����L�{y���+ʞϖg��0�/�c�7��T���|�Q0H���]�n�#�e��#��Ȱy���S�,���:�Ɨi�6,iY�٧��(���K�ҟ�s�M�B��� � w��&��R����D�*c2g�?j�ȔG��ޮ-LB�w�,�p�OA��O
`��bz���ᱟ>�N�ഷ�]��}��sHx(��Fb�d��a�x�r���	�
Ț�mΑP��9;�Ґ�-��T�����a#z ��LKG���=읱��A����jޟ��@T�=�8�ԍ�`�^�ʹ��E>���"�R������L��#r�荙"6L��=���N	��ÜZ��d���a^� �^F�~��)>SU�Q��3��2Ǆa� �ZAe�^2���D��ė3��S�<�z�t�<�O�f�[)��QqCu�A��_��V�O{��|ܧ��k��~f�a�b�8	ֿD�=t��6����>?#�ʍ�^�;o�P�M"x:ux�ۤ@��D	Q@'�_iP�`�����1�U-fb��e;����K�8%�����t�U(��$8��&���2��ד![�xV���v-[��f�V��GR;��d��
���uZ@�Ge��U�:[X��C�1�帎9��xeo+�J����m�pNX������2
I�s��3�V�!)7i��k��ݍ$�z��g�Ψo%��:we���~Ia򛙄D0hG�3x�d@{6�섉h,-ٷ�`�8���ثk��}�
��)M &.3bq_�5f�P����(^>�e��רC�3@u���V�,D��s��_���A����$M�CJ���X0�����Q�ܜ>��:�ڈ��M��K�I�Vw^;�t��G;e����N#�X����-
=5�͚�sgm@�<?�9�\��1�'��Ֆ�]���>IvFX;���1�3�i"�5k�f�i�A~�N_��&i��_�P��T*&�J�.=�g�"M�R�'ʸ(���h���wvh��?5�2�mnhBv�M�֓q1
~����8��Ợ��uH���
�bm�=�L�t4+Kڵ�X�d^�P�4�>(\���ޱU�i@��A�x���b���˽&�8-�Zje��V>�GNO	oL]�����Ίټ5Jҫצ��$�rKP�j���G�Ѧ�6����P�ϤJ�*�
]F(*Sd�la���kMk��O��Eu��]��G�_ޢ�ɡԤ��83�F�擃�/����)e��s���}$�c<�Z���j��= ��ڢm��P_nf?��`}����A�������YW���� ���۠�m�C*��=1Ȭ��U�������h3��/����?�4d���kھ�FRG|����%?���b:�.{�"T�WP?�g0�fA�Ȅ�9wu��G��6sư�`3 ;�M�Э������Vu��9�hI�G~�:@S恂)��'o1�k�5v��a*ܼW+e�7�a�y�tuX�5#΂BۂOz��d�3> �ă��0;�4Κ5���Il?f* �	��d�(���ao},��}'�C�Ak���+�Ѣ�Ej�
.ޞ�p0g9 :t|1J�H����1J���|����3���Vqׅ����F�I86�7`�f-�L�Jyi��ZV��rkv��F/��Nf|k8�N:�uek���d����ڒT���{�Q�D���E�?O@�ebl���ϺF}�h� #�J6gNߴ��ҹ�a�(a��'����ӹW��~�G���U��I�S�!ЍX�B-��ȷLR��*J��b~am����jjBi��,+�X/�
A@��#��Z�ٰ8�rN�zr�Yn��C��=+���gn�!���6�?󆫳�D`?������	9�3�~(�-�R��wN�!VX��15b\�o�h�&c�&R���9�a��m��_~���t��	ڇ���ʭ�i�q,n(��b�:�����
F�!�au��>�1,q�*���}*%�k�@��2u$_^�Y��zzdI{P���}�S��� ��Qos6G1��c��v��|�Y滃��s	A�D�,\��\�#�PA�
'A��A���ۦp^�\��;j�g�{�Z���c��-Κ�N:AhFS{Ƃ��/���떅���~e��0l_�DCxt܌��1�X7L���2�0����u���K�"�t����r�'P0�q���Fg)�H�u��M�"�[}F~�k*���Z��R9�\��y�m B��^��T2��x\��V�����[3���J�z�ť��Y�hN�C){6L��)� ��)N��л:ː�hI?��p!&
�z���dQ��^��Qt>�Ȣ�mV�R*뮐A��[e��2�u�Q�`4|�UNC� ��RpK�O�z�8\GoSѯ�g����W�&q�i��hp���;ՇK��)X�T�U9�b�U}&�������O��$�ZxD���i�8��I�N�,pJ�d�*g���GC:�77!4+#�$�����|������~��iZ����4�$��/'�Xz������a@�R�k��^XQor�V�k0��
U�d��[����|���UY���+���cݘ���S��k����3�<j�[�yڒ�b�"I�+�@��7���2I�T�<)*��B��钓�o*�u5�C��(�dnصMx�D�ԋR%B�Qh�~=Jo]�E��O��m�KD5k/�k�M�;^��i!>�ӡT,��t��`m���/�M#l�����T���T����Y���K>��A�H:&΀��i�F���J�3.������Cb�ѷ�c�^���}\Э�*+�ty{B�#(��l����J9m#���pGg����Ѵ�
��/���#K:����z�a�a�c������Pؕc�ؤ/v�é�_)�݇-N����$�"Jł@���l����4��Z(5p$On�i���]��#:�@��%&�ɿvͼ�I��������x��O�s�`�P3<�cR�"�3T.2�rP�iƐoT��ܹ^z�f�C�m���^����\��tX�mȟ2��|x��a������9�͏Q�q�m��9�+���$�b\�ʜKvI�e��]�Q�}�/����X�����%��u���,����6�j�Gb_����S:%Ѩ������a���5gOș�
�#/�S� ]�k�\gՑS�KYq�^8�* eC҄%=�m2]���?NP�2f���/�-��&��f��;�������=f���Z�۬3x��p!�^T� �{�ר/��<ہw&Q�?y�)Ӹ��3A@�|TX���2���-ܦ�|�n�/<ȗe0�@^��ʥWh��/�R�3qЏ�k؀�ΰt-��^�NP`b⋁o�$ꙍ,��D&x_��<���<c�`��t���8��s�j��Py�N"J֎�^H�;/@W�?��ۗF��~�J��$��=�����4�U8rt`/d�:cK,��y�{��P���;�Y>�_�+�5��"D�R�i���pw�J�)'�7?���b���.Ph�p�:����n^����(��Y�pPُ16Τ�@z���wW�Z8����|Dn�&��]CU{ļ�axgii|��=��aY������X>r�V}W���V`��Z��`6�'�����aN[�P��a�i-�G<|��(Xg�:s�-����n$S��Ρmvr�&	'
��U};sZմ�ϾК�ru����6XO������:�:��hq{q~\pj�?����j��"��바#yh��6��T�sc���:��s��×��p��k+�<��h�����ڇV�g���EYI��u�����%&<��.NW�S�D��A9=���r32-]	o�N���|=14}�x�T	�k꿒"ze�X9(7�}���߉n�@5��A��d��Azl�\����1/a,�$�]��d�ˁ�s�l&G�ņ�G(qSc�9�X���-�8�mf���E��?���A�z����c��t�,N2�_��jSUD�\�PwV���P�'���/;�zx4�XP��ג6�"�IF�z��cm���(eO��"�%��a�?U=����ߚ[�e��E�r�E��!%��"��~���i�\@�6����[���F����Ɛ�����f��M���.�iz��F9"��P��Ⱥ.�����(���;�Y��l̕0^J�l��>mGen�UŨ�׊Ɲn��0Y P��S��J2n�X��	�	�j�D�;��Z-���>��CL� sh���B\ܹ�P�(�,�6ZK.;Zb�Ӛ�ߜap9��`q�Fp���k������L�m"1��8�E���#hF�ҭ��G��@E��PI�Pdw�Vh�Yұ��}>�*l���,A��w����1&'T� .�.�׺_�Ǘ&�1fr����-�1��%.���N?��[�zQ���ی�,����m�ZL>ƀ7�����p�J5�Ka/������b�F-�"�:m��U0a��Mg�pݷ��$b#ne&n��#��M]�ժS���l0/9���KV8b3�1�l�����?��W��T�KV�����b�r|����4��ݭRJ�n���'�iX5���4�K\ Ӑ�ݷ�%��B��mn��VB�ZԹ���a��B�D.�쓩� P��LP�->>��������6_5����v��r}h�! �M�;�0>�l��/vC��pf��TUybj� ۔lj�xA���СȥlGv�+�.�-[��Vw��w3�LP Y�9��;�B1Ͳ�A1�Q�i�����2<���Y}���g�LQ��ؒ���P�j�o� |R�ha�l�5�02l�� �!���(	������۷Kk��=����t�����?�ؖ�WtqN���ς��G�ŭ�qF���<L�w����	�
��󽙦L�7n*$ާ��L5� �(h����Q`��?44�sT� @���$�~m}� v�և�%xD n�=cz�!��C���WJ��s9�r�.s���e{Rs��f�5�h)�M|7?*e]eB���E��j��Qo���AP}�l_ĔCu���?���+"����w�����aE���7��-��~���&���C\�8��@�?J5�_��>_��F���S	5��`���X�YYg�D����y������Nr�������rtٸ��;�d�Tx�01��"A=(����(^C�y~���n�sL�
�h���J�YE��4����$V��zN[-��~�����r��+���������s�M�X���V�1:���vu[?�,j�t�:zn�!rj�lu5x�W��\9u��kZ'ab[���"�B�"�tNj�Hay�a���4��,��_�X"\o�� SM���5���4��p�b��I9��:WȅSҭ[��AW^�&����v�|��Ύ����|R���9F)�w��N��c���/�є@y/�_ +|�*ZD��X�{z���d*�y��P���"˂����U�ᅸ�8�n�.��Bedy��d$T��~r�6����@�Kk+�QȐ�J�u�hz.�?!N�s�$�X�|�,�OEW�m���26*��S�^�U�_L��!�����x�$B�8��ǔ�i�6OC�sY�YjY���D��)q+Ťc�t�Ӓ������l5�x]Z��n����j�)]fxX�A��ܗN����ݭ#K�`yuRTC)6n��<��{�9�� ݖrFP���P-�MpTA����(������cC�h�B.����:p̷z��3h�ni����z65�k�8~�'W]e�u���W���b%!�!.�N���C4Αq�c��pYFل��c�ߪ�w�ڌ$�r��iC�`h������;f��Ĺ\*e�!���{𠏡�Z5���X�\��~��|*{U@Z8�ڐ,��6�w^#Ϣ�^G(c]<M!LWoy3r��L�Ȧs�9���>"/f�I��-J�wZ�Ϭe	��q�B��=Sj��1 ��~���I�c" ��V�Y��V�b8\�@�7�_	Y�p�=H�8f)�VB�( ʢ5��b�û�N"�ݠX�e�06D��Rv�9���g.H>��(ջW�X���u]��t�]��R���ٶaY�V�6��j�_�d�g��U��PS��+�dl��� Ld�p��k�Y�k��\�q*|A�Ҹ��\x�"(�"���ڦ�\�b���2�Ӄ��m�͌���Y�G?���@W������/=���գ�_�+ڬ��a!��V'4B����m#ӏJؠ#�-��)l�tbb-�
���������n�AF4�~��y�K�d�B���P��8�/��B�dSQ�CH��cP`���x��f��/TqN[�t�K����M|�5��:�Z�Z]�����{�[���}��$����/r������Q��S�p���arP�05���&tuWv���m��V��5��s���!hGAd�5�L�@����?�*h��g3H��_I�$����o*�� Iκ���[�b�n���E�α|�G�t�G�M,$_b, ��Y������)L���ecR� �fn_�)���&V�>!N�}A^�_���<��Zo��nne}�gms����+�ܮd�^��_���AL�.�Dۥ�c.(��"��F�!�=��%"��J53�+"y��"�'�5,�����F������&!0�>��]�1<����.{oB����
�Ԓ��%�;,~�陾D�ǝ)���w�k��5����Kz(�5�D/Z���6���vWn�)����T%��	�ȇ�V�1n�*�/'Vz�$p�� ���~��W0ʓp PXMؕ����[�ݫ_ '޺���rs]�B�9�:ԭ2�Gب!��n����� ��]���,\��\q��Rӓ��2��ru����圇g^{
�:����C������7nP���^�|�ӍE�~+{�S�"=E%����Z}��?�Q��	������Fu]��e|6 D�sݏ�o�E[|��~�xmZL�
��ޑȷW��Q�3�мg;NH}�(Z�-�1EK�v ��9ǝ�\4�������>~	rLʿ\��.��Ԅ.s;j��z�%��o��8wP.�������f��k��W���dU���!�X��.R 'j��}��[�`����OΑH���	m��#S�RM���N�O(0�h�k���2�������;�C9������aN��餓[�]*��9[QN���^;W2��t���'�ʇ�Aֳdû11RM�P��/bj�r��gG��T�&M.�c�8}���Ђ��\`�xh0�xWN��jN/�d�?Y�`�!	ˎ��V^�a�5f��}`oV���^
!�A��v)��x���]�mp&f�+���!!5ӻ��k҉�,�>��~J�e��풖�6i�ݒ��j
�m�r]{�S������>��pӾ����hfP��ϛ��A�Λ}�L߃��J�`��I��íy�54����/��sA��ܘhY�9�^���e�	y)�v�¦x��ʙp7Fb�_�]˘� SY��J��>���ν<���Y�|��W��ŷ�U�+�鈲>�~�@���ճ��ŗ�cv�!��� >APґ�\9q��ղ�6\�D�ߧC=K�z��*)�V��L6�}����=���j�]���y$����t�?{;���^%���c���DU��釃%hF	�J�-8��e��\��R" ��|�(w�h"IL�ɱ��Ē��|n���4�W��\O<]ژgxb���G�M��U�IFfT`3+��ۇ1���!N~ #)Ս��^��U2�lD�cHO�b���V�%k�|���[ %Gs����=3F�ڞ�_o�\�_�9j����`j5�>���d�6����c�R����4�m(��U}2A��������W�܎W�MA|�'ű�g�����Mj/�)y��>��Z9ό;�j'�˴�GϹ���t'ڂII�$�t�Q�5�� @Є�?���)�������lhQ�At��E5z1��V�UA,�B��hŰ���"�T荪/�Q����IP��4�*���+�a��$��灯��k���>�`Ī�d`���WU���0Z `"�m7�]��jB����h+59&�l�U'�W�1�P#�'�<�P�Uw"߫�ԏ2��c������/��cPr팒��I���^��>�=x�I�^��3J��}���e��dK����R*`��8���tRe2��c���)�i�G�т/��';�b����X���0O���>�'٤�h��AǕ��^��*��[eI�z�l(A��ˏ��4���0V�J��*�Rv�/���wf��?����ZEWu���u�{-����{����X2��&N�[
]	6��ݢ�n�%��Z�Д����o�o.rfZI�qΐ�tl{�F�Ѵ�_\>�q��4���RzC�������*��|c�f��M���Ս*�+�,�i}P���H�cϥ���Z4����Ky؈x*�Ag"�\�ƶ�E�Am��,�\zh%�N�o���	�ݔ#��Ԇ�r���������pֽ���m}|���Xp����r�.n?`��B���XD.�e�^RڹU�z��'��MhR#U�Z���t�ABЋ���1'x5L$y��{D!U�hMro�j��$'��͆����溪ر�%Z�c�a���1\9��i��O��u�s�����B���q����~�%^�|�n�+�;�H�9��CRה�h���H��������B�eO����������o�3������I~{8a��;�s����sSկ���
��g��	�҃S�?�	�Ԋ�̓�9� c5ȠGwh������Ь�9}J���gSMy]TZ�s,M�| �HS��u�������1�T	�J_&�B��O0�&hJ�h��Wg\�����/����+r3U�rN+��ީٱ�=С������ݴ������<�D�\*x/��K>`_�(l$�Pd��Y�>,�\��iӠ�a��SC�����W~ؕІ���镈Z��E��[d�X�AUL���^#<�E�ɚ~Y���n�gRHg[r�u��|�b5F�X26Y�.]rg�����.�9[��%��oM���=w��};����|�$6�]�"�]bWx�W�iRef\y}���#�F���G�d�A�������P��DeͪC�k��o6?�U��uы�)	F������L^�3��x��к"�1�_/���XG�Y�ڋ�����UER��Q�=�^���iꛯ�E�S'rؽnz\[6�I�����k�!�S@��a�k����V|���b*�y�G�J���c��Iz ���e2���s��:�A��!N��*�U��13�B���/���p�R��1�5��J�X*��|{Q�zt�g�R��x���]�$h�;v��x����%ڳ]XW	��+���Z��.� �vH�kh��% � fz�X�ŀ�h�=�� ���m��:�`�N��˗W��D��	�4�J�9m�7�Ah^yq��MK <G��2���G=-K�5v�.�\�L`��� Z���T>1��X���*Vʨ�դ�%͔�j�{����.��˲S�z�k��af2��Tńl�Ɛ�T1!Z�a�a��ǛU��-��do��0��ԕ�y��!��L��>����ǈ���CPed�����M��@=j�m$�b11��R����,��H}�����C���`����8fv�g�OA��M���A/MM~"-�1?L�b���������L��}�V�tE�"Bm����f�����\�խ#^�6K�׀�h���c���N��|�eK2A���P�L��b"��/�]œ�57l�Ҕdm� �����n�����[5�|l��Cc;�9�bYz	��˧�$�ٵ6\ڇz�
���H[Z]�f-I{p�:6�H~��X�d����!_:��Ћ&�����ʞ�k%5ty�I���Ɖ步����C�� �	� �q���V<�Ay��{���y�_hU�NQ�c�ލ�q���:��� �i�z��'#�M�0W~�Q8�y�e�&�_1�9jC�M��ᰡ� !3���˕���f���_(�7T+�r'[����8��7DHB�ٛ2�M��qk�w�쫐@����
�Yi�,s�܆5���s����V5������xW̤�l��ˬ�iv����aIҗ��*'��Yrpv���űȾJ=N�Q�z�J�w��H��콅/�u���ũhN_�
�BX_���`�Ų�L�z���A!4e!�q|o��V�� ���@�)�$�y���X0��c��?%�)+/�cX�]�%?g����>0��4�F��D�n�;Wܶ�,� ����Gw�|ؙ^��փ8��,�����5tuF����n��#�����]�uuv~�S{H���k�<忏V2���^�D�s\o�&q�HYV�:�Pn��h=Ɇ���0�)ߴC+F)���R����\�M�&�Y�9�o'א3=K��82�o%=���IF�n�iD�	�ĸ�y9���DM�deh��;�.ahÖ�n�ms��/B��$y��*���n�rB��W��]d�D!-l*C������ӻ�6�H_�Gv��k:1�� �Ί+�g2�,���ƠG�m������ON���M7�﬒p���@��R*d�̺Ǹ�&0y��~�98�|>���D;�Mi�BL�������g�(���Tu��+i/eƈs#��_O�L����D�C�G�F�^8��&��R����B��e�(3�_�mf+��+�:��
h0L-5׻����n��0�vȫ�,h�
'�gܽe�4���xC3�9��TWS�K���)@e �S���TfTyL�~ȏ����d'o�1M�[/��p��?��8�!XL%�⠙��p�>��E��{�D�>��<� ȜJ�1��Ca1Ҥ�GD���M�+����;Q��E(���Q,o� �6�ym�������� e�j����{���&=�0k��AD�9>/NC)������	=~O;��[�"b(�L��Ǩ��щ(%���/�i9k�l
Ћ��.�r�2�~F�?�qH��8��	��l��^Q�MVv}�8Y+J��0%bL�A��`��m�淮���$���$�*r���V3"��4��׊�'_G@�i��W>,��6I(߫g��	F͐���ʭ���h}��?X/�չJ�q���n8%l���N����d��V�r�C'��ހu�ٚts�> �7|``٫��+��H���#�>2M���n>�]"&��S�Iz�<',��.k �L,�	�!����8�`u0�?��?Ŕy�pT�<��L20.BceN����W�rh����,��'�Q�'N�W��Ὑ��xT���n� ���й���G�yh�MJ[jސ�Q������;�dG�9�z5�7��3K�ץȥ����b��/�8�� Z���{1�g+�&��/gZ5�e��U����c+Ga���&5J��`��!������[��һ��]S����/_�kmx�/~����ߐ*q�sUuKa�B�	{B���/�(�IZ�?�����S�,��8}ߖ�?�$ki;*ɴ�T_pEӪ�����nt��������1Y2�o���e%�nz쵭��e�`p�J��]M�y�2�MQar����������X��G2���J�lș֠g,hk�H81	�nej��3]��Ƕ�*H֣ϝ�����q�������)c������oJ��;{�!���Bn'����Z�r��_��._�����3 �������gF��s���>����pհ�鋚�r��<��[\����Q�F�Z���L�Jb�lD��^�Q ��Y��h8n/
ԟ�ֆP���+G�!����<��]R,�]8�ij��Q���G⯀�����~{v��0� �Q{F�/ğ����,�݅����lR\�v�C��(@7J����]~�6B����n�r�1P�H�n�vh�o�}nޅfx��"�4��mW��惹���������kT�[1�{�A�O���"8�{�/����o
X�|'V\5��?��;��>�T4!�ݡ�g�B�6Jc��ɦ�xu���9��y�]��?7/!���\���zy�r�ys��gL��*98=S5�t'`�&G2�A
4p�a@k�G�a_�s4���4��V��=|~f�߉�3S���گG&Â�7��<t�U��ҩ��-1��w�;	#Jy���/3#(��y�.~�l�g�O|�zcZ�ԑL-�>ٯE\c�z��2C�z���4:�w�F��L�ܬ�}(NS����T�Z.9c�˨��+����J����fE�G7���3\%�F6%i.�#���)Z�K,Ĳ�&�&�B[2�d�P�Hِ\��Ʒ��n��2� u�Ĺ������	�k��ގ�mC��y}�Pj�w���up)KX��#-x�V��[��:�J��5(A�����=7�r�v���}�r#�-��6	@m��;!�JݟaѬ�J�n�:SJ��� l5� �,��f��Z_o�F�C:R�c�櫁�D��/�`#�8tM��P|8q����W�n8�"�I��5Dju|ܯ�ԵYu�i�E��L3�lGM��1��
� ]*fkj��d �g���l���;}J���d�ϧ@�\�f���R�+�x����T$�9�~�8��QXB�[���Y|�r��S��n~)�ͤ6�l�y���0�~���@�;�\���,OIjR����3gG���Ɂl�r�C�>� �r�>�`����Y1�'j+�Y��")��/��6F@X�(�{ਝ+�exx��!{�-���)�)�˛Zh"�&��VR�L�-r��0�Fx���⾇*њ�
#��u�, $�w}�Г-1 �r5f�J��ԇ!�^~�%�{,]*�Y#L���%?�}��q�a�Ro��i'J+ٯ���a-��l��H '�ecc�9ޙ���?�����h����Ebߟȧ�^x�X1jLV���}�u����������F��N>�6��W�k&��x�9�n�c�F�}��	R!�S�;h{|�Z��wu�#�
�4��]B��Qһg�a�.4c��d�`�<��.'�v�{j��+
�|�{M%�c�"1uE!�����o�� 9Q%t(K����!�s�0�`��q/8��yo��W�oZ�B�x���	�p����)�Py1�����JG2��w�vX�:��DK��'lb�y�������XZ����8�/���d��K1� �D|�$���ę�l^��y&� h��7����m���g
aF�����L��!Psc���d�R��s1jj����p���B�'��P{����d#��JoOaD�ҏ�|.�%��ZQ*�^��(jA�<%�1wM�s�{���M}�(�&*C�%�/w��C&yy�	^*�]�s"�2�%�R3��n��:��gn�HB�Cv�.��/@���% O�7I&�I������}$��Юg�ճg�@�t0�����K�����2������@
>r�z]9��$�Ĝ?E�@?��=Y2z��`)���׽��y���̜��#���-�؉��&#�a�_�Gh�-C]�<����l�f�`���j/3̘Iv��s�jP	�2�r*�V�/l�ݑ=�����l:���e�}Z��j3�XxiD~>ڬ|�'ZTX�����X�%�?�:��m�����"�+絛?�U�Ǒ���"Ru��}$�rXF�s)H�g����"��C��[�'_��m�����r�)�=����PH��L_x`#-k'n���
�ctK��8��/Zl����u"����ݒ`��T�%$��Ru#a���-�\@�w��|�Z��v^yXT.���ȾʒL���}4H��(0���B��9%*ń1�ʨ�g��l���?�	Vڙ[�'��:�u��Z��蹾X�F��Nq��A���L��L �d[��j�S�4=�tw�=����V>4'^~W� ����..K����Z"w���>� ��z@oa�� ��u���'E�%��8������Mf�x�λ,PT8��2'C�|��E�I���"5���eIO�  ����R����F-V���Y�2/Ы��^�D������6�:��x`����v��!<U;A1��H�{sk�+:@��W� �f���0��@������&�}����I�ͤd�Up-����#
�׎�8����\�V@~o�f0E%8EG�?ם׻�bN�<��=d~�3
��J�А���Z'�I��b�RNK\	Te�ʀu?�Y���� ˁ�� Kq\9C���Քt��i����h"W�̼?�ɕ��E������FH��Hr�q6%F�bua̱��d�n���̨hWB�}ĄGA/�%;��,����#i�zMd=�Fg[  jeEPtWM�t���j��~X��~���0�����|��+�z���3*�\+,|�Ѯc�p3��)(�ǘ��nc�90X�%���n*\�C�����Ac���}�jU�a��+T�q�
#qӚ��2���S:N�A���3x+ir&A��΂�gH~XךR#��k�Z�|S%���1}��B>*�ɩ���#a�9�h:����x;*�[�vDsu��^ ��jVS��6���ZҨ��L\<���c�D�N廚�K6)%�y�Q�i��3ʰd��(����Q�:]�@�}�@��Tx.x��2Y ,�e�Ur�&�j�����e }&�G����z����{����R]:��1�Wٜ�f� p��h訒��*�X�\����m.O�A��{gd_���PP���B[�Ǝp��j���:1���b��5�.�H�J.���//�d�cQ�0x7T�����d#�0�_������U�X��;N�"J:GqFm���#�]P�h$�#<��������y�!	�Q�|s������� tl��}G�:H2�\Z�q5�ES���F�#)-pTz(_�Ŗu�n�} ه�#�t�Tf�u��<�~j���4��_E��$�#��2��z�����07rV��_�G�<Ǻoػ�|��Ǧ����V��{�N���nR�/�_�]��U}-^�x�}ʤ��0�X�(�m����dm���j��3q���@1�� 8Q�*'��K��f(��펲$���X�s�1���
�{�j���t����K6xH<i���o��`����P�}ә���H�bHk�ֹ|p�r�a�|�'!���	�i��j�e�Ƀ�U3И��ka�P@��.�L��⇾�_2���a�����"\�����py��U&�P�y7�MÄ4Y+��I"}�V�3"�6zShY�+�r5�����R��S:c|+�����k�A���w��*��2��1�������L���s�W�Z(�t�c���3�P�:��f�J�:���Ѿ�8�����p /� ��ri�f�(�YO��3��`�kD�ŵ��?zd4�i������]면�
�m��4��;�"X��]��"����җ�G�Q���.�M*$O�
�� m4�"�vCiJ`�-D�
;��2S��l���K����8S�=�G�*9_v��.���BIE3��I|,�.C�v�XZhr���e5�+Yԭ!�=�k�?^���k��bM��3!��焧���VJ�����IZl��$j�k�~�#*ͥ��ס�#�S��P;I�aF`��Y'(r����<�$h��πz�-]ܓq�N�;^�<a)̦cǷ{9J�g�T�,�55eܿ\D_[m*�R�؃���!_N�&r=T������Qe��zj�K=*��+G�O����/DI{���u�j tr����:�⾱�D4�G"W�s����W5���$I=�4�l�SN��Z�5���+�=q�!�=��!-[��_�s��tdr�vT��t~���L�ZX��1��Als��ͼG�M��T�#/�bk�9l(~c�^)W�ߖg����1�u������7�S�>����X�V��$eFY�!!�b-�nef�OX�6T�G���Eqo$���� �{�B��$I�MF��=�k-`1Dx&��SX���@��oɱ��R�ȽVn�]F�#�πc�r8�HV��
��)�"��OA��n�`̌<q�G$�<�)Oz=���ţ	���B�T� �~��f޴E,������ک��f��YnS �r����]��i2�/��1�~ESY��l�@�E����}\f�{?���/��e��1��VN������ݎ�F�(?u����A�O���e��dc-M���+�.�cs���i�Ӛ��^}�v�]ʞ.�p�*+�Ol#�2b}H_ʘ>��|�@���{�q|hl�]�5;�[8u3b06|)L��:��Q6�z�x�]��,޲'�N���!�ZH'n_y��g����@F���{)8����z�����8L�#�C�D�&_1<s�D@u.�2�+9*<ˆ�Z���h���pbA]����bQ��C�x��J��tw	��%�ƾ��HӲC=w��v�1G�%+�ٸ��"�-��Z��G��s�� ������vU&b�2=8��8��Uŕ��\��B�S� �qp�l����9��-�y�[�d9�%"��C�X��r7����/Y=;V�J�QN�X-�$e��X/�V?���5�!/j�`.���:;���¼K�z�Jr��,����hs�FM���!��Vo,d,�>���i�ށ�1��W�*}��P�]՛8˭�9gf���i�"&�����_C��fSX�dJZ҂�=�E��ܟ�޽�Vo�0\y��#���"�5�i��'UZQ��к�X�
I)�z��C�����v��P#u|%E>?Ovo�!:U�u���!�>s�-]�	v6�������\K�]��^�p L._R*��o���aݠCe*h}��R-� �U�B��5�mA�r+o� ����lt�o�Օ13��r�R�Ăɏ���5�uVc����"�)�N��ϧ��u�r�]=��z��(`�����]����j�-XEu$\�])�wo�g����)h�Ű:�.�x4�l��S��A��"
��(�.��ĻK�^�j��/#��qL��O�C���� c�g3�^����j$�PcpS�쓝u��"wOl5��"5�e�,��L�^l��i71���<�A��]��D�|�Dg��\��Ϙ���l��� �3�s�js1�D X�=μ}��>���U<�˿��[��"���>~sr,eѻ���Ji���G�o< �I$�3'�5�(��~�@�d!*���>M`�҄}������@�<�蟅*�E�b ��%�� K�0�x@4u��C��:(��χ=n���C��y_D�,�yI�ڗ�4֎ 0� Z�����V����|�6��!\�[�������s����]#o��^��nĀ��1��2/.4��w�E�C�%�I��_���B�w���籝����oml*~�1/Zk4e(�תG�2.�xm;ѥ(s`�4�"�c�>oKM��C�\��23w���Yk������@aa��sn/����7��r��t�AM�H�%g#S ��31 3�B�_���v:�c��c)����z=����P�����a.v��z7�c��4�"_�&���'bo��e1��E�\#FZ������D2�(U�ߥ	��.m��O��f/4�]��>��v_�ׂ��D�^8Ϲs�6�=�^���1k	�K|���q%A�.���2�2�8���6��X��Fhw�E��d��-�2�.M�^}�K��a�ovN�� <C6��\�_��8�f�WY%~l{�C��=`I��{�_�1=5��q,��<\�.ݱ������9��5����u��Nrp�O!�p߄�\1�D]
$���J�+���k�4\V�Q�Twk�	ʖ�?�6m]l���Z$T�F�^W�5�069�*,?[��@�I2s���4�g�g	� ˸C����V��^l(�+f+�hl��pu����I�� ��{��Tќ�Ϻ��((%��8����Mb�z*=}=ub��,�{�4�9a���q�����u#�8�7v>&.�ݏ�����u�Ȑ�nϡ�æ�7d�~��	e�
�*Ҳzj�*�X�b<���������������۪S���d-�|x|M$1��A�Xg��;yK2rw�,y�Q�Fږ-�°1��F$c'�l	��
�(�%S�RJ��g����;�b���ɩ�o<F�=�,<��u��Ȟ!C7��c9	3Av�P۶6t,?N<~�
sl$z�v�1�PxΉ���������>��\�����hY8����[bL� �������B�n閕�hꁚ��(d13^�f�	��0I�oɊ<>%�j+��1�r���	GG�m�p�����:��%%�1��q3'V�c�n�.l��3q��p�k�ע'3��dr�	AlTm��"��#���E� >E����w�I�z��y/3��b?7a- x�����'ƷS�A[mT"[rYS�X�ׂ�j<���hG[k�
��޼k�ꈋ�+|�o�fͥo�ec#;,a�bm�`������J���=��q�B��(�=W%1
۩�%����ͻ\��GDD��Ӏ�ɹ��mm�եO�u ��D�}O8��eo���po
���!T���A*�H'�튻�H�P�ǂ?ny�oI�i����[�:[&�6���T9���UƼ�z�-��uXS���,[�՝r�+n���?��݁���̂
��r���� !L���ͧ���s�������h�i�d����<G���Q��Q��W�G�-��-
Tf�B�2�%��d$UO���@�8He�Iڲ85���&�t��ߔ�)gj ���y�LPP�^�q;4En���&���uYJ��g���(y�N�(aY��ɺR�c�!6��N.�����!Mh���Yp�Тwۈ4��Ĵ\����t(�@h�A-Ɠ�͑Ӓ��)�o:T��M��4J����Y�Ǆ=9ů�[Qi(W�B����vU\����F5�t�D�H�]��,���]�ˉdf�8�tҧMS��
Xb�����Q�QWKG��b�ԥ�����xP�g��d�Ɛ���ϊC牬@ú��p�I�T��HM>�
Փ��X
�������9�&��t,r%����;&����Υ�U��BAP����gQ���IĀWO
��}����|��9G������N����~]��� ��� :�g��� ��Jl��j�'�����j&W�2T�ύ(:��M�Q>X�P2����M|-����w&�����=p�pXp�Y�b�Hǵ�`lJ첫�B`nB���eq֯o���p]���ܰ����z��v+q�q:鱯7��#��(:P$Aߚ G�����o�Dw�*x��vMk�`T�d�i�iǋ��y[/C�m����S§a:�<�y ғ��6\�V��m溨䩊i��S,:{H;FP7��H@�<�U�z����>���]MF^�ͳ۲��\C�5�_�ڦ�c=TX.K��Q.��Y�6-;�<{�D�����o���%6�^V�=���u�u�+�]$q�.f�߶���G���6p-u8��b��V�0�t�IH��|G���R�:��\aYԙ��$'�࿊p��t-\L�{�Q]���P��w"~�_
� �����X~l�݈���m����B��,����bj�Z��E��ܠ;�F��.��|�
���EM�iP_�Ԃ��u�n�5e�JC�@h���d�K�c��~QR�)��'؜��{���T�Ġ�ʂj�H��
��b���6hK(+�w؊O2a����j�x�yJ�2�}��Gǲ<{�Y�����+u�yu]v:��~ZB1�=,^�W3Gf���u��������r4�-�&6�r�&D@���n��w�+�[*>���8�H󜁈�0�v��JހL�/E%P�:���ډ��W������S�5���gg�m�(}b%?�͠)��O�%g����a ��A0�5l��}h��>�J֐���>��{�7�Y���p��8J1����Č�9�P>)xp!Z�y��X�����O��aP0IK��������6ʤ�El{&���>���'B!w"x���BM�2Fp���G�x����ipPX�>y�m7�#�^��(���y�.b>)������/���*�vY��ؒ�F��2M����v�<�ב��r��p���nC��p���J�':�`Q���u�`���~��IPVe��RlU^���Zf���1a�4�l��$qA�_�G��}3�=���4^5�U'��~Ҡ������I�r�	���j�_�0��T4c�7϶>�k����mo�BV�\�{c�<x,���3A�Id��d��K�dU��li!�xcI���?0Wsr_#�{Gc�U���u�	�H ��5��NǄ�3��?հ�n�L��Íy� ���@K�[��2ؔ (�/��5�Z?�/���l/)�jRt��k����2��q�|Jp�9l\�e��F��n~�KT��Y�S�����'����3Y X�J���$��p����4���z�/�U�A��)R�-t"���C;�:q���'����T_�A4���|<� Z�:0�.��rw饋��'���M~k{��&�g�۸gA$�2DS�VU�����,��U��ֻ^�k�y�￮kh�5$*m�W�����lՃX��<�O����dN�Z�l	���R���W��v��uY�c�.h���x�������<6N�i!���.��~�߭A�Iݨ">�!�>�b�X_��Y�oz!��r�v��a���lR7���hT��������[؝6\x�?>��|}:���O�ڢ�q$V�Y2M���N�:�_��O�W�y~ݖ��gvkT�ɑ����K����R��o<1�G�|S4���c;l"M5��l�_R��sp��{;.����|>�vd�x?uA��#�29l���A�Ŀڙ��z<��:L���N�躕��8�PR�/�
��
�y����}�)I��s��=x����s�݁�E�\i��x'{�n�k?�D�3��<|Tp7"�C��M?���X�c ��'��(�g�]� �zI/��G ��/�=���;��dYJ��bq��{ݸc_���eg�ܜd}F�	�F�؁��A�ψ��ſ:׶�BJ�b��ӫD��p�eyx��g,E�I��}�c�e�M�fM�g~�h�B׼-�_lWz�Fp��m�΢��9���Qm�y���1�a�d�.��T-�~�0�!�e'�
���/cs�Ł�|"����� d$��9!��h�T�M���WY-���уX�����)��-�΍
؀�.ߢ�,�0�}yQaz*9ٰā'W;��U،���B;��k��V�M����d�fz�U�s��~~�5��/�N�����V_R��V>|�;DX��j�֕�x���gT�-�K�!�JZ�T�e��C^�6<۩�Oin�Rr��� ��q��;� �R���.�p��]0�����ﵓ�z����uk��_v�]h�|�E۩���׆^��oݪ{�q����%��f��R�[��x������v��K���R/���*1�Ƒ�^����_O^]M��3�Ȩ��Ovd�0��B����{��-⎙q�?�2 ���8�c�*3���~]�Q�x�=����_Ӛa�yY	��OH�ʼ��CZ"Vƥ��V�ˡ ����4�"�ӻ�K���f�\��ih�Yd8�yN������S��|��H*;v�!� 	_�=_�b����`�i�!m�Il��Kɛy�(l��5�թ1����q����c�_Kd7��[���3p0�Z�\ SoE�`�N�K�S��`$A�u��I���箾c��\S�?�Q����j����?2�A��c��S�O��[>\�.��i�	?KW�ƙ����p2���m�����E��n\�0?����4�d��2�E���	�2ߗ*��fS����')��gѪ�&��H2���`�2��c�
mȵq<M�������aa�qRx���]~�h�6]��f2 c��*	��B~�}��恳���_���(�e�?��H'_麈�qj<�t6����.���1Vd�ʣ��0Q�3��s4����g�/�H�W	�KM���suT��b.o�{�0=w7��oSQoЄ�_���C��{ ��杞D��>���t��. W�'A����l���U��Rn?2c�"6�o�hV�^���j9χ�i���c�x�?f�xt
h8����L���IZ�	�A�`Թu��eь�� @]n�\�U*HǺ�D��.R��o"�����b��GR�
 f��`�s9���gJ�5+�.R�#����2ٚvh��+"k�$ua��c(�@{�]��9��I������j�'�:�3�j��PU`��ÀP�&�u����{F �m�-��j�׍�V#�'"T��5�E�Bd
���ܥ<�x�C���&)�{s����3홐�^S"��>h��dA�fk͛���$�ȁ$P���g�j��]8��v�A��6ո?�(NGr�?���E[�S׸�s����Q����
������!M{�M3�Ҥ�H��l@��?����٭<34Zv�Z�f�x�_��S��q^͖M�#%��{*ha��C��]��I���=�,0&b��'C:t	�K;H#扼x�j�:���Ӹ�i��Y��P� 4�S�A
�W��=�[�}�����_�x�<v>�g .������I�s~��������XHN�nGz.N�3\v��v�j�0*�D>[4]�$�l���v�8�&MI�\��&���ȭ�,����r�h\�2���љ&u�B>F-}_� ]�C��+�E@�ѳ襡��#*�ж����Wo���8�Ӹ��]��j4ӍOga�v-Tifw��T
Hȿ0�"7&�),�䍁���H�Ե�;Yᆡe��뼠�u��L��"9W�t[��e���$ƫǚ+ƞM�����i�/8*r���O��t��R����AL��W���T��b�\�2+��1�n6������QFXpU��D`{�Z�>��`�;��,9���JV�'�K�G�Lt},��}�E����(Y�7���l�`�z1ò'�����tl&���iYy9DyUP�[�K��_?�V�����#�<!�D�>P�ٙi��hv�jLv`@$.�� Z�k�X<����"��?�V�O���r���U%�/�j\\��[a�)N޴����*��J^7�n����Iw�<e��wr"�|Pŗ�o�l�~��R��6�Q�Zg�I�4���\��
����^�gF�<��ȵ�ah��"�V;�.��E�)$������"3����?l�SH�����j�ڦ%z�$r��ߓ�<a�p~�pk�UNM��au6o�7��2��D��F�Ef�P�D�-��<q��X�$Z�.�.PƧ�[��t�+)u��c]�G�@yU4�	YD�Z�'n��&s�݅��75q ���/�Gߒ	`mݱ�n�O͝�s�K�)��&����Xw,��}a��Z<6g��R�&7��~���/M��%,��5��g�Z��7�R��P�+o����P�_�e��J���	m��.5�����;���,FJ�a�`�l~��1Z��;-w2��$�E���{nkc%%Z���b�6�ݔ@ok��O�R<�H%2�͋��UN�\X�݀��V����\p�??Nc�9C�����8��5V� $�/�8֚��k�4��n��Y�&��p�Gi�Ya��b�����f�5=q���5-��<�&�4��
Vev�~��K)\�*b��ʍ�	鬅ڦ>�{.�|�@��ST$u�i�����ǯ��G���[,v��:�m�����݅��]�_<L��x��u*��ߓ�*�/�j֍�����Myȣ���.�K����k�4�u�E �D�������'�`'A2q���F�����c3���F�z�0�<�X���v��lxP�|�^� ��0�SY�:�w���9:���,7r�ny���d�v��ʡ��be(=ǋ�`�}�nקF�X����]��ȱ�bk~ae��KF�4��P
��^�|/�#�o�u��e��z�x����c|��54���Q���2(=�,䶼��	2���QI9�2@�u�1.�	�ǋ� ��{4Rн�$E���.��M����mU}���G����Q= ��H�IИ2��Ѓ�4G=�B�׳��1��J�>�ŷ�x�Zz/l)�9K��������G�}����`f����N,��W}�S8��K�{�-O��>ؼT�.��W[%�e��O�c�E�����5�v���{f5���j��p0�]�	{��>i/��R
0��ږVS�Ѯ�D��"j�B��FJ���6���%�<��g�Ѵ/�7�@�è�C��K��<�{�23�A�j�W�	Mi�I�5aF���'V�jЈt����*l�q�<n�>��5uJ���S��G�nNԑM��T��A���!BX0��>l�P|���g�6��<yV8D�ۀ���v��"�Ξs�Z�/�{�X�J_�� `F�e�+�j���v�'v�C�S�g���(Z�AN�<���ק|��Y�8`��n�S�N�09ɗ��x/�4�vd�.*���Bű���MK�L���7/`n����meT�v�?D�N���C�)�Kc��!���O��*x��Iy�3߃��-�o�`�tO��Kt�>�$�����L�`[���2���&)[O�+��qϳ�w7^˺^�ٓ��L-ڊ����{��P%�"r���T�9<�-���kyx�S�}�6�c]z2IXZͿDZ�Ņ���&NN��qr�b)������T�so��E"
:ۉP�|y�$�Y�f%UѝL��;Ha E��\ �(P��t)$�|ŃX�P�:fS�^����U�*����1fU��w�=���?BuW�].�A�y�+�� �\��61�����������R�������N}x��� 
Ԥ��\��	̫[�uN^�K�XWFɐ]�Օ��ʧ�Q�I=E��ε9 4/��������`�S����h"����5�φ/̦3�X�gb�yr������a`��:��ODq6�'�U, � '�Xz/�mÚ��ى���)&�򁴴Y��h-����A�/s�[�#J\��fn^�m�CF��3���Uj'�7bd��/ԄD�p�$�(�Ȕ:�X�/��F�@�6U�q�,�,yRn�`mM۱�Hs$$V������֮q/e#��+�
��"��0��9�ڡo_�� ��o�sR�49G]��U�S���X��dK�k��7*�a���_8�sX����"]h�8�Q�&�+.#l;��=B���k�&�T�{n-T��,7��d'[���:�$�P	#�p�y��M��%ʍ<F�j)��/�N� ,Ǘbs�~_E����XR$�
��.9Ll:��g�;��n��W2	f�f>�cD6垚�ސI_gv ���σ����\��4l�!�Ba�4�ߏ���vy�{�^6-���z�/�;�!!ÿgY0Wp����o�d��e���Kj���6*�P��$��#wwh��ӡ~�xU^�B�r���b�H���F��%V`)�j���a��bN?ؾ�B����3~ωt���i�2,��U)
A/���(�S��㜛NwO~�[��ϓ%* ׋�n�� &�Ww�c6toz����p���bйP��03Ζ�غ���"~�,o3>\}�߾Ѥ ��ݖ��&�_���e$gc��lb����h1�l��\��Q���r����a4�E�8�ӵ�S&�>D��8��;��o/H�1�����<Ń��q��5��K��o1�k\k����!"�)�1�f��^���rŇd���R�o��[x�#��Am���?�ј�C}��k<���>݋���&�C��7"l����9�FCW�w�v�
M��]ꜙ�;*�l����7`Y�Z�	��OJ)���z��ˡO_�)>��������I�ɪ��+1nb��mU��A��s-՝��<Wb���� �`��<8�RM|%*|ԡ�w�2]�T�EF�N�&�i���@���0땆��y @�*�f�������)"��}RX�4@Q]n�9��ǌ'D���i��ۢ�(�������{�1�w��+F�-Jd�K�6�f������H�nOJ1Mr3)fYn�Y�*�z�/����?70�l]��.���NI��@�@^8��/N+��?�C>ALSUN��G+g�e.>���'��D^�_���Fp7L��Nĭ��i���l���<�z�^B�`T%��tr����Ή]��ÿ��`2�Y$��V�A�����a�te~ĭ��|-|��7-焜� e�1
�H��bc���Ѧ�N�Y�^DS��S@E��~�:0^����w�W�,� }�,�E/ۼM����ϒ��1�ʰiZ�i���J��W��8���W�@B�PJ�q�gY�����b���������yN$S�N�W"�G���	}TTy��'8C�#�ap�$wS���ߨ��J���F	��� tg#�^�zx��HI�C����5���쭸���t��M�~ϓM&V[���;ah�܎�|���d��m�뗈��e�I������7"��2���MG��/Y=,P�5���;�8���aHM�equ�|02|�&���Ғ^�c5py�qU��v~�����.)q&��RdؑIK�u���� �|̯I�"7����@��؉�Ǘߎ��[DY�;N�ϏT��3��$��@��BӭR�����e��`"��**vJ�v��r
wh1�.��x��"�D+��~�6j�n��N��H-��k?�ӆ���}VϦ�"C��,���&eN�ckB����#��2R�=E�dȧ�e�?����S\��m��).\�qh��1\7�3��,�B2�t�������i��Bæ�oi}{�'P��
�~ko�z\�>�
��"�$�h	)��s���=;�zUi%t���~�jR��oIإ8x�O�`�lb�R���O�RD] �_�Xu������ ��MO��-�TGɶ��١�C��6��12�?U�oZk	�0��~��`����[x�gPU1���	_��4�J�m^?*�
% /�z��I�K7�����\7��Z��Q?�C�W���nhhW44w��G�9:q�Zَ�.sR���f��2��Y�2	��sX��L.�X��Ղ28\�x��3b��	Z�E�H�&FZ���l �*7X\��֖
���- W~΍K�h�)��)S��Ő��棸,�VYwYMGab@��9��,q#ˤr�cek0#`����bLP׍�Ļ�o|����hh2+6rT߉V�m���!l�� ���y��U~�������]Q=?~��tU���//h�D".5�Wq�6la��������(~[�	���aW�5���z��k�"�_�D����R2؅f`�m2E�A��5\os���Y5Һ��}��^��U�J�W���s|j!J�j"o�����JXqI^�"h���/��y�k��c�}j��a҈O�����9>��L@�C?(8t'��Lsi͇ӄ0](�Lsk�[��E�����e8[i��ʍ��p���(�]��@�W��+�8���͔]��F/`r��@G"��F����(��u]a�[��/������9%WOUV@Yo�7K	��f���Yp��+��$�_�`&U�ɆM������t@OuZU�
���K�7yh���*�ۣrN�Хl��^�B�m^p|s�-�� ީ��>'���Y *`g�A�����ZU�L���"�^�W��r�v�=��͕֮�p[pqT6��>/)N>�n
)��pWY��Qm���@��ބ��1��q���C���ˍ������M��O���"s� ���}���'�!BmF�V^9(y'��h�9a<�'FD�+g�-�s��n�a:5�>)���@J��28Kv�u�F�����* $������0��~[��͠,��|�B����k�����їT�aP}���P*I�Rq���~X��Sk�A�A8�5%<Y�q03�H�)��z�TǙ[�D1�W9x5��Sc�h��z&�������:�<*���(�B,TC�k���G�Υ��!]���	-��$�}D�K�mq���Z@�&ړ�N*g7��͍�c�(�f?l�t����xvޅ��`�+�L�u��RW��F���-�VКm����vFK�\�	M��s���1��
V�in)<�nBKhƬ/�qJ�-�oEMC~Y�馨�ٗX�-���-����_L�J���H�ݮ����"?J������1���t�����R�φժ���߈� �n��}�}�� \�gP	œg2�p]^�#N���� �C!"8$�ό��%â��K�ԯ���{���tOÙ����R�}�@3=��4��t�����X�d�rĬ_�E��fu�qU�Q4���,�7�F�#�?VE�$�*�切1.�=�n�/q�p��63clh�?�z{k��D�$�1'��vd��);���r��Y���pH~�<ib�'��W,�c.@�%^��4x�ZFg|_GV�� �qU�d��
ض���{`�#kh~KC	ll2&�����OS[�\)E��T:r�����G\[�~VUm<լ�� �<{HvV� �/�A,��gηIUn��x��g���qj��� fT8-&�sIm.T�	��7K>|�2���n���E>�(N=�1�$G���l=���T'P��c��W���S�m�G�U�2�rr��9Gu�j��ݐ* �[,�91��ˡ����G�g�x�j��Cy��7k�县H�jz<�
�7�,K����]\hA� '�3�'W��!�`Q��h"�?�����	�!˻���{�#L��mY�C��4�Ǟ,:E؀ ��àbq��<��Ӧ�輓�g���ie*+�m4�����u���|�����m|B=������-���e��N��q�o΅2S(]��E��j�Mq�Y�9
(���os�6�)�g�߉O�i#��`|1`�[�y!���RsQ���f�V���Z��,����@t���N�s�s.9�k`��S��L�L�PЏ����T�$I[� �n���Pa�����Sf_�*ۦ���.�k�b��h&5�V)�"O�>����� ��>��9ў��7�6��5A��B;����(�2R�Hr�bF@���z�REs� ��(xDU��I.9��it~����,c��[�;�G����m���h��� ���K`�q�5^��7��T�݃�
�4�29*g��}�V,+�B���Z�gʛ���;\��!�u���e�4�2�N�6y�	�	���t�
6
s�-�Z-�f@���LM����{D�ϋ�P=��ƺ���>C1����������(��(��w��ķ�Ck���a@Z��D���L��䠆0Ƴ��L�J|a���{�c.PN�(Dv�z��n2�)��V�"���H� ]�k_Ğ�`ٰ-Q0T��p�۬C�<�`j��1�Z���G�]�4���)����5�Tin>�!?A�˶yy�������>�ˡ��V�H���ko��.=ף���G-'r]ޕ�}-�*v5BS)��*���&л\�?����7GDm��SQ��W"E]��о�7�`ƣO��ya�zH��=r�U{l`aB%WK�'ح@H��N��qk��x��m�����	�͸hB��\FN�xr������0'��t+_����
D� ��]�zTZ񩍠�&*'��ș_�����w��i�"U��ozA�V"�f���BM|<��_�6����X�Q��uBff��Pe󢠄��9E�XN$�����[UO�ҽ�:�AUb	�xQ��~M�-yL��>� n����LP�@O��f����Қ�/������5>�n(�9W%j��gH�>pV���:�4�<�Y����C�|�[��E��ƽXrbƽK.���%Ǆ�%������ �`�(�BF�ꉹ���0�q���Y��ߥ]��C]�}�R�j�tr}zL%o��)��<��Cޥwt��#^*��l�e�Y�����/$�JO¿��?���Xb�W>�E�����:��S���ȼ�SXbQ���N�[Fk�ۺ�k��-0�@S4��&]'qzq�X%*9�dSm��縯���i���zuX��۽��L����Na|6�9�g�p��4̀Mx/�;(P�Гf�Hޓ ��E� �"Ӷa�2���+�W�q�ǡr�{��2���t<Vhs� �F��A���w�9�=z�#�q�z� _��D�96 ��f��Z@�kߠ��G��b{��W5�uP��x�K�� �y#���=��`7��A3�<U=��^Fxc��m\󳙺A����!t�M`���� �+DeyU�� ҫ�J���b��q΀�t�m���R�(�^�݄U"3!��5G��j.O����[+)n(u<v��&�+�x�0�@��u2|��Tj/�^�����(�/�O�F����C�c�4EHS����w�$@/��ȿ�J�H�	�SŶ��WF.h���$�L�0�0 � �sk/ÔL��8`����]��c�GĽ�e��GV�������3m۟^M�j��!�]QP
_Bg.���kV�-0LK�]���T�V/�6��L:ǔ�o㨋+�E�i�SSĘ��P1N��ƥb�����D.���Q�d}�p:*��^����P�1�A5�j�?W�@��W�)�@���.e�#�ȘnIM��ϐ޾Ĉ�ou�Yk�XbQ��hH�����[� ��ٍo��90xn���0��X��_E�}�De�]�K��rn|���d	��.����.�Э؂H��e$�����#��B t Ι,��^�p�i�4"W>$�Y71dy�v���\�-{'��Pj�WC��S�ݛu�¬v�院�����Sv��qK{b�S4Uw��?�@�e����]¾��;��+~�.C�}�)\��h�����0��\s|�J��$���NtOxQ����������F!t8w���!�q �`8�_*&#耞��6}�6%����cQ��q�h�oD�D�B�FO�%�w�8��a�ßZ���*Z�	��d�1G�_dzTD�|��� �ƫh���w��{YL�ݲ�-]5�D�Gŭ���}ыR1O(Fm��M�a1��+�.�A�BzPs��TF�N7H┑�4���.4��x�:b)�Ta�|G�ʄ�M�l�L�4�w��@ەp���MЌ�n�ɗGS���i|���A�����!׀*��"��9�RT�R�&l�;������� Y�E	�w�{�W�}�r y�[�H�_��A��҃	�3�nV6�]]T���v'�3�Ɉ�n�e�	mZ/Ҝk�U�`Hׅ[�fh\�������������V�?����%��	jB`�i�a̿���1a��c�I���G�qwPTT�n���S4Y'uK08Y82���4�(�01��~L"����R����O�U�7W���Jf
���a1#��^V�z���ZRǦ�&"�cq��I����(��Fއ���~V����F+p�Ic;����xyG��'r��&���˓ƽsMʿ���)��8����=O�t�ƬFw���Vӽ�%H���*�]zj��,n�v�O�o�M4r����~�����Ľ�Z�z?�^��2�8_�΁ǵ �"�H�]ͼ�J�� ��R?�g�e~w��hq:PeW\sy�P�i�(P�A�,P�����4�.�0���/�i+��@�}.��f�~��';��b�S�Q�2�ؿ-��!6���`�|���ؚ�09q���V�rb'c
5�@��Z��ɪp=�S��zc�&W�UK:��H�km��cðiF��\�W��]��r��$A+"22���w�X�.�- �y𿀭����%o�H^�{kJ8�W�g������:%���dK���P��O`�7�������b�3ۤi_FopDO,Z��j(�k\�H���ǵ�#`E�l�z`�h��Kv�6Xݥ� lz�2r���t�!�Z6�s-�܇)p�ē�W��/ Mp����3��e�mi50���Ѐ�/҆��ZiE�]ͮ$�u�'���s6Cw3M ��8F}�U<qv��{]Ӹ6��F0���Y^Q�!���E� �u�;q�`jB�&ȉJN��oǗ�qZ���8R���u���%1!��FxI[x.6h�s�&	7��x�|��u���r����(�HH�u�L��G$`�o��,���d^�Z�v���8b�Ro�􉜍�S��r�Ү��t��j.E@�t�Sw�Gf��n�\�u)���ė#��M��G��d;X����m:����8�D��Հ��Y�6�$��e{>�3�
Y
�|G�0U9�Q03��[Zя��e��ŀ��@�����D�,//£�:�>��Q� ����2R=D�h�����Fqg���V~U�]�Y����*o�����f�ۃ����F�k�:`�����r�k�_������d2Z%oo�3{Td�fX��>�͕�z�|3�wE�m
�r~`_��{+���DY���R�w�ެ��ȩʷ�/�ay��_R8Q\�J�l�%�E�[� �u�-W�AE�;�t���,����AN]��?V4m�4�����j�� Z 19��ݔY	l���:�-���y���ûR\�����M�=Y0j�s������E��X����}��˜^���Y��l�W�$ĥ���r�`B����8<4j�O�%EETxe�m���F��,�W�+�ۏa��u���槇���89�zu�Nei�&U�p���|9�!䶐��>T��u{��f7�����p�<)Ω���q�ï_<�Zp��Q_��҄�P������J�����'_�h%��
�-�1*���6�g*]B��	A�8�ʂ ,�r[#�PjA��:IGcf��H�ҝ߶/S�U��eu��t����(���o�}�MRL���{� U!�<�Ђe��o�H�3�#LL���4�A�Y{��yZ	�!�l��,��+��)Gl���n���Im�GvB�@��k��K^�$��d���g.Z�*����m�b�3U�_d��2���iM]��0��{Q��_�����ȷ�� K�"���o��{�7�v�q�A0c��g���~S ����N�u˜�F����:�-�Fn��?��e���D���H�w@�j��gqӡ�]m����a���}<���0�~�w�JF:`I����xo]ߗ���P�S�,���2��>�Xn 9/�R�m�b�F6��]Ô�
����'�0�����r����� �.�%�$����N�:y�Pv�/Q�����-Y��S�S�j��?qC��hj�$ ���bmu��w�dY�f��>oFx"�P�gK���8���	l�j�x�U�[C�]B4 y���W�M���b� �����""�c�~�͓_;�O _�A:c��G�u"���f��ͥ�́U�#I=9�vo���r��݊��י.����j��Հ�m���1��M+��7�B,WS�h����m���&{�9A9m��%����7���8U��2fǿ���~��]���SZT�AE��d��R0B�����$y�ud����쑶�U�߰z���C@]�nD|�o�Q��,�v9��oL���.�RcG�ƞ� �>��˖ ��4�A�W��;�K	Z�
�[6l���b��b��sQpS/u�5�P4�G{A�-����a�a=���0Ƶ�g��o��9nP�d�tzm���U?KU���:��T�\^��u�<��[�>�7Eď}7* j�HwH$��I\��r[��{��Y���	��ݼ�VDΝ���7����<��'�}�����(�A�̺盼ˇ��m7�I��$��b��s�R�}3�;�qJ,-��d�C�7A�bk(�"�� �s9�!�K���e7�7�i����3����b^��}L`�s;�t�� �z5���"IM�ҋ.Iͨ2 ��/}8wW��U�&�ku�d`!���F7[pO�{�s�u�hCvV4l���@�a�Lcĕ���K�ًr|⡢�*wfQ���4�@,=c��c\�����D;[�&�D@f^��	4#m�0��W���u#8��q�����(.�gK?��m��n�Ȫ)瘖���K�j��E�-��k',���1B�����z@Fb�ĥ�ҶYb2D�l�ޫ~�G�� �s�����Z�0���+�|���'�jv�R5��p�-��:���uF�b�����Y��F����_v�Xy��#'L���!gO�D�J�E���~bF�8��}w����3"C�W�Pc��8�'���HŊ*O����e�2F�\f�:�v̹
-ɩ`�Q�  >�"���㊐s��/2�e��u����])�6�>�|�v'aI(F�Hk3�]h�C�X��61�~��#�&<��z��"���b����n.bB��+�C��p8q9�"��֝?�+�"{�`��u-v�7G/�R̉��-�$dlIPu3~�Y�%#��zC=�N��\"��b�9 �{�f�F���q��j�j+�/3��\�o4XG5?��*�\��p,<�ɾ	d�)X�|=���7c�W,se�mX�~�^�1!�m!RHg��L�'(����d�wcH��n�ɫ�R#N�����:_�	5�R%�Q]�����QO<W�����;���} s��Y�s��ތ��&5mL:��)�P����[m�J���A
�N�L�����&�����ۺ�o���MN���vaT?�;��L`h���^Gp�ٴ:L	�E1װ�t�wt�����rO|���$��V�f<��g�(oZW�	I)�P[z�u��F�byD��K�!�1��j���S�)�~ܤ�)�=z�����O@���A=Z���2�&�I-��=f]�����$��D���%R�i�Ǭ7rӊq~U��fNm�C�\
^�{o;�Е�	I�\���J,[���q�������c�Ί˵�g�ַ����\#�.�P�~���^nȌ�޷��_�~��v��f��2v��u3��&�\���H�.�(x�yo� �E�0v1��k�+��x'� �@ڂ�ݬ��mTpoY�����_Y�7�\�2R�]���^а�꧹��A�ܞ\j��9D�ۊ<���W��O���
>�AѰ�p����e�L��x�-3��K4��lTI���Ϥ�q�C���̉���5��p�!V
�t�6[K���5$�B��FGB��NT;�;����Q�lNU����;l���5�B5��S�dj�3"�cG�W���Otr�Lb�3�'�hp�c<��L�&���5��M�^�Ŭ��� ��+���n:~�����_�
���!�U��(�7��fM��q���+�xm5$I���6�?�ݥ�(����6���Ug��x��1/r���C=^��(���ϝ >͌���3@����BU9�s;�g���_w"VT��;�q�q��ҳ�I3T�{D��a�6��"gs�v��6?�BT�\���>��@ٌ��y\�8����<��3R�"�!7tu�V���~���O����ͯ���-/;��mN��W���.���:N�-L�[�5S�
��M��$����T7I�g�]0�Z��qm��MF
�‬����Jzܡ��ԇ*�lx���T����cT��\����t�jp�f�s�.��m���ٲ��`�u�`�{�x/U���{�����9���_:�!mZx�ը�;��V����g`��T�T2�r�V�(x%��-�0�7-��+��u8��Yq
K�*=!*Y�y��!��r��_���r�N�4?7]D�����^�K-�$M��
fb�"Ps��?&t�%`��0be���۷N�hrpԾ�(Z�N�P���{6M�}���}����gk&0�̥2�֞�9���"ͅb�͇���Z�?*� �GVY�A�.7�*Dr�C�����I�ÒR/����`�;m� d�(�����DNR
}Z7T���^x0���F,��mZ'Կ@w:S�TQ���1a����֤%�r�Cd� �Q��l���w�I·
�N�^���uTҽ�N�R�R���X�c\j�2_l��k��< ƯLE+#&c1�?���'�d
_������Q��Y���S^�f�o풧g<_l��� }���(cy���ᒲ�]E�g7aa?�q�\}Y�aѰ ����6 �i�^AtF�%��P�	"������m����T��k�݊�q��wdg	|�K�k��X�s�AN:�wK9Ϫ�����E)<�(R��d0��԰��X�85-���7?LOi�Ղ��e��̈2�{�\����
���s��S�B��T�m���@|X�A^�{zG�_z��Z�o�`A��5*gw׽/x;[�@�_�����X�k�V@���[��aME2��E���]\o)".�fa�}<�#�A��+N�I�J���n#C"�7C֍6Fc�E�|�b{�?uM���b�p�A�Ez������L{��rH�r$�,rg�n<��(*��!�.�݄b������9`�����@@���dmg�0eSyJ{��O5��������&5�ό���S�.A�Q�uj5y�����4��2���$'i�S_ov����g���6J$�����ܓC�4[����s������&�J,���7�L3�P��^�*Vl��2���?B^Rh:O�S��7Z׈�~�]U�ߥ���"��Y�&�xp{�h��}+�ǈc��U#������U<;4#vz�$A`bdR����PV����?Y��we�"��Dv��>���4��q�Y 8��ۼZ!)�kS+Eή�'�2Բ���\�B��b$��Y,#(8��A\�+֓/M$۾zj�C�S�����������̾��Y�r�|*RR[��K��㡫�ÛM�1��$�$�]��Q��ȹ}u�ZN�nϰ=�a�1�5��=\!	0W|i�}a���DWO?�1���^�D�r���h���˵�'��VN*���a˿���
��=��`į�׻`ɰd���Q|�%)��P�q�D>�%jd0�A��qxU��z딏y7E��hi+ �D,�ܽ���3zXK����aw/���j�B ���rJD��:�=�3IE�@�ؠ�6�҇��e���i�"t�W��H�E�8^��P��>����Z�\�CR�hJG�=�|/�0<�n*����;w0Ӣ5ɋLĤ ��t
�y����z��]
�k	T~�EpL���cԗ�F��-��w�����$T�[����]�O�T1�!�!�^��/L�JB��
g����6��Y�'E�v���C����U識��l�����+r՛ {�} T'{�����%叛�H�s!��iwK2.v҃%i9��p�tza�5�A�(�����ANix:�Q��|��w(�3�3�7}���ݺ���z ���<W�'��$l�s��$]&.'�[�m%�6��i(�_��|�nS}�\��(��Xƽ�5�-�j����gn�j�s��P�2���:%`���~:��S\�p�$~R���ැ�ͬ(��>���hk�{s���Ј_�'��E���<����m������_�I9ʴhe<ɹ�.����S�S
�߆�.(��h5�M<� ���Fi�1s�A���ݙ���W����F`��f�伛���Sdʻ���<
mp����r@/�v������fW� 6����گr׃-�����_���6Ppɞ�V~�ܗ�<2 a�1ŽJ��(1I-q@l��G-ef0�߫���1���'V�; 3*!Yō��Z�r�9������i�A*�Pϋ]$�p�<��@\��˩��`6��y��n���j�%��C1��ӵ�_�[�	 �ӺT�/?(�'p
��ˠ�X�;>0N�f���$��J�����`�v�:@kcw�G�#��Yh�OԛWk�d��/LX0DK(5���bӃ�n���XѲI�H���ģެ�#��h�A^n� Urx�9�����D��<\J�y3�&��Ru�z��%���S��Y���}<�x�\P�S��O����H�Q3�Q���r��a�z��>���`�)Q�i$k �Xb��[�Y�-'�k�b���L�	�	c��=��	��ӆ�9[ʠ����<l`���CkN;�rwG\�bP}G+���F��s�`�K'h���c2?�8i�Y�g����k뷮�U����C����Rv��i)�2���Z�(O{��P��%{�ߺ�耇
�:��RF�ѼЏ
�M��VQ�V����*^z4t/{�U�:6\Cam~  .�OF[G�J+:�Y���D��>����m�<1�X{��b�d�R���k����E�MԊq_�_��fz�pӧ�9����g�+�F�1��'�p�&��~��pC%����Ж���7����v�h��2҂�zcr]?2�;�����v��ܿ��b���1v��/����" �-�ޔ��^[p�D�q-0��b�C�ؽSc
+%s0�+��
|�?,���Dg�(ފX�<,b��哮�!+������H-o�p;�uq?*���E�d�A[�E 's9��2����q�J�c� Ҹ��L}����#o<��d�A�V�e��~Q�b��س#��/���W���7���ݩX�2%vK_x������\V��F*�9�;�a?�{��S��d���ɓ�k*�CZ�6U����2�Mx�=�ڗ��@wM���w��_��4��)l�|��l4��E��Y�Wn�Q���n	��Z����+�쉴B2)�
�7�|�I�v��h�+Y3 �䃓�V��i�|+bZSk�t3�V�ш��/Jb�g:�'3�=�n�^5��p¼3=G�ͪ�ܝzصx/Vg�$oG���]��hV�~ ��Ϧ��*�Q]k�FO�쐡����b�Է�8{_N�uP�UܐkJ= ���Y��� ŅRn�Q�h�!������~�6!?j~A��v�p��n���}#,p� Ĭ�i�ln�tV����d!��`Q'�?�o��x+Ҫ�N�Q�Ѥo���l����k�d����	s뗹��2�(�_�9���#R�l�<���	���/$�C��L�T�Mz�۴*�M��xq@����q�`�ѡ8�=�F�D~cy�lB^*�zF�K����YM����T+Ljij�_Ab{�p&�C���g����O��������c��"����Wy���`KϩI(414��1Mnm %~ň�ZA��j�ӳN�׻���B7�5��&D�MǗ�A��3��IPrN�嫽\�ǛP�%PT(�ӈ�$��K+#���?���Xh��\O3ѐ,U<6�|d� �����v�n!)�waX��Va��@'T�/H�qp����U۴��!G���	׬%2�Q�L6�ʿ�pA_���=�:H�o��=+�\_$śI~� f�b�5j�!�ƌD��O���QBYjQ�~�R�W��;��[O������R�0w�5�g��x��������h�Ɲ!�[�ȡ?±C�)Se����t����N�/6>�i/$!�\�Þ塭*�A�HT��ƹ���Np�KD�C��p���@X���	�����ݞ�s �8A�d�%ٔ���C_����yLrL��J�����u�+���8�]!0i�}��x���6��ƀ�F+�9-��I]{@޻���;A����[�B�5����7-��][�<�iO�
<n(�:l�ʋaK+�S[�?�,ҟ���^D��f����qHS��N%]"K-�xq�P᪹����a"��AŢT�x�96�
[���ӳ�F�����JP��e��;��K9_��<֗OG���'��G�]�6��f5@���������z�ۜI�Y�ݧ6yw�����Ўq;�����-����Y��=���cl�j�1�{[�;��%UL�nh̠����/�f}v)pt"�UDY/�<ָmc�JD0�s�_�v"����M���?Xτ³�=4�kv�24DƏt�Nz*Jy�ެ?x�f	�,�'̼F$�pto��z��-�;C�nLZ��#�S7����>�����>.���^��_2�Տ�GN$,��{����˵��M9����K��:0��j�P���A*r�j��vM��90�&a���O�Y}6%sm�.M�˦�\)��Ce�F�[6�8M��}+����k9%NUk����{�������^y��7`�R~�Smy�� �#��v��IЖ*u�S2J�|�f*���>S�R�RASNQ[�i�㒬���T;f��:�I ;�09���*�SUB�9&�<���]U�^��ʌ�@�n� ��C=��>)ݝ@M��<����.񟆉B|Oe*۟<ͅr�K��	%E�����Yo�O/�B�G1�������|���Ɵ���ݘr�T������̍ٶ̦��+���Β�{�D���~%g��_��D��g7��_���
�+�7R�]&����)�|��&�l5¦wx����e�����,��1s1T����֩� �y��F?���/uD��u;t#�G���X#]�Uڰ:�_�-�	HfG�۴�0H]�t�����b	$�+��K�s��!��n��%9j�T	{ԍ1sK6m���#�S�u CY�����DV��j㣅Tx��UEl+����ݲ��[В����#�2M�=��G��J��*�� ���G(�=�T�FboA�@/) �*5-c���%�ՂNݦőAG��'a�j4�U��Y�ն���BBح��g�@�����*l�G��9����q���փާ̀`�
[���TpN��S����m��0����<a�>{\�jD+7`A��������>.��2Z�'��:�_qp�0�@-bGS���#s�0���H� !�*E��
p!������P�d0���o��	��w�JnG�6���&paҺr��@t�dީm��>]f!1�r}t(� 7��w]�h�U X�������U�,�s���$ϳ�g��ߣ��$w:u[։���ĩ�Z��2,v�ˤG���{��>�7�o��� _5^6>(����j)tx	5ȴ�k����=-���t5�
��Se�|=��� &�R�$��ю��F�wL����Z���4R�s䏀T�BϔU�����$�4�B���a9 ���� �WU0�D���3�?�͚�����"���9���J�-�1��T4�w'z�!��`~�2�Ԑ�Zk���#3�T�)�EK~]����<�t�⇒U���w�}yz-Hie$���I�+�92�-����Az��!�����(y��<PvjIS�Âr	�}�d��\b̫0���!��Nv0�`W1r�U.��W6���q���[��s����5uB��M��XIi�6�0	��[�#�kV����>С�#g�mQ�m��ғQ$�cz����t/��ݥ7��|�l��|��F�E��tKT�;#��s��Rx"�/�\��XU�������z<2le�|o�a��2K4H���OL������g��:���]�t����q9{�	�aR�rlS STo�Z��O�	Ԙ��|��U���Xs�Vh�
+M����r A�N�[�3ޫ�6�\w)�v��OM>����Rt���F|˭?�aȪ���)r��'�O���P��N����J ,���> �䭎4r)V(�À6w����y� ���N�:�;T�^|Gv?V����D���.VyU�脾��q<,���憒��k�T���1 WJQG�cp[�S�Np�	l{�$��hӕ��������`��êA-�����V��I���Q0`m,?�[��lK?}>�
����R}�]�4X��N��Bk��+�d��S˭Q�r�yhfR. ֶ^x�m`kĴ�ҹ�^h�����9�e0�d�-��l�#������лz�L�-�Gaq���T!*�/�%I5�+9�xX��O�8�:�ŏ����@�5 ��z�9���n�Нۂ�s��ףJF\`��[�N�@t�?��G\��z�K�;��(v�\NxE����8��C���y��!0�q��~b)�dɠ6rsЭ�v�(A=+(q���o䮻s����R�I~H3����B�����姲���W�F�bKl�й�k��I��EyG9JZ8�BZ� Tx�/�3V�:$+Uh�z���h���5ǘ�駅 a�Ļ��Y�J���钛=��1c�J�q,�� ̻^��Ƶ1#Z�f��p��H�Lм�����uǢWϲS�Wk����3�7'*�f��o���R�Du�����H[�����l���G�mݞC�+5-����]3����c���F7}�[r��O(��{7�N���9/�
պ;Cgtפ2Z��	�&�|����=Im~Y���=�5	������tU����L�����9a�e'AО�-�,�J� ��¥��d})�?Q�@���JS���YӅ�c�߈�0����%��yd�˺Gײ��J� ����k��rG����_�hTۅ���M?���V�����I�$-Ù ӎ$��<8~ޮዔ�,G�N=���V�[E����N���N��k��sO�r	F bih��gxԳ�~�T����/�Z}������j�G �%d��WlB	�G�	�-�+�M�-��J*0dDe�%r�A��tJ�m�<:շGHU��s^TѰLՑR��-����zfYs8%�߆�̀~)��,���j�b���y� Ɵ��\Q�a�&�<~�������i�+ ,��jc!�MS���g�M�,�z�m��δ���{q�0y:�c��ǒ)��ɀ�ѰR���0e����BX�C��Jh4#p��B���]3'\��1z�P�;�
R���z��:Frf�R9�7aQ
ђ�h��a�O��7*@�|֯����QXM�&�9��/��[���`୕Rڕ�����d�v�1p��B����C+^&��܉���pV����K?����Q8�\����l�s�1�"*����E���_���M���ߚ��F��z�"�Pߏu*���i�qZp�.:�9  0���,�ȎMG�)$wDRV����T��q1����F��r��I�3`^�������}����Z�7ٺ��n��4%�n�3n�F�� Rd�ӝT�F$腚9n�,<���5D���*���
���+�c��6��y��z�����
��3�֬�KEW:2���`�:Ɲ��W� T��S�c�  �O^}?�'�(��*.+��2�m}�j�����c��_�` 5�8�K�kkԋ�]�'hڝǓzXd�����Ep�+,�!�oQ���Ң6g������O��"�H8{�R�0q"�,�BA^�D�u�hZ���|�Hұ�l~�o��\���������{�*b�S�,���P��J0�1-侥�z�i���V��6K��usx��F�vVBt���ƞ�ed���+av�<��C�,!��̵��xOT�Wk�4�h�aǊ4�~����"'�|���O6W�d[[�%�qS�f������_a���5w1����i�a�MC��Y+ڌk�I�YġSh���TMRRGys#:I����ŢY��˿_"vv�f���ǣ�_�ę����ұ�����k��?�Uc,��:�ʴ�"8�U�ԆjN��J.��5`
����v�U~d�Ԍ��2$:HWZ���9�c�,����$�������4�v���^��=7�p����>�Ɖ� WE�G�$5w�$oE�W0�y� ����<��%�pw�A��R�^�U"�0HJH�{�O��[j�hW�D�+���!���o�ZQ�$��nm؂���;/�8�r�D;<�M1#�;�2���6���	�Y����pۃ}s�d�CvD�Ų�2ay��c��؇&�(��u����z�j����Ci8Z\%8�I��>@���w�=�'D��0C%Y�7@U�%N����\�T��꺹��!���/[�fxEc`D�ޡg�$��UfbqA�y�O��U�����'&�1핼*�v���z�g��DW���1��=���7��n#E�6��lm��Й���P�t���A�/�E���ʳ�Z�a@u��B-���ü^a���(9y6hn�6=C�U��_�%�ےd8S��yԄ�!���{Y�����A��B����������q`h���5����C x���{��t��j�^��׫0nTJB�����]���~�e��!��A���� [>���<��i^t�����]��R(������� ?s�O�<��ꌎT��WD����"4�<� �'�E�#(u���8�)Hu3�/"g��s]��I��2f#�$E��2u�:�Y�=�:d����~a
�ø�=�ay����X��V�w/_�em��c^)S*\%׆���.@�ݔ�_����"V��K ����2R����w�0�(��6+:�����L�h2�Ʊ����yKN㋀�$l�U���]���2]�!���� ��$f����L]hy��A+�{�����ju��7�?�鏦������n%����j�mʽ����ХF��F)�����n+6d�餒j���O���T�c|�ZEh\Ș1\��R$��=�#���	+�R�����]�򄴤��Q��i�������o��8�:n��-\r F��+#�'��KQ����8�_��f��p���m����ѯI����љO*О���F'];肙#��w�5Q�4F)sTҕ1Y�buqH~��TΟ5`UH���{3��z���1`o�E�v����d��;��.v񊰤]In��5��h@Sg�Uƾy���������
�E1�,�$NZ;e[�0������H� qB���O��:�3���<#Eku%��F¸>�1���:�V�q�sU�M�1�N��Q[��O�0����6�*��@�kd_�"�^��(���<��h>��h���ʔ2��U\�^�V�l;�G�כƮ?j�a_f<V�q*�2ݑMs�q�6#����1�]�E�tX�ФO�L���H�U����=DN�ֆ )� ���ɿ~�s�=�(��>* �n$��	��(|xx}���/�(E��:�̈ĉ�9�mp"M���ORx�5A�kA=\���`±D{�O�:�~a�Jcwy���<П�3�S�؋��G'�y�cY�Q��$��䲭s@���>����&��P0���� w���;�$�����,���C�c��A����!�a���xC���8B,r���K�%w��K�������9�в&zyed�F�?n::^����Gq�f�Z� 4{e"�/	\�(h	"�{,v�u�r�5���B�Wi�
ro]o>�+�s�9���f6�l!���^���$�\�N�iLX�Q�؆�?���6�؅�����A�n�+TCI,�X �W�����!�y�%���-{1�sW�ݷ��-�g�Ma�1��"�@p�u���_j����v��'��"7R|���$��WK���m��U�Q�]
Jy��<�����G(%!��:�]T�O~�e�vCnS�#g&I�`�{��^;E�-�C��W��Zc�|�oQ��5}��{=!��.��P�U��Ч�_�u/N�\]���!����~�/l��u%��s�`���.���_@���	�"uJN�+�-��NN��~�E���$�Z�\�ugH�l���sh����'�CO' �JC��<�1����wu��l���؇8�Ϩ�e��(hiS��x#� 1�<Q��&)	�6��H[��.⮘�'8Cd�ˉl�TjE;0i�	�PP��~]6�/ǣ�e[�k2�9�� ��X���ѹ��t���X>�L���[�2���-HzT��W>��W��{�_DO�>/c7��QE��P|$o/���/�W�]�����6�CSs+֍Þ���k^l���P9���i�B;��LC�}�j���P���8k�����sƆ�w�?1����A�^U'Y��Q�,��tmRq���Z�i�ֺ�w�>�/�gԿ�q�Lᾖ�`�>���؞��j�W�y�rm"3��š��Q�֌�as��P-<�7�aL�e�M�?�!�<��s��2�EB�K%L�Ki��yr��d�b����z��Y��N�a��D��à�>/S�^�r2�]Ii
.ƕj�FcU~w�{�0nCA�0�3����D�cWןl-aG)P>\G���S�͞}���+��8e{�T%�a�
Y��uo���{'��#7�����SO~u�^�ɹ#��}���?�m����0��W�s�ϖ)�팞v�I���J��}���pj����pa�=E 3�_]�K���7�To׍�x+K�X�Y����x�3��L_&����<%�Sn�;RV�����6��9��k����*��`�'�#���O�:�JIt�Ѽ�&�^Tb����r�����ͽ�N�/-A�O�`��;�)�Я�S�gɕ!bgA(��˻����!�g~ӹ�������&��%��|C��*�/l�+�x6Է+G��O
0�|�(<w�d��y�W[<0���A��v=����"!����z[ ׻x�M�W��[�z�o�E7	@��1��K��v&�u�չ�����!l���q���ER���~��*>��c�*s���#�xEU��U9.9��Ko�����>2�7��e�F�.}�d�V�������i����VK���y�&���<�琻#��z>�$Z�X�8�`��t,'R�	�2�!�B���3�[�v����qoҬ��xt /v�h��J����z��h�o{������=3���$x~2ZA�Ί��w�[��&찳f��].��
A��InO��a�S�����z]D�*�*
ᬠ��/���]����X�t�����I�%h���1lݾN����e_����1��/�U��AFM
k�s��*�ˋI�z����SG���?ó��7�%q=��м5ý#� <���3JΆm�W]���: &��+;��[�Rn�<���k�|�*'��.}��6u���H"u"���p�:;n�*�O�풫}���"����,�w���p�����n�V?g��xY�l[�6�<�AG����{l��sCy3V��������^�:w.��纕:KE}��6��zEoqV:�=5e�'�޶�l��#t��5��_����^h�7۩jq� ����F�<6�U۴��~�{������{n���B�>�C+��9>��Í��!�T��lI�N~��(1��8��������KV����<��+Wv}�~�A����LH��|�w T	z�m1�"��vy����pڞ~�R?k�(n���W�شN����ݻ���b����Ն�6Q��B��O�W��D �⚓ϱ����j��[r�$��[��������RAl�إ�P>��[�cY�_"$`��u���]�>j�ʢ�F�;&�r���uh�?[�>��R��Zy�R|�u��9�-��T+�"Ee�QV�IS��1y�Klk7ԑ����FY<�ߣq��o������͙Ɉ�*�&�üa��{��p�g$.���q�M����&����A���k��8�y�i��*��h�	��yW�#�|yG�>F�a�Z���T9�'�g�����j����R��ֻ���
�j#8�P(-ޝ��W6>u�ʣ�0Xc��N�FÌS@Y�!��'��������-�n�7E�o�<�S�)|IP�_>��o�G�Kd�D`%T������H�y7F҂�u��I3
�	�[�X��P�6h)SD����}��Lf�%X�_j�)�;>pK)8D`��'/�S"��t A��	�v���ݘRː�`�vd���8_�R~~WgK%��Ej'|�;��̭�����q'c�V��B�ŗ܌E���8�% ��������z@�
f��.���1�f`��F�O�a<��-�t��&R�<���v�\_�`b(�~�<�}��e�Uo:������Q�ٹ+��"mff�˶6X��*X�t��˴6}7Qo��B-�BzuQ�yb[�ݞ�I���৛�^<�4�M>9D	�i�jy�"����W;EZs��P׀�����'S�ϝ��5�a*.ˠqG�%�-�v�O��B|
=̀�f[3Ԭ ۡ��UAJ��4�o�,�oc������O���D�̲�d��=``�Lذ=�,˔�����B0��>)��0<�8�*j��*|RJ��f7�i�IaVb�e�K��ih�������
��xOO�F��t��U��H�����iR�)]6DW8/��|����fy�B"�y��n�i�}�JV�Ӣ�N���"|�$�p)��\���cZ��?�A��꣠�w9j�7P%���0�>�dV��/�Z�� X
5�ۏl��4
t�|�ț�׼C���GR�Z�.��]ên�N��e�quiwQ(	2=�.���|�����4�+�uA9���z3h�Vf�v4D�}�/c�BE^/���Q�<o��E��0b�.���bKc�����b��C��G�}�jw�> ���j�6���@	N�j�����K}�����O|�Ȋha�޲��,�C2������X����[G2���3�����=�f�����H\�6���5s@���{����c��y �9SYը� -��;�Z=��}:ͦ���ݬ ��\\��|G�_xy�ǃ���������q���^/+]�� Kz���V��#}�g�P�~^��4V��(�5�C�˦��Fj����(�Q�{H��ޗt��u��2�Td������Ԍ	�_��*���U��h�҆_�際j�
lc��ZΡ���?'�#��,	�(u �h�����[�2+��D#uU��jBX��}�'	$Z����u�\d�;��R3՜��&�Ψ�Pӷ�7�1�ȸfN�=T�@�k60��Ԕ4��� >o��Jo��Sz�<��q<�g�~�����^�������;�U��A�P�V\A1�Dk�Y�S3U�B�ai�����{P��P�vs��I*-�t�@[.���G�؉9�@�"�(lǻK�qїG�s�[}d����mn�X8����I\YWK�[	¥X=�Mݫ����
�w�ł����eZMks��$�
��L~=�3��`O�ARZsC��E�q���N��b%?m�b���d�n6��s����:z��;޳e��H�t썹RQ�'E�/&�qe	��<�p�N@��C�����[.^&C;D��B`�"�����D�ǚ4��䃅�HEw�cϾ���O�3"�vϓ�s���	,��X?���m��E)s
� B:����7u=cQ��_����X�t*�]�e �[_�D���,��Լ��'[��!������3�K�3��a,���љQD�t����;�ǹ�f��iA��0�w���^8B�m��#�w���C
H�_�"�3��
�r=��'9�~�mRx���>�`l+�̃A��a�
�ʱ���A��C]=TiԳ'F�ay'e��3���wϋ*�{S���~��)��x�ي��fG����@�ǈ2�|g�����O�Ee@8 cC/����o�ǲ0j��f�#�w���|�5�l1�)�f<4��X9�-fn�C�D��Qo��Ղk\Q �^2U���OCy������?�v����*P���øI��4FeK�rG��0�r���\&|���(;�#=.��dP�4�̎��cN��g�W��!b:�ݣ��_��>B�,^Q!�#�����69,��i4�=�c�K�_��r��dg��*�3W8���7)����Nk���F�v!�ͿM�[��\;�{w-0c�{���n��XQS�~9���Ʈ%h����P�>��ԇ�gye��9�F	o�l��&%E��A�4|�<Ol��x3��2HV��G��PD(�>v���㖋1L���������(��5���[��.�����r�����ˮT��L��FT�Gu!�k��,�I{2~h'�6=�쒡�pF��2l͘n��D�mTH��]C�Y���a����;v�8A�S
42㻝=�:������.�\�I�u�a{�Z��0�[�w>�n
P���?�O�牉����P���M,ȥh���ڳ�&�G�+�
��V$�2Wۇ�����~���ֶc	��
��su<Ь����⎟w�U	�G��s�Gf��B>�,��Ue�୷�L�Iu�x���7���,U�T����%�*x:#����m�vT��+�����W?[��9�o!���-&iS�;,��LH^�f$1��#�0�t�c�Q�;��� ��Kn�NіF�9�UD�`��r�i�a��A!���*�K��s�N����T8�)�y��`�aѯr4����=z�ը�k.��P�������H�xK'���N��$2����|V(��QC+T$}�n��j�Zd����о���Zo}(�Ig@!�{W�Y�ᜇ�%� �#���r�W�-N�:��[n�nF?��O��R�e##RO���E?�;��m�]��<��
���HY�A�z��<�5XƤ�K&DшB��^��y��O*�I�kQ�W35n��X�ӟ��ˉ�Cq�=\ӊ᫵}\��7���ѵ�m9��s}��
,Q�|frɺ�n[:�T�S���$�:d_Ijs�9)��[Y�D+e��h#K�.SfqD���ю���z��{�;�m9nݝ.�r���^����sR��WS�j�� $0��|ZH�#��]�{7"�(܉9��Ǚ�h�X���C�X�'�1����b�gw[#�&�[����O����j/�(�,H�be:��Mss#dQX҅o��~wmD���`�|: �M�ڨm)�����*'��^�|]Hp��9�N��lS��w�N� ɮG@1ʤ\)���+6ֱ��;ѣ�(L�Tn�~��]�e�
���s�v8*�m�����"�z���h�]R�T{_ i��x)�"ǧ&�����M��P�5��b?�1&G� ÅAꔱt�R*�7x��+ ��o ���b��72z12���n�Y@{�E/=u7�3����Q��޹��B�=�v&m�I,Ŵ�t���W�j?�,l��*
m�x�1���hua��|��[�ف:�S{Ʈ�^��!��/7v����4&�#��V� S�!�}�}�XO����4W$$����鼉���c��%'���̪��%��=�z?�F�Bؤ����̛��eI���3�W�}��O�4�(Ndo�7t6(3���4=̈́��u�K����jq���d��So�aB"s�o���;%!��GG�|�ʢJ8��h;Xe*�8��%����x���5�T���B���� B`�&g�+yRUKQ$a)V�}�l�G��m���n����|/_V/�"[�f�;�zn�s:J6�~�=�ZҳOw�x��f�*���_a�w%������I���
�7��L��)Rp�S��`G�_m}a��c�r[5��9�p��iΡ��J�0 ��g��U�`y,���"��\�����斢Ξ1}���R~s�|�u�"f�fgN=��Iw�l��8�T7�.��)�
PF)��S���X�����h��G��\Q'Y	^m�m��a����	{�˟hO!<�s �p�]O�v�op�T;߽��X#����"��`P;~;Z%��#��K��iWU� =M����E����NE^�9��_��OP�����*��E���U�<��3�Bܑʦss?�uv��������85�"����ͺu��c	�#,���6DQ�@���%�@\7?�g���9��Q�W��o���f�+�M�*�1]��Bh��S2"�@����߉�"r�M��&�db�ν�>�P]�_ta�25�W��`��0���)����G	СT�D!R�^\���eZԆّ���c�?�r��rX�rRH	����A}�{�,�Jp��>�0�p�ա�G�:3��������F�B'9���Ra�&\����	��[�{��w��ſ/����$�nQ6e;��>�s�9�.(3�74ooY���Y^c�9�+���uc)E|��=�⁇ݞ�.�G[�X���>�E����i�8�����BuVqn����i_��v��_F���k�
�4(f#[2��_һw��]������<�g�Q��N�>���;i+�Hg��k�B;��;�`��1z&K�8��x%�d�3۬�%��$�;k5�lK�F� nֻ���,�6.�솢Ǹ�3��	S�zn����'*j�$����bo��S���o�q�c��S���?#��5NC^��^�Y�l�5I
}�4��{{I�*갷r(WKb.���Nz�L�6��ӷ6����-
@���I����W����u�f��MIdh��� ˨gر�j�M[*�$��x�)�Y����c�4��!�&��A����+b�e$e�a��SL	��5��k��N=�r})�|���ߺ��#�8�xf�P#�Ml���زK�"�;��s�k�x��L�O$/�r|}F�x�U<�0m༖O0^ebh0Ⱥ֕�QH��Ϛ�����+�1a@\�B�>v�O�ڱJ����]�D$�z�@�sŽփ2�(�;�m��@�A��7�(��U,G�R���z�N%A�lz->K ����@.�l �P	��~E��j,��a�T6uH2� �dy�yT��?�'��R`v�3�xa ы�áި2l�53�����ow���Kc�+k��`+t�.O�M��k�"�&��(?��[�H��4i�ɱ�Ġ�x!1����S�/���*���|�%_��q�:].�wNE�:�b�Y�̰�$�{��.!J����_ftP˹�-cpm���].FT�m�#�����^��_}�1%ݛY��٠EQnĿ�1��sfB8�Ϡ"��W<��u���E�����
e�Ln>���򚲳�T߁��Nr̝���D�<<�N�'ZwARC~+iel��)�Ғ�ш6}2Eg�rFc-��"�/�Y��wd'쟉�|F+�RA�n���R�ի ��ք�9qR]AVo��'}7��߁I��9EGb+�uJt �Zl��ߝ{�zA���vq�P�2xo�tjR4�@���*p��F��-:t�����ߢr��I#��: � ��>oNmPc��Ȗr�����)�NZa?��"wj�5 �����	�c_���
�Q��V���x��[c$�үyH�mn�q���>F�]�������PW��"�s�U�?�|����CbĖ��������m�#01s��/��8cW���m�v�
�6�t��o���^_.�&���"�e:�!nM�-kS��;s+���f�EU�
�+'$�I�Hʸs��k������.��?������Q� �`�B�7`
�p4�rlcu�Q��P�d�^$e�BH�j裹�.�T����/�S�A2Z�����JV"�Yh�]�pb�eL�v,���h?_a���W�5oB�p[��>�i��^P�K�@�V�%B�4��a�#oFCO�ܖʇi#�.����:+�j�JSy�f���/h~6(�%��s�ҿw�+ɾɔ��̸`Ǵ��P$G�%Zxw	��N_�̕��51{k?�IV�}~�!͋���̋	�idX�O����V����P��c�k�d�#(/)V��g,^ЭH{4����%<?w�����ڔr�K[R@߹%��`W� .(�V���o=�S�*�}��L �����Y�����aƿ�<鞵��Br��Tݽ��jbNZd��)�Hcw��?"�80�v����b�f%P��[�7��5��G���3S����:�fF�5��C'@�x٪�"�1-LHw��-7�hF���Ȫ�"�;��߳�����C��e����$!��kV�#�S��C�C��� ������B?ti���4̿��5//�;%�A*������%Q'��It�"E��<C*Ä��Z��TFѕ��aқ"�|E���MUO�LYB��h���2<T��7���n�|*�?�\6,��p�����+}��~1F>�K�W����Q��
b��f���~� Hl�t��:�S	�g��5 ��c��@��"� ѐ�����-	p#'��:���DkB'އb�7������t�Ko��-߬Ԧ����uo.�m����]�&�f�{�xYE��d�8tsF������������7X̚�N������+6w�Y�F�%:H
%@��-�l�{��>Vl�ۢ-��<(@jQ~�
;�a:���X,M�	 �^�]D�.1� �d��b����M+��@��X�{�ZHV�:1��5����GÃv�0��h�-�Em�(��qj4���[�D��#�s�X�A���`����VW#�����P�u��+ab%3(V�;>G��J�b5��7Vw�g��/.�3J��7�jp��	��М����f�4���}='�yH'm�	C@Qx�]�!����t��e挨ஒ���~ʄ'����˥�=OR*� ��7�0'�-D\T�w�x����b�wZ�8�h�v{b�B��:^�ѥ�2�O�.�LuĽKf�-!��*u�)>��������?����Eƣ{EF���:s�ߗ�y�[� �K!�P. ��)dH=���u6��M^�z�JeiLli;?Ҟ���P�/5�0��Y�����w�&Z�&7��@�@�^�T�g-S�� �ۗ���^܆q[�~1��@9�����<��*�RD�X�ZSMA�^Δ��Kw5���P���:�+����(s0�4M'
E�]6N�t�+VzAgv�S6��9riP:��V�y09c�亵��;�L^/+��X�j�Cڎ�J���6s���/�qpFN���G������W�/�#���'�@v�8뢠=j��P��t�����G��{#YF:��.i�g+��A�(~��Da�b\`�������A�4��˂� ǟ�N��J��ãr_�/�\L�x����K���h�>� �v��f��ݱ�r�P����?�)���.��_����nb�������-�w�7L?E�����������.�e��)4�PT�L�y�<%R��Ʒ�3��Aç����:�'f@Ñ�b����?��h(�b9IKn���r�A�S�W�
�ZVb��P�`Seٽ�?+W�?�s~�cé�ci���r�+ �6�FՍ�5�m��Ta�i�3%�Rx�-����%��m�6�x�2�4D�0m����(�Bo͇!��:kXY l�>زd[_dV����lb8�N� �90�l�{-PM�-d��U�}!L�!��o����J���������b�O�B�I�h�B���l�;�{���'�
�=��J��C�� 5�+B�_/,n�+v>0����j[8�cg-����r���F��bA��[jv�惫y�6.{��%|���^a�?�F�$���-�9�+V�c�}FA���O-z�KE��9��2�� ��7{X݉��c�"�h3P�Q���d9�y�Ɖ�TW������_�>�Qk�����CL�>h��(�P���P������։ ��L�Z��TK�^ �A���T���UK3]����j�v�6��� �D�E$�;I7&���%���Q3p���m:��e�D%�avh�����ɦW�#�(�/���+a��D�Z�^ԥ�;ã��k����G�f4�j���]�z����v�e�N��g��avy��>��T�=7sS���6v�������L������Y�Z�q��-�s��ՃlL7Q�sfL�UU�͸�ڒ��9��O6JITR�,�;��ܗ�'�	�p>��x�U��e:�X�8�y��,��ǃt�����7R�����T�f~����%�z����6�*L2z��?�Ҙ�����ܠ}{���bbwl����X]�yZ�]8K�0�|����GI	GӾk�mcM�ܵ�lӯ�E��`&���I��YB?D����f�;L��[��B�HG">u���	��x18Jk�4�*jR�w����o�!�DK��H:YH��V���W����Z�溏�tnR�2�>p��Y�~���j���%*c����3&,��W���]����q\%4]�m\/�+|Rۅ]I���?;(ӡ;2�
�
uMX!�^ȗ�$S���hO�+i�|s˶� �V��k8�߭�� �0O�l�����w
��?�B�F�8NC����`<��=��x��s���܍|�j�`xh�	.B��%@�����{�c�-�.�[A�n�,�����y����*��sW���R���F<U�uj���p�|��K��\X���Y���ޯߙ�zmoWɜn��e]��%l�n\,�ZI[9߳���Vͼ�l
��Mz��n���s��W�<3�?��+�h�L� T�X�ܺ)�%�)!�	�.(V�w�����L*t���\2%:�L-o��͘ �8ڧ.�����-6I3O'��6�~}�	o�㍁���U㜡��2�~`.�+&)�~Z��oҲQ5����:M�(�K��լ�a��c�H��>@�r ����ɧ�i�
d g����Rc�%a��b҇P�&�n���І��w��*O[�5^$}����w_�Q��bk��}
؋�l;�g�[F���0yܩ���j���i��O�S
�rs�.�O�IMy9�1��:�+�a�A�D�F�Kn�j �\\�l0�]\��z1E�J}��<�v\)p��Gt����ԏ�`2�����+/9R�[��zb������!/���^�}X��ҳ�El>EZ���N
W��ոZ=�(N �8�<Q�9� q�_�&�:y���n6C�{�je�JUU�f�Z��P���{��\����P��ivt�9��p�Cڎ�D������mIX�e<jZ} �杵�A��������
c��>��P�{�\'��*��	�l��哯��5��}υ����_1W���j�Y��`����w�V�^seE�CP��ԯ^[�;X�1��Մ���Z�e��5q�<2pQ���w2&:pa��.�J��
u�yI��kNc�g��IN�ir���/ri���\+�b3���xl;
�%�Z�H?	���URn���XU�_<�F	Y��D�>������*��d��0Fw�V��{����hκ���2�鴹ګ�����sv�MC����C��oo��#���9�w�x��]ԅM
�b���kT�LL-�Ln���3��J�)0��N�\�D�-
0��c=�+VF�E�8��+Y���Q��B���c&1�Y��R�c'��N���x�j7��TV�)J�f^'��qF��H1�`20�����f,H�<���n��;:a�ۍ$ǌ��ƌ���M����=ދ�����ŉ��N��< K5��<�w��'בά=�#^�T5gO�/ۃ(�/jH)���Y�����q�ZjbW�'c���(}{�w�H�Ѿ�V �E��A�IH��U/�r�>3�$F��Y٨��PJ�]�~��Eh�K���\�)�X��Rr�BL�9��%���>���2��M���%�M�@���b�[J�����MRr� ]��E�S�a�'=F0�9
�A�.�|�k�:�����Չ���B��F�6n�{x���\~��99��pt���s/�ep����X�9����@RÏ���?�T�t�}-�[)i��$F�Lju��R��k{���#9�9�e��S4hO�o���;� �r�����h��K!;�a�^�,���^W��sj��3���T��kv��ͨ,�A{�~z����X��q*�Sb�'6Y�'�ߠ�ntdR�w
��(�����G��2/�8�mK%߻���N���de������.)���I��Kny��Ӧ�͂�4��qͿ�CU陉���I"������v��zN9���{�|���y��̳�[�~�y���J)8������a��䧚�ϡ�к��w@))L�����v�`�R�~O8��࣭8�Ƀqb]�������Q)��f���M�opva�Ί�b9����)��%��'�����[[�2�lwH ����.d�=5�px�I���Du��l-$�ӲOZ����O|Q������D�[���foA�6��L%I��O}��8T�h)�g7��JM�W�W����zo,��L&��<���!�kgǴ���g����y���)�t���+K>����㝔�Vʈ�F��;��(�Fa"��t4�E}�64qOlxjK�yMv�o�<�~�dj˫���W]�b�,��f-��L�>���k�:�<$�뽎��e�	=F��#���F��Kޚ�8��Do�b�\!��!կv���R�G�N�$p��F/㾌3/.���\���dS��!!��!�\`��܃��س�wϓQ;a�h�M����(Ԓ�� P k��a�w��n� ɀ���T�e����ע��Nn}f�)�P���D��Ǟ䪱*�yѤsz}�,���w�k�=�0�g|���B�� d��Y���,a0�Z��1���� B���/���*�`"x��2Q.�g����$��o/�����4�lAP�|����P^G��I$#$)f���ˡ�|�0>�?���с�eP�
��8�"� !���|-�+W��#����h�d���"<zȶ7�T���������f]�_�c��1fr'd5��obQ�xL=�2`� 톾�7�W�He�M���F���z=��1W΀�R��I��<~�of:T7ؼx�2v-�Ҷ���V��"�cȘ��e��
�ls8ƹ/��I�l8-�H��&�{W8¬o�$v�/&���fDji�#w�h��j|�z�!�����Nt�L�z�f�*�H�v��pP�������#󺫺��:@B�-�IPq��v�jX`wt����1�c��'�7�#8X�9��l�:"L%Ҍ8=��o��b�޸h�������;s_kƛ�M����d����i������T��=b!���7vֻ0?#Z-�aЮ,��̲����;ӳ�{j$�;$�����ZI!�5{{�.��C�p)����Ļ0��d��J��6���$C��R<_ȿ�ڎ���u�FӃqQ�&U��.�����&֛i2ϋ;l.�){��V�����zR;
�.�wM���d��6qʼE�Uh�IP�.�n�ι�8��.А��t{Yd�'x���l¤͓e���"��|&@�KO���d�,W.���m��,K}���N�xl�͵{�Ë�}��](%sS�����Sc��Hi�eG�P�[a@B��ƪK�խe�3�{(#�us��}x��Dg#�2b�Q��l�� �?�,vSt5�������|^�� #���y>��u�7PpY"��N�\�t�-ޑ��s��40�wH��̔]�}K	=�XY
8E����`�Q�]�w�����wa���2��
�#iW4%�a�h��n3�#s���N�B�f���c�0���7��E�{δ��L�!�{̙6�tg��2����1i��O@E��h��g{B2&���m�"�=������?(�^(@�A*���5! �O�0r���̫�A�bJ�PW�gl/��?c��;�L������RrT8���c� 3��,$�F��3pJ�&>i�9��cd#�h����CSF�� Z&P��yذ7d˹��3|��[�3�����p}� �	pRY�y�1TO=�$k�:_�,P�V���kf���		�d�� r_�2�.YN)X��[��r(��&�"��"�
�{ɕ������N�
�>B�U�i��<	���������������W�CI����Q
`��>�T�q5�����Sw{w,����%��%&�ƽp��zx�0�WMC�E"�@-΢��@_�S"��j�/0Ã��C��r�j"�z��̺u�)�l5øā�`jд�V��������$.���rꜰ}�]���e�5pJe������k�g�tO �h��NE��G����_%���Gn6t}l�]�|G}/��d`W2�9W�{Z�&��Y��D����i�.�����F1���M/0�n4h1
\��=`C6���L�>����)���^�Nj���)mH�7��[!�����'�9!��4ܵTKwm�f�I���7��ن<�!���Rk���y��>yo:��F�<W��L<�����R����� ?�����|�s�F��3x�·ÐF�	6֓��l w��%�$'߽�7�r�t�&4BVOE�{�����r��{�Ϳ����_� �
ڪ?�-e����DD�.|^i��	x	�:D�\w��R���ōQ���@Э�Y;���a�?`�.�D��t�xM�1�9��f����A����"�y�'>��"A&+F���� ����xz�ZO7�HD[�H�7&�V�4_.J_���G��H��u)�7�>3�SxL��硪�O�Q���ДK��M.���h��k���B�O�f ���aB�8�gB����Yv׷�x��g��� A2J��·`����n��4��lc5�aH;�#��x��n!=�?������9x#G#�z08�uǆ�������qW�a���K�s��^�������%L�˗fNHc�D2�}DQ�,<w���1%��=l Rnn���<Xq�B�`e�G�����˼�D���j8W>i04T�{�G��i�kW܁Kɝ��xm���Jrϥ��tR���q��0F���(}5<!�2�o�-�����fy͡��tբM��{vsT�d�}Y�8{b#���۳��7�R6k���F�v�1FF.uRh(���œ���i����,N�!'��?�5j�j���+�����PPvX�I�b�4��0�1$ԁZL��[D�H�����pP�9ꖪ�#��j5a:gLV|m��A	4����p$�䥣߾UL#��ר�r�e��QDS��^�D� Hx�xs� ��Őx�i�$�t�e�5��/A��Y8�D�r+M�<W��E�r� �A�R��W;�	R�V�c'���1��)U=��ڢ)�ݵC>��
�����@,����I"�l���4�NS'��M#�0[C��9"=�0l���8.L���R� S��K�������RY����I
�n��ehai����s,�Y �8��yEU���WR7aV���<7�������׶��I9Z�3JA�U$�q�0C�s���	� ��eI薿�w�,�7��2����)@PlFXj�P�C啤$�=���=g��]�T��ȋ��2;��N��6�a�P�4�FT�W�9r�ci�$���}����1 2z�����X�Bj{�i��ל��������`!�'!Ay>�`�u����2� ���S��?NG5�x�z�U���7ύ��aR��r����r�|�V�R���߆�cY��g��0LQq0ߧ�C�F�xW)k�#�4�틽�*��/Qp}9gZY鋾��O����X"B.�q#��}_ ǒ����[��F�Eog�4�q��u�C,�&rf��CI�+���j1wk�vR��� 9[���kq�an�~�"�E����:{#I�r�3,7>�-d����;5.��Jɋg�t(���/h�D�)Ps�	�������pLAT�[�C)^��뙮�K�/3��ѓٱX������5mI��Rc���A���bk�*Q�g����j�H���͚��m��[Ƃ���O�f%���븊���::qօe�l	卻i�y�_��;���Z>��SJ��I�����W�'�8Ş������r���XQ�Oˤ~�����T���z	��Ƥ�8PBk֋��.��Gf��\Zk��Mm�<S��/��wҿ7q��)!�L�}��TkVU�
$�_܎�J~��]p�ݩ�������� ����:F��X��ֿ3�J��ȘR�n�^��L���8G
��Ԅ�T(��,HP�`,��Ή#m)äx�"&��N#r�8|D��8��ʓZ�Y-��*)��yp
��4e��(�\J�]p�P(׺�َ�����M����X0}q#��'�L�m�����&�&[�i������æ�(�U��\��ӎ�.��	#�o�A���lq���˭v�����x�+8�K�z��P�wt��Υ�d�a����CG��}�s� �@H-�mYEK�K��aN�'T������l��}��O6x��1��u�v$�O��Y���Zb�"�,��[,P�ec��N�bC�u�J*��U��g|E��_��\�p���0�P�O�a�P(U��N����y"�||�deJ����V�;��0̰�7�;�z 5�����<GWd[ŧ�u��.�[�Rց�����#��a�~s��Ƅ<����,�
�K��9���b�=��i�.�Y�T	:�{�?�W>lXo+�a����C�r����1�*j�
J!��t�,W�x��&��J���jTm�5�n��#�m�W37��^����g�����Le��4����-
�� z�̪��'�F�%����=�Dc��D�}�uL�>�A�+y�LOUמh�*b�������6?=a���=�����Dz�޽��C4�l�j(�2ڈ�A��j���^S�HG헡 ���Ք��ׇp��P���=y�V7�se�����.�/�
�:�r�-t����6z��A�=T�ǚ<+�+�
e��;�E��V��qE<�⥸���B����h�eM ��"@G/��rAt��T����A�N�p�nn�*���[����`|Z�~<���3�Z@�]��x����+���ۻپ��h`T����5gFD}[	�J� Y,��3q�1���Ģ\����9(�U�͏��Z�Dı!��.z��ooui��X}*M-ѡ�Y5�8j�"G�r����K�C�NkЈ�k�CMo�W��O&.�*8_;9ZM��)�|j��l��.d� �%�L������z�gƘ*�1�)�����%���4o��a*]���s�
�!�N�85��L�j�3�K�F̩+W0,_ϴŘf�iF�h�JI��Z"�����[XI$k��<BT�?�b�(�:s����	���6"��L7�5;��'dsrV�\JϢ?�N�?� }B�D�_��A���*�5E�ƨNOE�[R��@٦YV?EC�/El��F�m�?+Խqζ(���yQJ�u˔��eY6��薰:#�0dDF�%6���H�Ɍ׆���3�ʸL� ƥ;����(�[�KO�0KI���r�(���~�'ф0���-3 ��y�&�:?u��	z��j�(:5/�9�N�QM�h�i~�<�}��)���0���]�����U3ܹ���c�v��w��-7VM�
:�b�O��&jB<�^؜s���w�����BJ/-|���D'�HAv9�φy��U"�v5��]��7���Eb+Qm�.GG����w���?w �݇M�冄3�7�6�N�Z0F;�<ѩ�LZ�������z���a�
$*�8��ؙ�n#�l5M�К4����;s�߫^(e���0��]��h��L�(���I�~�K	q]:���
yQK�=�NyV7O5��= ��"���]�?7a:C�qT�/PZa_<��JN�/rj*��%|٩�e�^�>_ �B��}εiI��z�D�8���K=b4I�y�+��h���G�hf�b�]#d͹z�	EM��P����2�'�T�ͪw������d�#�T�e�xD��]�Oߜ�A��&����K�9�ϛ�+�'�U[D�ʻ��d'TE��l?�4�5������8)���y���Ѕ�dkS�n�cR���]U�Qx���Oן��2=�6.��HM�b �E�^a>^�(؇����X���ȕ�����`2e�R1!L���?�:8~��3vxCY�t{���m���}�զ��^Db	��=I�V-ݢ�g`�o���DL��J�p�Yq�W`$�Y�"��F�`Jn�Ղ��e�Ջ���*�1@yϢ���ª��%����m�Wԡ�:�A����
�����|����{�>W/��g�>�y@�b����	r����	��//T�����0/�"N�g�����_�T���^{ �?����5�
f�7����b�l%��ZM� ��6�uU�Yu�B?匕/�Vp���&�&a����B��%���X2﷟�����>���8ܞ-QǤn���|1��ɯ[����³~��[��2w��.� ��4��^��� f,ޤ�A<ڄ%�,�o��B������$kG������(�Z{��B�����ດǫi#�\r��8]��_�ˎ\[�!�
h�:N�z������7R;|O���gex�����?m��tB6�8����ݯT`�l)��G��Eҭ5���d��~���*c|Pj�E*Җ��-$���S��2W\U��hj׫� ��h��Pb)�Q[ � ;Ģe����X��N�eKN��T�a�]0U��i����ye�K	%Y�쯾4�6��*�ʘ����&gەF�G�&(�?t���� ��)٧��1��,K��36��g���[�s����Fʾמ	y����Sb[���K����u��w-L�=";�wTx��$��Ek[��b=4bA���u9�L��!���z9x��F������U7C"�53q�X'U���L�g�N���p��5fǯQ�J��B{@�B��=EN����G.�0��7U�E����o���w#N��$�*����B��X��U>���^"�]����	�!UV�K��������' �!�m[��Y2 ��������M&+Ŷ϶\ս n��\s��z�7iO7���h�LnwTL�������Վw�UH���$i���hD�~�ú^�ٛڼ�pZ�qY�ۂ�Ҁ�����ON+$ ��XG�	�2�5,���޷�`���*��zsA�?S�S+�l�E�
?�F�8�c�~ׯ���4^jܬЙ�/U~�V���)�@zqu6Qw�Y�l�̴i�&v�@��S�R�����j�j)Z����z��V��u�ȸD��N��.Ҧi�&�YJ��!(���Wy�X�e�?���P������k8����1���{b��X_m���ãn�EC������mikDTXω�+�	6�"}9��?��'�B��D��z�����R�_Ed8��'�����Y�Y9PsMf1�1��m=	�l�N_�@��T��s�9�d�r@n�����4�)��G��tP�{�g�o"��4_���f�b���J�W�}zP>IH�b��f�'��F�:N�?�.������ȸ�rl0���6פe����e`O��fN.9���gŪ|�>$u�u�4V���]y�އ� �羯ai9#�>���"����l�͡�{�+���[u��\����ET	qt�"����ʣXqִ�����?�+W���~���-Y�4ʜ�̛�Q9�,f r���o���}��^��vړ��/����=F�թwu�V�Yģ��g�
+@^J�K����P1����<��	���y.�۾i�s�S�C>��k�f�:�y�K]�Y}�l�T��K�hr+JYG�nLQ'6U� ��|Z���z��J~����θ��]��<��]��6 ������[)�R��UmPi���\k~^)���I��"I�F�#_���lu�L�;]	NX�Mg&�	ۃ�^yvB|O�g��I�]��x=>�B'�� ��g��go�xo�Ҳ���h� ���#�0oN�J�_Py4e۴�
�[�Y�pOU���>���5y��l��|��:�Ad��U����B*tǧ� 3	C!6%�Zk�f��D���)_���1#��l@��x��b2Ͼ*(����i�A����������q�q�ߑ������lwa���������d4:�M܆�\�*�Zo'^�/)a9}Ur����Q�6OM�9��������}K$?���l�6(ɠf�V�)+�T���S�f�z���)��5�`1]�K/mMh$F�È$�f��+��f����O �3��#�.��V�2�_��¢N�]��a��ф'�X�Yb,(��.�m M�'9n��;�|_d�~����=�T`���p�1��}ĢB~.�7Ԃ7�[^�|,��P��`�si;q5�0+gNƎ�]���:�e"��2���c�����Wl��@��b��s;�c�ރ�euH;�}5싙�ՈA�?��;���O�-T
MU��6��� �j;���mP�T���D�8���>�K��5	��b����e������B���m&��M��9/��\�ZT�,W��c�p��B��ޏ&���i�n182F�u�8�S��?^z�7v-+�7xg�	�5%w�]?Zh�5E�.�L	���pH�8��iG6ˊ�Õ,�zH���-�Pڣ�;�*�W�G[��W�d��A6��`�-��摮m��$�Ǌ��:���Ĭ����<碇�c~�0��y�<İ�| ZQ_�i�8���{��e�;V�-I��R�!T�Z���G��lￛG��O^��&��P۽.��5�[���C �����1�X���C��4CT�y��'��%~�Y���[u
��N���"3<A��K�7s�e�Ƒm��s���*Y걉Cb�)�h�&��#�bJkE_���9����%��da4~�'��e1!A�a���
oB�H������i�	 ;���*����2����Κ���(���jD�F'0�b�~��@�;�+��[�kf]jd���z�Wa*M��\��Ϊ� �u��N�"���X!S{�%�LNg� �h�s�W�BMO�@z�^l7<�*T�ؑy<S/�,	iO����Q�^�DN����*9!O�L!�֑��u2���T]�"��P>9�^�'6g�<i����<��x�4�ƙ���~d{&%�5QxX����A��=q��r1K�p#+]��צ�T\�����n=��1$W����o��2��
`Ѵ�Ċl2́��A��SO��c���3� ��
=�/}d�;"�|��(�������w`H����N��29�I$^ʦc|1����5�U)>w|\.6N�~�C�4�����W7T$�;�{���wѭ��?$֤W+�C�9[���c��K]ǂy:�V��
��3@D0��DUn�9l<x��Ce�ס�ہ��f��*d�!:�������%��s������	�qDK��Yu߇T��+#.|[z��a�.)�]��(��N�L�Y{�Zh!�w��pÎ������]�u����̏���O�,�l��G��&/�J�G�3�H? � ����������Y%�pюuӇ�����?]]nC�\J��_5��3Y��R�����W\q�q��r\KM���0PTг�3*�C%�Q�"����lr����h��Mxf����4�
�=J�7�m�Z��i?�eh.��v ��]j���+V˵�ʌ��[#�$�ؠ��"Ji�vim�%n�1CvKY5^6>���ʧ���C�p��j��@%c�yD�di�a�5�w�-7M]�6ޅ�Z�����^�����p$b1��i�q�~���MV��0�bhAG,'q�h���(o9Z-��Vs��g��*��)#��%R']�R�	R$��_��%!�x���vb,�i�b��`x�>��V��<���@Ʉ���$��B^��|��2���%�W*3tKKQ�'=��1L��EEy�6<�_�4|�I��T�dq��pM)�do���ʑG\�2p�>5�nS��;T���)��S6k���lg1���Z0��
�0i�ۀ�{��'�)h��|�q��l�A����('��%	X��nH�"z\��R��M �������M���SsYJ����kl��ܨM����Mն�3 ��E4�o�c]����!;����<�ڡv'y
$��%���ϵ���}痗�nn0Y*1,�E���z�'���,$Ƌ�&���Л6���;��;ڬ��6?�� �W��`vp�3�T=ß�<�������s�%��sc��a�Uf�u���;�#�q�XK��FM(�\ENh���_k_�R�%�?�{�PK^l`G��K=%.��� �����Ԭ�{ȣuZZ���`��%����+��_�4��Wt�_M����l)D2�!0z[���?P�yT�������MQ}�p��3q�c�$�#jfhf�W��~�?�B�m8�J������tcǡ�:@�+�t-����5YVP�z��"��AG[��z=��w��D���SĘ��{�7JMscE`K��z҈)���pXI%�/�9�Un��+A� Ets�AQ�Z�l�.���,�ۮ�p�o�򺂇��q7,��"�����{B4)�-�;4n-đ[׷Z�x��c�WT}r�ʐC�#����Dt���fLt#��렻v�a'����8ge�ڪ%ͨ&( �4�O\��Z7�v���긁d]��a������%#��XzR1��v���D�5��|D6��XĞ�e�y1$� D��u:M3�!]����a4����S��g��SLuƄ��������u�����+j�����|`a��uv:=﷛�0��u"E��kc|�����xVl�*�a����4w3���b6�hd4 \<}!n#��	1>4zw�����![�Q�0E�	�� �`S&!ɣ1���H[�5��RF���e����Wd��6]������FotD7��~�O�# b�¦bc�����x1Nq�w- P��o�F'�/���h�Z�3vF��.K�?c�7'�X6����ӏʄ%����u��h��������,GV�w�
�nx*�[�袍rtA����Y��.�.q�z�1��k-[lg0��,v�Lh�.XVER\���a7�P�Ul�je��Q���.^F
��W 4p;��/pU(�kSa��%����}(Eu,0�'���8&I�6P�f���A�5o��B����A ���[��¥͒���T��UnN�X�;���U�OC[B=�f*;��f���'0{
'��$�W��U�C���� ��n�K��g��vo��>�pS|������W&��k ����	�,�G����?f� {�2s+��L�w������0�+8���(z V�����>�b���  j�r�⓳�\F��n������%�`כ��(��2��u�2
��5��oS��.�ձny�I�ŨT�C�/o�Vpmfdχ�R�eA��'���Cۯ��1�/
R-)(�[[���$��~x��*a��Ӿ���N�H�=zT�]q>%6�3�X�:�I$�-
-.*��U(�G��Xp�����u��&A�� �3�3
��K9��.�Ϯ�!�����ݚ������*���Ф����H��۷v��$�4�#��i�{�~9S��-u%�Ǳ�\iSJ�@�����Uq12�. Q�J~���e+�������l�3Ί�u(�w©���De
YJR�H>�.��Л�ۢy �4>��UoT�T!��ޒq:��?�w��?��)�󰿼�a�(AUtҎ=�|��Q;��A��kr�F{�^�-C|�xI�_D�)P`^����5{���~Gqyx������h������L8y��$8��+{�ՊE�6��������C(1�~���h�\��Z�9(�1��B��8�}8H����ߝ��0���C}��uK(Wˀ��Z��m���꽚���j�؂!�N�ޢ���F��#4l��%���&a���+"dD���r�^�m��%����q�7�\�$_f��^b��u�ߔ�_J�$Om@ʙ4`�H�&����w{�͍��\t������gjo�
|H4��q� L���H�'����-�����sΊC|
�E���0�oϺ���( w�F+P��Ư��&1f"��DS�H5�qk7DSI����5#���gw���>S���}�G�Œ��RڧK��.�G�z��&����S�bZH��,ں"î $)�]m(C���7��Dzuk��E?�z�RI%�����Am����Zc�%vJA��n�C��.��Gq�,����*�è-�v�ֶ��j�3�q�Z,qT�h�{�R~C ����U��p�50�u��s*�_Y�Z1��_�S�>���y�}�dO�1j&�)��f4y�����|ʛ��#�vܺPǒ���-=�L�h��I�������RT��m۠��|�5S�����zZ7��s�NJ8��"K ���w��(��YuH����E��K�^U��D+�_�C0���*]�";c���N���Z�e΃^Nq�8 ������g>!j��@�n�i��b���")��Ć��r
��ꓚ�p���9��"m@�o4)���Ec��F�?��݉����\g��{�X��{�>�1����C��6��u�x�{�A�S!�� �Ɔh�L��9O��$���I ��2��^/��Wq��ZD�,|~ٝ��"�z��	)����/�*�1���S�/�Bt<-�`�Si��x����ߥ0"{1�R��c�e��f�A¨H�C����E��ť85�[��C�����b�8�m3�&���/��N��5(����1��g������ %�Ee���>X���B�0�����U��G����a;�x�Я�x�B����@)�	�K�>�d��9u��*��=�u���#6�j��|[�]�ix"D:WdO|�3��<�i��-)wtv����2�o���
�'��?�/*���jhWIP3��N�S��;P;�xJW��.�/�jI�u�Rw3����%��{��t�)��C�U���C/@BP�Omj(��E��;�����)rbˈ~�Sk��luOW�i���C����2�M����z�ݐz������s,��(�PK\���ޅ��F��j3MlQ{@����F��ɯ�)�U���+��u�w�OH�p]��%Q;oH��*p���x���R�ϯ5��J���T:?��_bm��iN�W(7�3iY*ۊX8�9�8x��z6�^��F��摑!'�'�,�(񘍤z&���o񱃷S$_��{��D�[N���2i��9cV��}��gl�Y���'Л�dm$�l,��{r�4�Ȏ�+
H.�6�Y��`��h�B݃&=��?\�ǬMT�����K�H����w<�CQIˡ<�N�ۿ�A�\��H,/@�	��UZ��L�H4Ұ�P��Nc�
d�V��1x��h���K���a�uȵ)/t*5	�P1�ʊ��� ��,Ul�M��v���ք~J�Ê�T��6D�k|����r3���5�oaL����~��D]i,ca+&��&C;� �f�c�༙
m�&G$_v<��)�e����5G���G�%�W+�oY�N���ً�&sb��5��y��t`�|��A��ܘ�,oy��:Vv�m
<�@��{E��U9:]4c����;xv�5o�P�B��z�?��:i���F�_�vo����_�i�kE�mFs1 g�kB~�U��}����Y%��<
��b>F
���ك��ZIN��]ח�o���jUQ� ���x{Cɕ�)�1U�3���C��z��<�#��
�����NK�>X��W�Pk\-*1�|}����4�����L��G�����S^<��¡��N@��b-����D���wn��)qFˣ)h����!�u�,�Ӟ�x�w�S�cṯ�?z};�hbSK���5���ŨYq �(8��>#>;R��B5m]�z9����Jj��к,��J��,"��9ŒK|���b���æ�Q^S���?�d��bZ��D���͝���=YJ�D�q
YE�w���l�l��h�[��5�n��X���p��6�H\dB��vpXKFJpZ f$j�,�Ϳ������H�DBa-%`�8��uv����Q��*��?�T�F�|D��;��8eh�&{�r5�8�A�=d��m O��炠u�OG��{��3K�{��w�nR���?���r�H̖0t�<�)�&Ȑ@�"��H�)<C|�o�<68�2PP�|36�2&bz2�<�l,;�4�kv�Ng����!�k�@P��F~!���M���Dc$�讀�e���3��W�d�^��V�����Q���}=�rl3�?bLVzh��(��+?-s�vU3�b9 x�MF�Nج�x��mʡWYK0|u�i�[��w�{d��d5k3Be{�[�QL!f4��-rbD?�$���K�t,�n_�Fr��rt��a�^��G74$ߢg�@t�ػ�ހ��y����7X��(KS�"��T5%�vnjp�)��r����d��?��i|�`�%3ԫ���gc$���\F�?�
)����ݩԊ�m�N���.7��sg�R�2�>sK��{���f8L����~K�(���/^ޟG���VH`�)�a�vK"޸��Q<�9,Ƹ��?]WZ=z�FvZ��u���_� HB'��6c��s�P}�`�j)��ac��DU��`%���:�6�͞�+��z�����J������B���N�$���;�2ē}���N�u����Γ�2ɈLlRZs���N�]ovW���}b�V(��\��P
�+�
a9{>�fY��b$'ܯ�~Q��u)�ٚ��ذ�~���M@U�(O��fdcPr
���>O�����n':f+S��oD�NO��1�(Q/�NGҌ������fWÒ�x�>/�rj�+}�9 �]O�x\�\�����@d�FuI���Uun�i�)S"l%gHO9���b�T/��)y jx�I;����ݨ��
Ϟq�j7t�I�x�`�	
p�߇��=&��<����6�ɭ�3׸�jěY���;m�=����jx����K�^y��]�̘��R�u����_х +%=�yGR�?^� B�����3�Ә+>7�h+�"1�J�L͊{�Z؃����<=�G�A.2���66,��J�7,F5
?���	�C���B���$���l��Y�
Q[�߃��Q&��:gP�B�18#�z���F�C���̣͕���v	[k$�\aV���T �]ُ�x�+:-R�tL�n�#Z��h�o+�bKi6�L=?�&��GPO������3��c}"ȵfV�0�HR� ��*۟�� t��پV��fU*��`�/|1�2�_���"��d1�a%A#��ŋ8����f���	8���ֆ�зX��P���aQOW�m��Xq%�|ƻο/s�y7q:���f~ͬ��0��iJ���'���ӽ�&[P�7d��c^H�#X8���E�s�嬡�����)��T�d�yYw�w �b�\�<1Z�t�i��>A���=�� l�$H/��g��N������-���ŕË�P�g�9 ��.� ��8��)e���8#�5X%Ͽ�Q��-��l�	�4���)�dR��md�a"�Qk>v��O ��7�#C.l��z`����g��,���@T}�1�����a+uz �cU�s�v^4�yI9�h�Ӎ���)��B��7�dK.7�֩nW� �.���{<Q=�϶�J� ��HB�{�l�_���v�r��)��y ��
�:��)���״`:��h�cj��b��І�3�<]
�O�r��y,(�� Y��<Q޲�ɚ�/8�N�b&�c���k�הA��,c��֋�u�Ӯ�->$)��n�=�v�,�4���B0���C��?6M�K�a����>�����^�OpM��FH³�7���Q���W2T�&۹�<���G7�$���r(�*@N�a�<O2䶨[���v��'�������QI%jNɊ8?���&v�|`�7fO��jt��4րy�C�	˂r����;�}��dM��ȇ5X��C�.u����Ȱv��b]G�?���U�³7yd7z��^�$�U���23��sHPp��s@ڲ�4�56r�9~	8��q&H�F��v��G�щ	���cґ.���3������拞dE�8UOnH{�||�Y�zw^]УA�	�����/yIW��N���{12|z���K���*�S��}�Gy>GV����;�^	 �  �!B��4��N~J5�����&�^r��a��MW�Ȕ��N� AgC�Ԃc'7�y�\��[@
�C��Ζ��A�.�v���+�d�y}�L2�O̱^?�"0>�B8��]�\�A��d�G���u|N�m�A���ϊcu11Y�>��D�ɭ +�����U�̯�ؚ��J$|x���	{��� �0�� Wn��(M��p��p�����^��^̲8���kc]�X��U`U�o]i^sW�P�����(/g�f��u��
�����rmӅ��崪� ���G�s3B�N3G�%�M\}+���}S� `�J�[���h���J��Sܖ���<�,*v�| ���kA�/�g����$I�n��B�x�L�'L��W`������	#�u�Ƴ�m�.�J�-�B���������p��-�Ȇr�t�?��,rc��J���]�d� �͘G�����B�LGG�焨�&@A�: l���?J�ջFf�L�፹�&�(��KA�^�S<�U���)��m���t��ƾ�����B�R#�(-u��dA�ȩ:}<9�[39�O�7�T���fA(�g�6
�P"��b���Hy��σ	pkF��oZN�]G�\��C�o`|D�Ļ��͇r`!�@ 45��s,Ҁh��1�E�(�^=d(��Ɓ�����:Vf0�o����5O��[�����߹�U�+xJ���yv��\���<��1��"S��H��2)��R��E�7e�45�a��vT�/՛� ��ν�$�]��:
�f�X��:	#	 *����D\�n�O���xZ�<U,�pX]P>��7e�;w��<��C������@�j�&��mf֨��7.Bt�ה}���3�ot�񶎄�<�Fl>��T3�b���m��P�+`�g��ҿE"�+ Et������'����H������vX$��6��h�پ��jI���|����t:g%�uF�*�}�I|W��k��df鮚Lejn�C�>բ�dռ��i������D����*�\J+�Ƣw�J@�=�g�+W�s�H�A����]��s�~�̍�΄��L�V���	�	F�ZF��b���P��>&yf�Ǜ��i����hZ;��B֋�ͼ�ܕ��|��jtd��r�$����e�V�V�����p�`[� �|��:3���k�İ���m�癪e�U�d坒#��\�?���tG}���NhCj���U��[AS�j,����Cˡ��s�V�Urt��Yߓ|I�����-�t~�L�d�o^�c��+�ϣ���/��<b=^�t�������ю�A��NN���Ѕ%a ;�	�Tf)I��|�!�%f�`J�*'����Hݦf�FZ�,e��d|�dG�,(��|φҜ��3 hv]@��h�+(5&����Q��Z s�&4����@����c\G�C��.ʂ��!���Չ�OB��.<Ӝ2"��N����OV��oYCz��/Y;كl`uI I�����b�8u����k�
|t;��Y!ٙ�)GOv�w�QD��HK��(d��a�/6"S��*�_�_��]-��5�V��;�=y����!��
��#�-�6n���Mړ�T�-����`��tс��{��p3J<�hl�H3���Ԣ�y��G��ba�^�`�L�d /��~�2��N�qH|W@.IG��^���\Q6?)�+,���C*���M�\��R�� ,��|�x#a�@�%+#�l��F�=\�.��w,%䭓&�0��\B���S��E��H��)������i�s(��/.��ΰ�{냷l�4����<X^[�K�R ���C��"��5����7Q��;̓1A��Zݷ�=�,2��Me��qc(R��ֹ�̨���/'�n ��<���M��B�p����{�u�����4�4���]��)»(G�`WީȔ:3ڄo^t9��
�
O��;���u�T�Pu�����t���N�J<G�"	1a�F<e,;5��=�����R�.��ۺ�7�7]`�`�����a�
A�����J��'��]ZnI��Ƥ��m���^�gǙ߶5���_C��oW`��V�M:Rtc�R7�N\��ݡ���+�㨤U�<����� �U��$V��>�������B)%K�te���~�~�tOC�c��p�W�!��M�TrzH���ܚf$�LUcP���/ax�F�WH����i���4ȧb{�XG�B�b����hv��Ŭ��&��
v�T,�J���I>��n9�xT�_���e_���Ru�6���@�A��	R�u����X؜gy-$���>��:��l�]�V�jqFe��:�B��,~�_BFٴ|Q�a��`�h�̙���M�����*�d�x��\|�"�t��?O�K�����]�;.E1�Tjd�z�Dp`����#`)��G�g_��Ki���bh���F��*���ua���{4�c����h��U����4��E4�	r+j޵U������eD+��K����w�kv��uֻ!�~����P��*��!� ��IY�~�G=8��)�hƍ�FpP*�:;ĵQpI���.�M����Ҁ�aC��&#Ҹ�����`;��j�����Y���J�� M*��Eb��:��G'��{lWsq����n�P-�v�)�7�i�葵�1	O�%��sEpv��0ϓ�A���˅�> u��6c��*m��h���o���,�j�Q��Qv��P� �{~Bv�Ivƙ����;�o���;=�0�\�/�y����{�����zA�1�G����'\(B�C~��}�܅��'
��͔����Ł�?�yٶ�\}.	��(�''�]��`5�i6NP�鮘@D��4$�Dy���:�Iq�x�<�dN��Y��z�0�d�6H��=�a�FแE�S)����k�m���erU��]�j�p$���|�H�� T�&� ���s✅f�~mQ��ԙv.;zzݞp��P֣d�+�P���4��Ɔ�L3��>`�0Z��xfժQ���t��C0<9��}�d*[��}�©j@�'���o�DO�ނ�������E�3��v�J~��<őr!<=CW�S��\tU�"��5OQ&��of�ǟߪ;9��ȿ�/G��i�ە���K�[��E��/�7��c8H���h��c�嘏� �#We'�>�-p�Qb�����uCJ�%�4�S����w�Xż���a��q�2&�[�7��kٕu&m�2b4��o�(�]�,��V�F�g�L��!�,b1�W�>C�&B�/��>��u$Ѷh`����=�B3�L�G,`����V�������l�y��fj;-?��;���)X��|q�֒�,[g�@��2h�=��r�{��Zqsr�(�`��Nz�h8G�{я�&��Y^^��m����+w�d����i��a(���`� ��
0a���RO����^2lxDȔcNK�Kb�E�l�y�lo�`N%�K��J͗3��
���j1HPK��=}Ŀ������?�˹���Z�c.P�.'�2/͕U��P�mXq��r+�<�na[�pkt��D�`	����wR�Y�⍂���j�Kd6��u}��f�/��s�v�u�r)��AJ�����-�3r� ���hѪ\���7cQ�	&�%����p�R�b���\�2�mx�*/���uwKf`�O��*Ip�ȭ��`%t5��F�S;L���E�J�m�,؈���F�hy���Ef����낽�뷜�R���Lu�JP�,'m��K���8DY��&���]��i��|��!�]�K���L��Rq�V<R�+�<�~�g�8KxR�&������:ۜ^7S�>j��l�'���P� ��_�M4
6����"$�(y�s��H����o۷�?�x���VgE0@���N,m_x�%)8�ǆ� q�m2,ۮx������9���uEP�"��z�j?��sڌ���I�f�I�~�.i*Y��,p�v�qAJ��rb8�$�#��¥`'?q�Y)��(&F��r,�����!K� �?ԧ4��e?�r�>(a�{[��e�@$T���G�:x��+й�u��k�/��ᐿՖ`�h� �<�l�8G�c�Z*}�M�\�"�c)���:)�!�ßwH?�Q�L����E�Z3de;�����2�,,�����K�����i�q��w労��`�uT�����T��L�g����&�W4�@��鯍�on���*�Y|�B�D�4�͟�Dt�R��5|�Ԟ�oB<�yz��:ƃ`��y����4�G`�Ps���L�|o?�,������f�"j��XX�g}��I�dS�������}�h�\p����4��xe>,�HہFᕒ_���xS��X�𒶨Gp�jaz?W�%����J�����k�7�b�JϷ*�Q_ٯ�n`�deK�D��p�Z ~��$h�h��T^����7�h� ��R�.�*�v�P[�Kя�%:��q�hKW�rHU�䐧a�tIY�]����� �K��"�s|\`�|H� @��Tr�@��q'$���ƣ�L!�~��W�QߓP�쐫63/l,rF��2�����Z�>�<?-�ne&�N��6�An����;�����7�������K��>Y��®��ǌ��c���.Fؒ"Z�</���(�)���ObN�Yƫ$�Z�fT'-��Q|�2
������&�F��;c$�b'���\�9����S:�)��-v���.��Ht��]������,�4.~��ą�_Z�ҿ�`�L�S89?�O.%3$Rj��"�iމ� c(`�<�Cݵ��ɐˇ���ڣ���.X�{ r�6�y�P2�$K0W&]Dc�L�N��M�xZf���CӃ�]�P��K5틲���M*i7ݽ���N�x���ʚn�o�Nѓ�:�����cbʤ_��B�m~%Y&�_���G>8�}��(�a_-����1�jڄd�b�"*e�h`�J��,{�r%9��,�~klM����$�[�ض&�:�u��F@>4/���t���^>�."�^aZ�+�2~B.wY�U�=�Ps
(l[r[o$>�z�^�����`�sW*&��FQ%�Qj̗"�C��Q���b������`{�iqyVs�0^E��\����Z�4!GpSMxW�eA��r���_p��i��#�"��x_�3�ljk�p�t��o|lgv�	�)��~U���h]A1�����'��S.�I�_���g8Q�v'g^Q����>K|s�zV9�
��Q1���*�]���}��Ԑ��3jO]\#�HA�x<�@�d3<c��ĺu;��)����G�����<��U���KZgU��mp���H�K����%�0��Zg���Y�d�J��d�"�����0d�^�C����ʋ5y}s�P�sqN��S�G����|V���9��R�{Q?���S�6�W�^�Ч����0�Wc�.Bq#��I��9rU��,�f�i���:����3v�JP�G7���*��m�!e�8DJ�lA�I9i�=Vc;7�Tz_	[��k��P�OϠ�SZo)\>���?J��?hܼ&6�ȴv�8���Z�Z�����@�#��5�0o�~�(�����Izȫ!8ȩǸ��
WR9A�ZS�P���8c�P���� E��a�z׾��p|�/���+�?(Ҁ�QHM����s�H0W�{�p��#����Hvf�K��Y�]�얜q*2zz�Uⵖ�U��s�O�͎+�,��{��*��V|>SY����'�o3��>�Y(4��#FZ4l�o@'�j�b?^�(齌��z���+"w�j�*c�r��r�%焠os�W �bH��E9�	�k��l	%%W�j���h�$u�PFz���t����;�Q����QY�ڄLu��1�|� �{����ɢ2{F��R�J�tu���v��uJ�	�^�������4�f�$�'\;��7��i�u���T�t��R���� �㺵��򘕆�'s�9�����W�>�V��4�8&�#��F���MW�wk;@�A��J��	��F��M"pwZy��)@���e*�P��9�5�O�e�27��xq��Њ�S�(<��#�ܪ�Vs}:��8Lg��yEMU+!�ĄFJR\\��0؄ܖ�^)E&��21i-y��'���}�7]�W8�Z_�05����g��&�!m�	)�j~3A�ޚ�E�WÚ�-��h�3���ʇ��Ò�i�������ݖ{��ɍ�\�U'�i��=z=O��q�ʟ���'Yf�Pd��ɚ�HT�������-�f�0Z^��BDǡ*�e���-����U�]� '��T�h�}�q�7���L�� V.r@����؝�{��Z�V{�)E߭A�������пT����[��\P�[�7`�df�9�Rp�[B�b�s��s{�?|�qv��p	L������:]��	:,�&��O��&��&_@q���vY�/ٛ��{?�4TY�F����+�P��8�*ch�C����fE���zZ�������<a�_" I�
w`�������	G� &bo,�Z�:jwHrX� gh3M㕍$\FrM�#�U�s����O��+�Z�J�ۘ�t>�Lx�Qs{+>؅ҵ�N�IּBi�`���wA��TT��@��z;
��1!Y��=8�V8���w�;z�ܕ0a^0?��~	�-�Y2���D�R��cܙ�������u�M�Bg���J�tUø� O�?\p���#��#�.���� L7�����]s� �4#��(sf6x1k!x�cg�04q'ǫA52^h.)�O����J�Y�	���r��������T@s�J��hT~:���e>R
� �0�P�I���b��,�Xؠ����Q��mi�T��=R����v"mg���o�# ������Yb6m�J�a��1?u:�J�g�_?�ʘ�o��ܙ���10ak8��#�����ܴ��ݏ\�=}su�c�b򟵈�3|�6�:��*�q��ַ��P.J�ٿP��L�>C���Uڕ���ǯY#�7�j0�6{����XQB�]?��C�6q*�b!�Xu�i�^�xx7!�@1)޴%7Ѹ����
�9��dd%N���'�Wb�7uI��l��A>��J�_�>Ƀ�\Y�pf5'����֗&W%#��yӯ'vԪ˞��Č;�p���*�����o�䟠
Ϊ�a@�W�tW�He�dv�]�޽�I�d��'mmf���X|�G.��c�(�!�1J٠"?����4?`z[ϼ�Z�.qF�����)��-�H!b�Z*��6Nf B.ؐTb��0x��)��/5���7�zG�ox��u5� ����ӨP��+���v�^U"8+Zt֮�ɶA�2���"�V3�U��Z�ie�Z�]���;~�mwU�HHz��4	{mI�P�-t5Du��@��U��ө�G�T�A�Z�_�*q��LROڈT�}\��Y��&	�h0o���e�i���]��w���.���ug��ѡ�~3P������z�&τ��N`�u�[֥���Y6]oG�0bŖ����(P���Q��ё�0�=�	�s���"sؕ�k&R�/�=!$������tr�������k,���:Y�S�U��-�K_��WnY*��P�����A//PC�/ G����-���ڛ������\P�5o;�x�ݸ��,�r.��@�T���-�f�3�DK{2��,ܯ呑\���;�z^KV�,���G���>����L8:��/`Ƥ�.���)��~fZ� 1y�ܹ�cw-3a^��K�2̋o2Fd9a�Y�@E�y4��8͝'��	�)��2�ҏ��2��X��Q�4��Tk}T�uY��%�A6����K)���y/�P�(W`��J�	*k�Il�uȻf���ԺsV��
�o>���ҷ���W�"O&>kυ���p���j���yуP���#\d&�efM��Z��>�z-۔ln#s�Ez<�iN��R����U�j�P6o��ӳ}YX��Q�,q2��N�r	�S��C�F�R&�p�<���GE����\��b���;�ޔ�M����Rt��>��0�+Si
x7�V*�-$�i�k��%آ�N�*ڽ��K�>����-�#�T��&ź��TQ%���ƽ�%[k����O	�=�Uq�YJ�%�-����9�	�����?�V�T`N7�)T�B��V���W�Ui��B3Pr�(<���7C�N�-
C(_,�W����D�)�I�_��PT�����!�ج�b
�h~=�5��Z�3W�����Y�>�gS�"�����.g��Ix�ԅ#�5�u�
��Z+ �/������c��G�j���ѵ���]�� �G��Y��<Z�F�`�I��]ʎN�5�|��9Iz�k%�H{� �@��s�~�ޑ
Ý�7/�3��%�KV�X�x�E�0-$<g�k�]z��E�� 髐�{g.�c9�I�1CL�����̽p�=1��z`�ݕ`������R��C����2��O�5����f�A\�j��_F���N¢�)Z`�D��c3w,�Mv�m����FP�r����#��5�	4W��y�*���RR%�Ӷ1�)�XKjŸܗpQ��M�0\�X���a)�`���雇�=Լ������#F� �ǯc(��5��p���b�^�s���dOH-�E|$�l�f����"��][+��A4B.���1a����%�d^�w~V�=�qs!1�8a��I,� �c.�'�N�F"ځȱ��5]��w�)v�"F�]��!vyq/�6�9�^-�n;��ݧ3U��AO�|�J�Dq�X
�Eϳ��e0�����lZ����(�2Ki���U�
$���H E�-E^�v� d� ��J�+F�2J�E���+��qw ��G��=Y�j,-��Z��~�>��F��j&�l{h��`mz��7�m؂B	C�Y#Bw>}�h��;d0X��u����6x��L���ac��|C�]j�Eg5���
�.`J�x:pD�墄�D �R��փ��X0��7)�#c�Y��Jb�:	�^�3Qm�R�%nY�_�p.u�2�6Ü�hd�b̡��4܂F�p�?�|�����|$*ڬi��r�,6[�L�X!>;��r;4����,�DY�o��r�#z������Sر>,�!�cf����`6�}*�3�H��F�ps(����l=p|k���2d-@v��æ�%��%�]��Ad���9r7�?��%.$�����pC���z��N�&�7h��X�kЧƦ�|�@�K��+��־���7R��Xq˗�`g�eec+���un�8݉lT;�}`\M��F�J�*���F� cә��7���X�fw^wd�&���a��#T���m�-'S�._����J|�\ r�����9r�96�~�q�`9��Ǝ����E.��RE���<�H 	ky�UuyN� ��rf�IF�v�>�L,���5.�N��>6�|������W[$1Xc���M^���ei�i"s�G�x~��rXG\!Yk�b��^�(�U��r�U���"N�\ؿ���1w��z���3�5F�d~�B��p�W������t�'f���x�Y�w4�O���맶O*k��>�s�Q9�T���*��H~�I�����|���>P�dQmSk�G�c$;�T��Ź �A�Y�L4�Hk�����M��KsC�d�ڇ{.��4#���1^3_!��� zP���ٷj�@�{Z�c���=��ٔ(G�S����d�FTؓ/��;��x���5p鬓F�	��ڭ7�o숯VGҺ�aa|˪�y%"���(*�g`�ӆe�S��_­��OՓAS;�(�R���7dO2Ǖ_�,�8?���״�B}�dЇUY��k騅S���.�/?�oKڂ�J+�)�𙚓.���_:�6���d/�Z�B���T��\��L,���þh�8�V�����O����֊�4U7
���ɋD���LQ�i+��	�F(�~���J<�h�F�F׺"�������g�����ȪGr��#��.�*���1X��_�	��^�5����=���h&�S�)�#p(H�~�lnBvw�B�7�;-y�>�pc��s�)|�@C�Yy�>�䔲v��A�v���� 5f.�Q�Y�"���������qid�4�����ܨ��S���j�Js�HK�ʅ1˖,���"��1b<^����3er��nI� �l��'�.�EU
�W�̂�ש~�Cm�c���l9E��c�S%��G�YT��m��}@͇�S�9H�cZ���wߋ��W�L|���v���&q
FçL[Y��A��7;�z�я9S_��� ��}�#�L��Y��6�����N��u1'i47��wf��$`(�v=6A���&v��&�a [�[yt�r�Y�V�����	W�Bs�t� ��G�Na��RY����R�p�����y�t�{'�]���菩���Uf:s��b�	��bb�!9\����k�l�4	�B��?m$�Q�[j@꤇Lӎ^־�n&pJqe���Q�g�Cg����uJ3��*.J��X��!r��#~gF������ߍ_�@���,*1
����F��ZYM:;Ăb��{�ŵ���ʘ1���	�%&�H@J�W����@�]u����.�1nf�[�`��IG���1?6ү�?F�)���|1B��4��JO�i����QV<fەX�U��)���+m���.�XEirg]-�Ô�d�T��c@k8�?�)w�٧c������6�Z���5u���`7^g�LPKǾ"{>��[PlBw;�~��n"J}��wml�n��Ȅ{cw�󍜡� �e48�t{�ȖZ�M�4��O"�ԏ�n�%�I��s9fvúm�Ŕa��"�s�53�<Q��@]g7�����d�I!�pФ�h����u���C,�����jHh��j(�f*0��,ou0�Py� 
��Ȫ��i�P�)u����I��rYvc�r���B/��ŏ"��e�]�ABfZ��ܕ��":�Fv)Bܢ�%�@#�ĳ��6s,W�i0�r�'t���K$�~ipG���Ъ���T�ch��2T����;)?�'���N���	�n����uǱ&�e�s�yF����0���R1�0o�m-�{0*�N\4
��	�un�D�z����0{���~&UӲ��9�ިL�c��;�����{���G<R�J���4Ф�������8�Ee��	Ф�.G������5��S~u��~�YZO�,�Hs)�֐w �&����j���H>�L)�x\5��-,JW�is6~ZT��('�_qr�v��ۑ,��Pp�{ϷHqL�)E��~��ܒ���|�m��z=���|��\g���[,9�L|ZA���X���C�'1'+��z�����pG�4�/��}�DHZ���J�/�n &�����<�F���}xI����T*zL��Q�~&UU3�D�WBq�Æ>���<�v��K{�ə'��C�mo}b,�\�l�����)	��xwk{^*�G�ߕ6ki���R���#C)}T�#g�	��u��g�I��l���K 7:������Y���Y�c77f�h�� y9��Z3���l��~8��A���ܫNВGnp_�2ݝK�f�����s��]~���4�����2�U]�d��GH)A�5D.�<���)<8F���uI���4����*��%��<��<G�ȷM����JV�S`��5K��q���7�atJ�{Dl����a,Q p��I���|џ�թ�6�.�myM�տ^�<�  p~��z��U�?��>~�w�;wx�f$b��jB��
�����b p�Gê���Xx�E�]��,�����֠���B����+���q ��MTkbCq�z�M�Չ�7"~�<�g�̫R��_(��X�_�N�%�26b���<�X�#p�v�aDUDO�<$=jc��c~[(����b��� �ֲ�� k�/��"���� �gh�������@}^Sh͐CV�(/��+%K�*�3L�ak��o]���V����)��*���#�~?gk�f�ձ��i�nZ�˱͂�|87���U�+V�N��<kU�|� �MK��(�=K"�o8Ӑ�S�������$�"�1u��%�Y~n�1�wYq���"�x���o�^�c�9��R���E�~��{~(#�T-���8֍<)�I��JxD�`#�^�aP��1ݓX�`T�ɺ�����q$j&ՂGQ���/����z�E��[Ia�>v8p���4ʸ�Q�%�#-d�9R�1��;jwJej`ĥ8Z"J�,O�ā��&����X�Ǐ
�ݳuK�XxμL��)݁Pg�q��CH������Xq�����c(vk`�j�:�"�>�B�)�A� Ņh���9�)��OX���N���A���"G>���
�i
 ��+�]A�6�욗�bIHV�Y�4 �K��ɘ<����X|q���V)�+T��4�o��B?~ v��%�d!Ya�/n0�a�u؁�L�WM��M7�X�2��i����ɟ����5�m������@W;t�:[+��>e��oN�7�Ks5�5>�'HHVv(Ϭc5:��S����b���m�>D6RV�W2�V��0E!��+�0��+Aqe�A�$1����?a�T�<�L-&��Y���O/ʴ�D(�a2���8/�*V�R��4�R�����E���i8�oj�4�����4���ώ��[R:���3C��j�A*�����I�V��_�A>�>Um��GmB�i�6�r����C�E�V �;��%�x����������,iM��]݅4A��w���ݑ^R�k��3u�,����X�l�y�i�f�p�*o
t)n��������9����A�lu�,�R�Qn,+��4
�5�,kt�"��TŨ� �����!4C�^����XX�U�_|6s��f��X~S��#x�<j9�"Oq�f�}ɝ�[nzG׭��r%�_sS�z6`R\|�*{�	em�3AIdsqk����Ҳ4�s��:�ۤ�G��.����&s��{��'
��'������79?،�egYK?�x�I�W�Rg�'8���P4Ř��X��5�����=�B�&����C����TK&I�X6	F�f�z�}�J2��z��Ü�>Z��kx��A���~���]p *W@
>jel��0������-�&��g�K�&j�i��w���S\��E�9y�Q;e	q=$(��@2H�}�A��X>�~�s�<��p�#�
W�[��x!�S��e�?���T�=�v���M |֜�]�Ym�1G���Y��D�cSw�ܫq����lV8)�H������&SybR����hIT��̀'�E�bSb辶�Ё��(U=�:��*�\P����)$Bd]���KVk�&T�hZR(�F�T�;Ǚ���ޔ��+l>'�J�K�X�����e���s$�Fi"5%�8��_�t�m_x�R�#�bu@�8�^K(K��#�[8�d��RBf\�]
�'ǰo.����&n1�X�̯�w��Y+h�7aX�A�]J펂mN�6��|�j� J�#S�Zl�G��}��Vx�qB�&ɴ�'WD�GZ�H�|�|S&�z�A�c���M�k���G����lΖx��_ΰk*�Y�dݗ
��~b(ؕ�ë4*9�\e���v�:�W�GIXL;ʒ�U�5N��u��l��)F�v��)^��wE��|�e�f�4:�q�A�gI\��k׷v
d!`qۃ�5o������@h�����*��&se%|�b����0 �/E�v��ֆ���D����б��d��u���3�z�
cC�/2�}���>q}Aho�r7x���T`E�4��Q�8]�N����炊����{#����r8�K��CGx䀱��Q���]l�7#���~�pq��\)��X�;���IӬg� R䒅U?]��g۔�ۈ;}A"ߖ�>;�� A��ri��A�I�jS�O�]����ۤfzD�2�b����t�`�OqOm�7�kj/Ա��EWfk�Nt$�d)�@�a����̪�%	d�Sd�?X$��$S7y<����t\��sy9��ķ�[��Y��~i$�Z'��p�=��W�g/��59=B�P9,Q���Ӭ����繽G��i�B�_��c%
���%,k�����O$���k����8yek寘��e�g?����nP'/��eǧQ\\e5�4������U���ډ��
;�։[g�0]_�k�m���c��4N��+Xhb���R�Jt1�/�?� �әf'���~�/�e�qs	$��t�5�4􎛲)������Fi�N��cӧ�� A�Iq+��Uw�Sb���Gf�
��p3��aq��[jJ�!���{<4ư߹a��9jں�!W�����5� ܔ��,��Y�������q����rv�������q�ȸ%�v�/�ے�ӆ�I$R��}�ɔ7��&'#��~� ����[TG�Ԭ<�[��V s?� r�#t�ZԎ(�D6gE\]�t7��U�$���M�l�[U�S/�pl���	��y���pX�\��$��-j1������7DFٲ^u�F���Nz��E���^�O����e-��]}7�/���~�+���ZrC;��n�ۨ��C�5Ca�s|��s���(i����B���Mv�r 3���"\�j�� ���R%ceu���p�S�́������ �)؛^4�Z��(F��!�S�&3"�.�8X}�F��I���[5|��9;2�x49�X��xRj��q�=ŉx����NC~wG$%�*g��/4 �Ȥ>��Q$D��q"V�b=�	���(�h�����M2��{x{�^(�������^����CB#�m
�#)�	�A���d!	��� ���L��@u���*���>��:
mEu?�נ����-�j:���K�F��������ê��GX�� �Joۊl���e��0tS`c8:�9K�d�6���6	��ʻ�v���h�]��{�+�)�I�b̔ťJf�ZS5�UO嬾Yw��j �UE�!;uV��5��^*t&�NR
']c� ���o�����a0Խ؀��?Tv7
Q�V��� ���w�e�k?�W��=���u���ۈT �SWW�����w��|Ӈl�A�-y۪�h�T�.4}(�؇H��������5�F
�����Q�D\]+'XJ�u���5_���o$�0'����p�	DD�}.d=�0i��L��7�] x[�?j{�D���oǅ���n'����i-���� \����2E�,�~]�8g�.ʧφ��U
�;e��X60n�/�XdSJ'I�%���f�ޑ%�m��s�F��8w�ʘ��?׶q����b�K��#���4g�:LQ%�<�.�$s��#�9Ο1l�=x�Y[Y�pcɾ�E����򿙎�٨"\��o��{��r��F6���b"��4�$���:�,V��d8��"�Q~G�^nMj�|E��齲쒃���Ɯ^�'>�]26Ў��,2}.��	{%c�@�j t׋�7p�Fvw����"��m�ѩ�[��*�vi�@Q�7��cd,A�K�s����k�:� f�k5�L��N�#i-\z=?��fY ��P�Po�+b�?���������jX"�2�B���[ ������8��6��b��/"�H�򆾡]4e;��Q���M4�rЄz��o.j&�}����?�x2���--mpm���s��E�fA��#�&�~�ٛZ�.��-j�#���q�u��eԞ/O��de�Y����1�Q'�5&���6��w�"x����M*�n�RaJ�S��՜�0��6G�&-��$dq+/+�E��b�~5��ȢT�4<������o�
>��,Ȭ/�Dx�f(���T	��'�ʬ{���߭b���������!�qi��r��{=g������t$�O$57@�k�7M}+�����~֣̎V)���g���Uy�����ϰ�e�em�'��LN�_�j�J���0�/�\�*�)X���хyfj�!����,!�6��@Ø5��Д�:=�Twn���db��x���Y+�u��0'�uy��1�R��
O�GMVs@�;^�_��ш�߽�*G��E�.vR*�T�K}5R���Ĝ�e�6��L��G��d�Z:���}�D"�7�b�:.𑄽w_��U܎'@� �*�*��vr����2MJߧZ%Ȑ����<Zy���p`Aՠc�fI��w���1�k!���:�����u�	�M�� ˝ԮG��:�/��>��TJP�x)��TKt�G��п!���>guP��-��Cǭ��ɰ���u�AA){��ۥ{������J�n7�P���a��%�$ª�I 
�}�Pa1adI���aHB���٫a�w
���(����,X2;$�v"����hG��(E����/2��#M0-sjZf��	��o������^��ٝ����>������X��x�CjH6�����6ܸ�^�~�a�b����?�������dq2�7O���$c��"�*����%�Y*����M�:]o�ݖ��_�wÄ���X(D���b����J�Z�9�;0�@
�&U�GU�]��}�����G���8�����J7S�5���D<��V9��oH#��{�Zl{�f�(ٶ�3f����6Y"�> ��RH�u��|�el:��8�R�����\YF����`6_J��h� �sE�c���tqS�4 �Y�_�Sx�qM`��ߍ�:�`Gt<�`��3��+��n�i��c=�����y��R3�6�}�e����@:�m��Ξ�x�B�Ȟv���&�V��j
������h"�Wڄ<���|(����X��us��&���������z�L��Up�hog���~K3��p���E]���0!1o�ŋ��KOTM������,}Fx9���)M�����:�����Ð`}�0`>7�����M(\I����MSI�	X|�q��'�p�d�5=����u��:���"�� 9�����n�=��N���{�y�ȕ�F����S�#$����>�ZB��j�u��"#�}�n�aJ�-b�cΨ'5c�1���8%�@�M��A>g���h/6TXVl.���[� Z	��!�����Y�f��Kľ)�cA���a�ɚM`�6h!�g8'�j�	������|c�.S�mX'<t6"gF������XJu}���Ѓ�6'��s\��\�K<�vP˧d1dh��'1?�_��5�O�c.3��YF}�j�U����Y�;�J}�A���H���S�!��-�r|��֏}��(�:U(�L&"]�ӎJ����!Fπi֏x㨈���k���*�Ky���]kr��qe�L�NY�����@?ʬI��V�}����$Д�^��b�)��>��g��Yr�c�q��fR�HAʹ	μ��sio8!�}���a�!�g4b�u8��s��Wܼ�Op��R����H~���Y���q�6#���hf�;޲��T���Ȍ 1M�*�9ܸM��-2��hZ�^��u �%ʓ�js�O<�*�x��u�  ��ž���x�
i�RL��DZ7�/.*�P��;E�xe�b�uj�!h;qI,G�_Bh�����T`=Q�`���̷Qa�X����%�;Mp��t�M�5Q?�;�@k19��B3V�E����U�l�t���0��Z��ӑ�O�*3��x�H�!������=���ɨR�B{f�ie�����b�Q��<:���!-�*7���D5��I|	�����.ŕCՉ����U��~�$N|	/J�֭�Gٍ���A�����QZ�s�����8@MΡh*����y�O~q�H(%g��N46/f a�q�]FV��z�2 M�ٌo�N�@`��b�G���W?#wiXX�/}�O�K�(q�����z�w��J��I���Y�]���P���{���aQ�|�Q.tZ0a����c}=+�3��:3����zj����	�}���3H1C[K�TP�d�o���/{E�bO�	���-p/��%��ĩ�Ԣ�!��c�x�!،�P��wݠ���<�/f,v<uݑ�:X�k��d���s��%3F����J��2x
�-����V��7\�\��&fi�M[�?f���� �j�`��W+�Y>N����3��qb<�X�s�(vk���O�f��Y�t�ƣ��d@�cX�`ԝ�􆕇���HZ8����W�X��'E��2Ŏ��%�r�EH�Y��=��~�mSt��;hiװL3c���S�b�h��Q�1��4,& �CC$����fm%,��xx�N��v	��։`�����,L�W���ۗ�A�W�(�������ܖd�7�"�~�a�RT��ى���S�Y����NZ���_h6��:1~����� �����9����t���(i��3ݽ��"3���vJzf��Z|�_�r�bF8|_$p��h��y�����Ddb�x�|E��>�c���M�^�Mh+'��ҲØ���?*�ܹ(�����K�I���-JۅʠN�Ж�\��5&�jG�3k��s�������P���]�R#�~�Q6�N?�����^M�ҷ�r8���x���b0I	|�
�����9��s>�3�D�-���A{,7^i����7Lj�Zf���W<By�&"���bɶvd�8:!e)��� �˺W�+'��bczU�q���t�jڳ�%��6=�VR�hG�u@\����g�+4��uQPR�<�̈́��؇Id�E�>�Y�����Z��8�Vr�х;�La�AF�8Ҏ��i-�ƌMFغvR�9u�����
�_ЇF�>�ń�A7��ZK�h��ȝ� (�.T/��owb���bߚQ��߅�@G�x}1i��e��Qgi����FGW�'����A�V>�9�4�l�@-�vc��b������d�xN{�]��e		LlE��by�:8���Ȭ����e`Is`��Շ�B'�VSU:��}�n�P2X8��E�t?h�W����|�2��xq��]ݾ^cL���� �Hk�Sg�qPw��Y*h�r�z~�F��C2p�\H������אb������ ��z�ڧײs3M����g���v��?�.�8�ɳFǌv��!�A墁��@��������Z:	i�E� VI��;(�<P�f�q�D|y�s7W;�^�98�{��+֩������խ<H��( �V��1.�UV]��3J礿ɀ�1�@͓X�"r@�� �	":���)�!�f����3T�Ti�3��φ��a+W'#��B��^�]=�-��$��},!0w'�D5��;u��#.��R�IMTQ:�#�;S�����G\wg��1!i�v}t���1�]6�Fi�o%��L㈫��R����) _-I�Fm�Q��>GPA�1��W���7ba���x�O����L2�b
a�'Y��v{���������Gn@O��|^��(bH�rV�����Ӕ,�^����4ǲ0hwS<7��_�=I��p���o[8�fR�N�}���H@>��V����B�#O��3�W�K~U��&O�Z��˘��@����]�}>�,�>;V_+
,��i��:�� ��-?+mA�+2	[����Y1��U��g��ڌ���$V+��!��I��9��焘���6�}�1I2�c�J$ ��3��j	����v��`�z��5�!]ۀq!�jz�	h�EfuԷG��������]�md�t�޾}�l^6"4�_^ �4�~��z�?Q1V�`���L�Y"�I��s����S8�L�8xJ�����5����=�e�;�@�2RW��"�Q��!��??�.��3�#~)9�'X�уO�ƤFL���z���PKԶ1)ph�M+{9|`>��>���	��jA�Z���ί��h�	���C��h���/�&�	�6RR�]�$A�{����T���9�"��ǂ�y�ա��ɀ3����n�Ig�8�7M�?�	�%:�c�Z�	��^@xb^��وg(� ��_H$S�����B�S!Ok����{N'g�y�)�W��:��)�JYrt�����[��U�"`((��tO,aϦ���X][�)��@�7����!��X�
����W�����fxjU�(����t���D20.�蟌^ h�g�0}����(,�����X���"�����E��׼f߃9��23�?�T�5q����' (����1�U��S)!�͚čKywG��M�|�uה��2�����s ��8��y֟����:Z�lj�[`2-Ϝ��t�Ԓ�G�D��k�d먀��F�����.+s�n�O��Ogyoԋ��a�en���]�Ck�0��?��
pS��B+�����i����I�N?��}��i��5@8K]�Gܤ;���w׵Y���^�F� ������#pͪ8�1�R��4�V�A;�#^��~b�����,
k-
)I�K:]�,TA���� (�Q���kე&b�5��B��.ԩ~9��Ȗ��VM_� d��^2�d�D3����0}��#E���	/z��ڎb��so<sJ&"��Y����� ��+שĹ��p. YA��q�m�2Pz�0^�v�3Fէ�;��QbZ�K[�ᘆ���9�@A-g�cL��q�������J\c��ckt��iju�ꡍ��X���k�U��m&���c))k\{E��v������.�������o��@3|�`P�R9��s݊u�o���.��k�j��Z� �	Y�P�֨��^Z/ȼ:?~r�����>��%H���4�W��랈���emx��$�@��V�}bQ�S4^���A��7Cx����XP��LC���P~����Vʉn��,���1�j�a�\e{W��2��^:#���*��H�����=lQK��\^���w�6?��`;ݩo�@F�o�ah!m�ֿч<���k�����jۈ��}�յ�F��BҸ�K���������N~{"o#l�z]:�b���AIwI�(n��"���O�ʧ뗗����:����,��NTÊ���J�$'nM�C���Ki2�b����mT҈���g}G�/3�n��25�n��-��H�y��qU�t��ߢ����^]�ڤ�T67��\�*R�'i��I�K���A>�|.�ë�9��8����E�����3jA��]+���MP�4�؛/��^E�B
옻�L�o�MI�qI�Cą��8C��yB`9�ί�/�Kg�������k��'�2uE:��f�`O(�VOÅ��7چ7��"��d�����)�}1��]ݘ�ߚ����q�b�Jk�G�e�8���-�1�;v�l�s�h�,
����JG0`��_�!Ө�=��_+��乥v��Y�,K��Y�"(�'��˚�Ftw��G���Q��x�%`����ᨦP�h� mʹ�JN['�ɶ={ZBj/�>��Ԝ�0
�ǀ�FD��^��OL��۸�4�2X�Me��zH,�N$�}"��������%�}����C��ہ=������\�a��h���ea���Z@)�w�K������
����� � ��0�t�����W)eI�<�;K㚿��,��:���d��ZG��=�Yg}�Xg�t��u�d�s�6�6~��a�=��³$��ȁ��7!��Fxsx=aX��<�i8>��]�5##E��,�֟S�6m���t�����cJ~�(��|�P^�5A��u��|٤���4L��V��
e�`9���o�m�;xm�Pc���k�F�ɞܔ���(2K��<�[[�K�)��F�>����5|��@&sZZ����L�i,���8�^�k�b+������	x�KY�l�m�K�+�x�Lbַg~l�~�)�0D�D�����9��X!���]%�Y̩�3�����<��)`�Ε�|>%#��������g� \b��<��X�3���y�7[	��jlaf5��8f}+��?�&�ؒ�qv�C�6§p���I�
e��c�;�������w).g�M�;����+=�2�`�Q��w��0�'�	��a�lP�8\�(�QCTźj�1�;�^Z�Zn>�f�	d��b��L8<c^�sO��F�CvE�}G�y�)3ulg���]p�/a���a썜�t���Qw[��b&���5jȚ�S"{W��_�g��x��j�6�B�8��ե%�h�w��H<^n{p��<����NP��D���J|���7	s��팫��q���?��7D�<g�m:�=�Tl����{O��K2Bv��!Z��ADZ �]�Lo8����[��E�sLO8��F�&4`�-+�!�![�lbľ��p�k�R���ȏ	��ǵ���#Vg��8
�ȏ��M�F�����vU�a>cx�z��FUQ��YI瞈�� f@����r���~$�rl��hZޥJq)��'��D��j�t�#SY#�EQ�s(c�q��#��S��9����tnM�G��Es{���k�͝:F����Ee�Qf}��Rn����{���j(_����3�AY^�üZ�3��o΀��A}.qI߰�p�N���+�pU�z�7�'t$�rA�ME�tM>�l����E��&.�ݟ�P�V+5�Y����<{�k��ЁrVM�$�7�>�ɫ���c�^���L,[Q���ɨRX�E�e�k���������q�#H�2��UI�d*Z�ڥ���G�e�~���v��B�H�#����a�S�*Y��K��(�\%��zi��j�0�y��4�I�QY�o��}}>�E��l(�M����Ɣ*�h>�Ҋ�Xa����_�Έ�Gg�� ��y�����_�|����IV�(����֛L�y���u��w�;9+ľMv�^Gc��h���^K���� 9��	ӭK\jg@0�l7ͩr4�b��g�5����w�9����`�`�o "'��t�_��p����q'���T,�J���[�XOb-���
��f~U�8S��Cr�/��F�$,{.�s'�p8����Pt�AHΜ��9��E�i��" �ağ<,���� �>��������*��H{�Eԡ��#�tL�:^TX��a�"���(f��y�LZ:NDi���ZW�!3���G4<����C؍�* g^���~7G.|8��
�44��������A
�~@:��kp���+�oA�?�#���ӫɔ�:�+��oA�'��Ɉh���"@��B���j��g�bmnƾ�fYrR�,��P̿���}ͣ���~��%2�:�/��^[:ζ����T�:�?d�Ö���/F�23̪7���Is=�Ƹ���u����$(�8�Xf =��G��Z�n/��e	���{���{�>)�m��,���J��5�;$����_��_NΆ ���Ӗ)�����w��e i��N���H���9Y/Q�(�^���q?����'u+f,2,�`l(Ie�Io�a:����FBY	?��������U�ޮ~�Ui����WD7@=#�������n'.e�[�G��r=�Q05SR]�v����ו�!�������$� �J�����7^D(���n7���q<E+���岾��!/h=�������M�0��^M|�Q�ߛU`į�f8W�p�.N-<p���d�V�ؠ�S�:iK(�����OK 2x7@��0�O�sݻ��)�&h��r՞�e:	qi�.���=�/݂�'`>��4{N��[�RVT\K�*�y�3����SJ}��"7em,���k��E!!W�.����:���n^9�B;���"�n�.�3f.<$ �]�K[;	'64�z������Y�O�GvS���h��k�ɾ�P��
���g�S�ȴ��f�0�[l��_��x����>}Ǭo���9��4#r~����}dh\�B�+&�ƂU���1i鶘o릛���?�"i�픝i�]ǎom�c%p��]vna�]Sh��Bȧ\��}?88���H=t}6_�_*8Ru�>?��A��hߊ��7�`f�L���l,|��Y:]��[��%r~3C�N�
E��b�<�N���	F�n�ߏ��Ѩ��-�n�#B�@O!�)��E|4�$�*�[�(t�:��OMtŠ墾��,�ߚf�1�zbȨ,���`�q��3O2d'ZKɕ�D��_Ie���հ��ʽX�T(�xn�}���X�:��/s�*#�P�R�==K�;n�s[��k���	{=��N,t��3-�3)��,���v�8�|,:�9�&�՝a{����QGfb���r� h�a�ZٛAzk�x3l�١X�nx+�߯�E$�dp�߿	��7�:Q3��4s��oѐe��0�������~�A�p\���PJO��,�1�$u�⋗k҅AO����0�;�Ƅ!���d�r��s1��lf���WJ]#����˃������l�2�c�m���r��n�d�?��1#5�2��o��5����g `?Vm���O��^���M���Cq��
k�N�����)#ɳ�<i,��-�9�}0�S����w�)�wU^�
�AI��n+�WQ���n��<�gJ�#E�}_2�V���z�Vۙ�f�U�5��P荈a@���y�P�i�si�J�Y�)ԞIQ��[Y�n�u=<Nr�6
s>�B�ʣ�0�S$жTq�8c��WK��$���br� �D'�"��-�i�	�wm���l��"/qvz�Ww��z��'&�ު�]g��c��*��3`�c���)�t��]p�d_{�<ڈ3p���]D�=��bm�`�F}vJ�Q��# ��[�(�bմ��h9@B��r�!��t�{�(�fx���J���� b��]�Y��v���<�z@��s�S�	�����Q�~��2���+*��ywl��;M�cMݝO�O�Ez�z��:���%:�Z(^LxO��ij�H���������J���Is%q�7�A��6*$�Ǥ�H?��.n^�z<�T׈��,��FF��ԙ[	�'��/n%��4[�B���y|;! �{���Z}pXl�C�����
E�B�k�}�BP�B��\�0UR�d��06��;J�^-�F�4wwf��&6���l<�y�(�|�h��jb��\�Y����<=n���"	>�����-�[���df���2:$�L�����(T@�dQ�٥EҒ=�yT��5�Ȗ^�����f�R��1�R<�;q��B���~RaE��Pk�P8�\,3T��TW+f7+��	�D�y��d���{�Oz�-�<0+�d������I���o�Ѹ�ˇ�-f������8����r]L�Y���1{�. ��7Pe��8�,�[W|w���9��B�~�-$�(�<8� ���fa�vw��]0�R"�j�x��{/�e��bJ����ҡ�ͰdI��a
UQ\�}_ρ@��
g_��X=1""��,��������4PW���TE)�s�8- ֫q���^��
�-���1Z� �:©E�Ф��6���6����(��$r=e�h�d1ߕ��능s�H�e|��r5tl����p)_��`�Z�#�{��[��ea���X �"���TFx/��w�6�>�f�,��	c�"��XiV���4��R�.����]$L��`�U���y,�[�u���r>�hU )ض�e�k����Q�{���Ӈ�͋�Ȋ.T�}TD#�a���x��a�>�&�4;N�:�N �;� �&������]�N��o����-5_DBM�j��2�GB�����g���R3d�5��p�$6��p4
jUr@eK���S���Z�zd�����|zzT�b+����b�nO�n�i������r\�h'ʎPܷ6��Yr�F���|�օ�r�b���kT�:Ժt��^]9�q����wˁ��9]b5ʍ)�Z����[���7}���NnC@g��p�H�bZ�D�y�c�sOV:�������|��Ky�_���Qp��	�f��}��qH���x[��Pk�TG��%��D ���n�QAE&18m��߅���TI��ӏ��k��GL���h�q�������N�����G�h���F� v�'����Z�h�妋@)N�`��� �TX�0�uEя[����Ѐ��{�"Th_J��N�?���Q�շ �q.�gʘygfi���u2WΔ�[�,T�j3͆a��.�'�T@s�P�19�nh��'$|�o��Wm�{���h49Äj��}��P��(VԂ�`��n��$>�<4*�9�
>紙O;���	P},�� ����_iN����4�B��-��)�	�B^2��0���1�L�x\|*����gpuxw���K�P��x
�3��%%��<�>˟��n��ef�	�m�ܻf&Y� ������F���L��$��� H+8x�-�vNF���U�nu!�� �5�H����\�'����'��}��'G�����	o  Q��V#�}�iW��)��	���u�30��g�Aȡrf'�j�5��z�M�I2r��{�뢫��ݾ�˻^�p,�T}Ȫ��Gu��ϳɠxC�ʿ�)
�9�e���lE�:��䋥�17�?gF=mI����e ���6�0Y���~y��=s�ݲ��+!T����tEc���s�&��b@�C����#��������.ki�(^DI��[5��6�`��t���-]nW�,TKkS�[�g7���p�R��!uj�Ah����nrf(�f:^�^	�#6���9tPv\2r�|E2�%[���>���B�V��	�Bi�_C�3r`�_>x3��qzV1.�������٭�0�d�__iYN�9,f�������$�J�+��dm���*`�r��s]<���GY�Og��_�����Z��w�N)��`�ic_(Z�#��m�Oݎ�@���Hd6�#®t�bЧ��,�Qq�6�b���]YC��_�X��<�\��1N�L�y��lK����>6׭�A�=y��밇����O�{r���g�6j�DL.�Q���=R�Ͼ$�C�ɀ����l��W�}��p�A�(�qb��HpoyX~�e�r�MB;#=Q����i���[d��1I�y[��^� ��0�}D�2X�� ��47�>&�����
jir�6~D��w�������������Ǻ�D(�8�]��K��|����&&� 7K���0�=>��}�Z�UI!*�I/D2|�Ϭ�$�ԍ�9HD�\��V.�*��ȋ�w��K��u��r��L�⮩ad���)̂�Y�ѯ���V�B̕|�,З����D��Le�=܇�W]��d[��F�vuf#���g���\sĖG}�P�@���C�G�[a�SI�Ұ�>��a�jsH��;��CEl���k�E��7'�n~�Æ����Ⴐ����`Q��z��)����ѹ�W�D��y�s򳾂]�c�o���+�@vԽ�5���&��$����^�KUP�܈k�v��)���6�	4tg����Uը	
��2�p��hC����PF�Xl�7,�i����hqzV�O��Ce��#�*w�k���S:�#��$�1"wE-�V.�t�]-Ql��-���1}���a��σ������!�ꢋ����Z�c;�C�F(
�����p�yZ�^�Up����!(L���?��n�m'�7�#6�z%��`Y�����%
X�cZ���1p�ƾ���\H�2�N�??�q�ߗE��53F"�������
l� 2���V�v��z��w�y0�Ζe�,�/L��/'E�q���Ш�{x��Q�y�Y�0[�{��7��u�P=5ĶX{�0؍�6��;�2;��%#[hliس�($b�X�:B�K��G�x}�D.�s�?�B]�oiH�:D��q��7�:��� �nxj>��Q�Bȫ��d	2[�B��W�*9w��xٿ۰����1��������b�ЩK�˃�s1�
�ξJ�ۅ���y��o���� �G�v*�=����#���>�&uY��i���[��U7{����-'��Z�x�"4��Zdz��|�L\�	�ȑ	�ym��K"�7@)^��*��;��hk��ڱV�Ux��<�%��7䵧���I��s�6o+1�m%yp�����5�qR�N�$Xh�N3A�wЂ^u?w�r+�R�F�ar$_+z�����M5���Y��O;��t�e$#�P*�F4�Β|��U�"���6b�3��i]32W�F<v��� s��7ֶ���2F�`��,���JS��\��/7�q!��N�M1�{�Iw��Ӯ�M�-T��[CY���B�2��q-��Y�����l���]�
$9��9�P�ёI������k�͎��Q�\��í�t�>��+�C��jb"EB���.ޒ�!-���Gw�b�ՀIƥ�����"\�����Α�:�� p��>���U�Y�����T�rh-�uek����\Z��_��q#5���?)�	~:o�T�'��&6�]X@��Ϝ5��$԰=)ʽ͏�fM�j3���ӳz,[�T�x<�%lly��X�A[�������**�j7���:�,d@��>$� �׿���I����~e1�	���*b���5���
W�|�?�--�c�� x�?��R ����t{iꏫ� @�ж��d�BD�N�w
�X�~��2m����F<�q�V���'�@Ĭ�`O0���)���`����ӻ !�J����q�ԃ�*N�����������p�E�-ب�-^�$����S�������&�AB63%d|�X�4�W �|#�8�~~{�~͹��������CXx�#�м!P��9�Ԃ�&{tM���_�>[���>h�ՁKQ�z�[$�h3��~(���] ?��(pG�Iȧ�B��NH_���NO(�^�b� Nߴ�&����� }V����C&�o��V�W=��V'�6
�_Ύo:��
�g[:�G� <��긙��x-症�k����W��8;3*bs�r�!�a_i�|���e�Xmց����'iS��S�d�i��)��26�j��9/}8�jp���n7���RS��WR�E�
��V {�@ާ��8�:�P~� 
i��ا�%&/�y�N>��T� �,:�e���nea/L�K�X��'��j��-w}�ى�হ��h�M�!v�d�'��\�s���F��0Ðw�� �1)��/��u7�%���`�TTu��$k����CrS��Yd�ME�<^v���+{���]��hu��|��3*b�!M�`hz���.m��cu�c)�!�;q�-�Ѩ�?���\���G�>Y�]��r�C�I��8	-��g�����?�����i��x���4��-<�,e��0�O���Նִ޴ȇ�c���/��7+�Wz(ƅ�3u�#՛_J��7^�+'Ÿ;�Mً�/��O�]�(gN�}H!��]�"���(���o�������|�PҖx�4�|�wß�w�t�6����h���oT�/��ٺ���R�T2S>��*!�3��ɆK �R���=C��o�5Hk�������cU	�r�,J�dR�:)}m^�'31i^:.B��w�Ed5���>[ ��*	��;�^p��&��j|��p��m$�s��^����_{Q��C"ޢ.4�N�]�$�\��4-�=oKv�snQ��j��Q��� ل.#��\���{���m>�t��@�.$n�]NO&7��H),��A8�c��=����;��q/!AG
}�$���S�f@s�/�>�*�{ӂ��6�J��D�&CJ�
��/Q<�Mփ��X�S��c�"a���ɟ�Տ�;��>����޽�:x�\(���CK��
c�X@��|c^q�E��3m�$PG%=[�
sԣہ�u���֙pkE�b�o�`@a��VI�?Ś���QL�6��%3{��TQo����>q�����·'\�8�?�gZ3m�<����O<r.��J�־��,`����c��Ϩ����ߢ�4c�����xK��c�|<��;\�t�l쬆_���_KS���5�A5{V���Y��L��O�����Az3'��7��$�&���c�xn��m;�Lg��
�����<��9�5�s_M2��+�v*���3D�%�7ؓ�������y~�jѫ�t��0�Vì-�t��w+���tN��B������_�h��,h�5��4v/���_i��ĀcV�l	1{��ь�V�C��R�F��tU�I���2�M��b��n>�HD���H�yV3�e�ݤ�dq(=�;
���Bz�W���ؾS���{gY/0u�N��L�~N��ufV"���x�ORd=���o
�!�F>@l�>E����5L�a�T�@�I.�d��-�`�$N_kL���LGe�-�����✁-��FY���#�O�̋�W����rS#�O����O������[&3�n�9]�xh��ߣ���]<".�<����N�+LY~=���#,�����4G1�qMJ�c��z���L��������2q)s�K�'�0�.��2+p��cU��GX�m�&��'����@�3<Tz8���%3nÄ���H4Q�\��r�~P�rPt�F�Ο^��v���/O"�;
^bD� ����Ҫw���j, ?�J+ъ8;u/7���܁!�������+D8�6(�C����B\�'F�I�A��{9���քu?j����K� �%+�M�^S�����˨"��j�z�Hw�`�}��3�V���Z�׼
�������洫]1}4+9�3�n���р��G�tG2x�P�o���j�مq%5�6C���5î0�vq��	��9�;�w����qA���!{�l��*4��pMgR�W����{Z;�Q��:�Hbf 8Z�@^(���U����Z�UU����W%,t1.3����|5 G\/�[�A2(:�IK���YO�iBxD��[�$IVi�sA���ݘ.����~G<}W��6�!�(��6L�]`|���pF������Y#�_�0@ӉA���ؤ �vŤi��'\>ZnV�eJ�=q�|��[Π,`^�1*it�j� �������w���q�}��1gB�/�S,�w�ݽ2Br�p�Ɓ�/���vP��x5|��dVd���<"�����^>d��b�D&�� �;�s���o�1�����(� ����)�����r2Tؐ�9^@�2��1�mǒ��y\VH晏�?��0�5��A��4,gv>����h��ڣ?P���3k@臀��۔��������7�Ԯ�D��=Ϫ"�{ D�rJ�'ֽ�@*�*���{"�L�X�Ֆ�я�-�E��z(�'}����]�F��%����a�e�Ho��+�ۣ
�[�g�j�����ɋ8L�oќ_��ԓ��_���5MHe��F�����ʏ�X�n�X>��E��ڨsU��mP��$ʕl�i����?�p��5{�M�	o4���?�>�.�O�B�U|��N�iB���2�+Q�-sv����&�����@_m�j�kRd�ˍ3=;��̅v�-�|�V�BdP��/�l�ę�����HJ�,(!^M�N[I�|�$f�?�-�e.����tn�3&��'��DC(7�����n\�t��3�*$?R�1	;�B�n�v������T=��r	��p.��v��/$�ɳ�2�@Rd�s����A���)�,��q��AqK��	���4�0��s5a�Չ��Z�m`��qC&���(�l�bk%4�>��d���]>�,#�<���i�o��-���� YN�й�=���7�p��� <����~�JՠJ�ET�h.���渕�8h�TP�Z9A��+`}�T�6/�ϨrB�&�	�`�9��9�*�R5{�69au�2�VYb�k�Ѣo��u���3�k+��J�Z�/W�!��3���a� ٚ���K�1�y/��@��C:c���]��9C��HTUb�p0[Y>����ߖ�Y ���)�Ӡ���O�����&Ԓ�27+�e�Ҭ�ܻ�h�(�,�H��Y��l��.]���-�bV(���'/b���=�����c��j�Y�P�;�bh@q����_D�y	�N�C�`-l�,�]a�zeS�4�ZN8WHh꒞|T�w�_�إ~����}S�lY�������K(��_�Yo���,�s���<ÄVf1�A� )E'���|�G�oơLuTFﴧ[�� hK��g\��Fs�����ϴ��:�X�R��fc�G�n��--��G��.�16�����1���L#��$��$"5��_�� Mj-R o��`i}2z!����~N�qN���ʧ�LT�~w�!�k�Ē3��淪N�
�y};{�7��K��>dn85�lp]���.1�����*�>�=�D� ���W�Um���V����۝U_���U��y�F�4]��<9���%D/�j����FM7y(�:������m<@E@̳��h���Db��@T�^	�XVXأF��������3�u��=�W3�o��)�w�������<��gmQ�Z�(0�#q��?!p��Y;�eښ�49����-��,BHS�y翠��e��7d5��ʃL#y+��z䴒~{f:���ɦ����j{9����o�:$��/���<d���y��개P6��-�d��&���jĚ��xߵ��z^���>�(�@���Ǹ��2�"$o��3c�����?����=��O��H۠?��7WP����{[1E�}>��x��^�u4�IbmjA��Y���O+퐟��z���G�Ϯ�LT�,���{�?�������5%3��E�Ñ�x+��*Oc�Ɏ��T��Y�$s.}��8;ʚ�҉�ШE��]]��$���I���K$��Nć1�H8a8塵�l���e�SƘX%!
q�*���l��?y�H�cR\�MW ��=0`���K�����g}Q*/�J���h��:��F�k����!����y\mX���7 ��0*�d�$��H�O��O���e�z�E�&+Bt��O���Dau�<Z�[r��C//:L���8Y�H�G�i�t�	I>O���K&���˼˓1g<�R`��s@�['X��ؐC*9e���jm��y.� �7��'{p����ٗ4���EŜ4����A�e��4-�8ۘ�`RD&Δ�JR��w�-W��i�ڏK��3��;�m(Oָ��Z�c+�U ����֏vA�9}� ?O�u&���c�	�,Q�F��+�,N�/��6;s���k�cB�� U˸5�<[�0,ddl�0��?#���>���zI���g\��=z�P�,�j�+���PNԝ.�4L��n��Uo��P���l�AG�ɣ�3ȬRGPJi�.�u�?O�v'��~5f<f �`S���k�M�t�N��
-�����ؒ��v_Z�f����@�3���;}�V	N4�f.5�7�n�Wu�7��PR�E�ڿ�����d[�q��5Yt�G��#R_�w^b-����-�FF�I���#� �;��A�y�P�>�mS
��K?��xFk<w���Ҏ:`%�{<P��w�k��1t}��NPW��+�C�:��wK��|'��"�	7ϣ�
YN"��{v��p��~�,�B��Ǆ�=�f�`F�^�h�`lӁ9�����ש¾N=@���Jy�b��/S��Kc� ��l�ˉV\}0�M�t3���ܧm܃���ÜM:ܤ����1�Ӽ��g��1��P�P��i�U�C�$��e�Ǚ����ϯhl�7����F9�[�@+�𓍻�dh�Ď*����p�T�eI`�e�)�e�D��X�Q�*V������	@�����й<	�?��*�_�C��;���]ͦՃ3�r\Q����'/c��߭�2Lk�?�D���.F@�"&��+���y�8H���7��O��L#@��(�=l���0�{܅ �m���?W�n �U�3x.��~3 �	D�l��B<���VO;
k�'��Y]���2�*�ز_]Q:��\�M�G��8�G�eI��9V:-D�6;�����R�Э�OjϢ�-iK�Cn皨�"	x�v!�*Tl���a�u%�+�{ 4A(�꓾�j�}%�P���ߣ��9<�&g�����" L���PL��r��L�wd���Q2(w��%�'�ֹ��[����e���9��;ʵ�G1���%��T���-��x�����a ��8�/ң���d���LVY���̕,��t��+U�M��	6��⽃W��{>�"�h���0����o�6�4�CMD`��Vm$1�5��_@k͞��<m��<�IS|���GeO������������~w���t6w�yWE��c �S֜蔜��Xl�8���g���r ��:�L��k��F]�����%߭�}`�vӒxQ�0�*���GH�ƔO�S�5�+�
�ǡ�ѭ�"�M�ۤ�J(af��������g�6��l��%^g�����d�nn箃�r]�BQj���>[Ă�2�#J:��0������M�6 ���99���<�%wcPŽ��2%�Ku���8�������i��46t��;TN�ktE�[��u���놃~=o�-k��%xv#��n.>%����de����.��i�E�!?�}a|3Ɛ�C2xj]M��5�3���g�	��<p�5E�� ;n�>]3ERPmT�7�tL��L��"�{R"UH�"z&s�D6���@�Up�9�1<�BDS=���#�5$�nPi�H|q�4�H������)�z#0��)8�tÂw'���<]u�ls	���ƫt��Rs<��J�`���M�Ԧ�6?�A(�`�d���ƃ��`�Z!a�ȇ�F�a�����/T��c�G����$�����%�w�O0|�$��T6r���"S��O��8N��3�Q��O7�՟{�z6.,BZ�mB?0�D ��Ej�2#|���r�J����Z�kd�`n�[d�6��I�	Q�0���%K�&_huR��m�[{���s����y�����A���Q��r�IX�1�Ő�otmy �f���;�F!�(�x�,:�;+�E�Aδ���J,�妵��K�����K�f�i$�Bj�� ��&|����SڰoyXڮ,?���tr�{���G��Qɓ �����@	jU��X�;t��j��c_L�U-LFg�V��Q�������+5VB!��ѯt�h��]�%l�������X9gX�n��H�hy�Y%7�m��SⰔ,�	��t
5L�P���>o�ƻP��lI�����H&St[CqA@[鎚(i)�bN��.�S#�)���=��3zĽp(�<���b���2Ud����l�v��(��ι�F��`�jY��yfR!�� ���`z��t�W�تQ\=�E^$�4ح�&�뽘S��v=��pg:�a�Kj��xUB��07�ůwV�7�G�Sџ�T!���@&H�E(�5��/X�{�5�'���!�����,�߹�*�����K6��X<Ƨ\R����,����j�����|�B����h��Hn���9]<��K4K(j`���աP9b;���\�;�O����!��GX���$�E�I���_����\&c��e���9�+U��7,!��#x��}k`N6�V���E�xM��h����E�;ŒoL_R�f�Mq�	�����Pw-�Y�X��~�J%����t憧.�5=�W⯅|]k*I�L~�J�Ʈ��"����n-R��7l�0��[<��s�'K	G��mg�z���\���ׄ��(#8��ߠ�6�}(�������"9��l0�HW����CD�6��v����.�AA�:�g��K[?(���>@������ul�pO�%�S���`y��7�S����6�/�ţQ�)5:9����Q\s���3�oq�'�.C�&
'0�
l���$����o6uaڶ/z ?�P��$b
|��`�3��������x��	;�į� 3�� �2�PKl?����.7
1��w�����~���%s����c�/�x�0�l�s��&�#{ձ�Ʃ�3�a�*S�=��٭����w$������X��"-l��,��f+�U<��h�V�A��K4K[�����݆��-v
�U�R_~�D+��U#����*`2�$���R�K��4p�!�&n�F�@Z�fu�yv�֦���ߪ9�{��to�+!�˨R�wᘙ˂����W��z�Qx��)4����HPV��-�*���KvؗT��A�9��-�Əo�ѭփy��\ ��!��S����F�b
i"�4�q� ��k��kI��ܻwW�u����D���A�րuN���9l���aG�Կ�YKO����`/��#Q���ù��s��u����v�;�ѿ�K�M�>"1��U+8�hG�V9� ��Rb�.�W<<핍�k�P�, �ǯ��x��/�V}�{"B}H��u ���0D���$Q��:�� �<4&����Qm�砲l���+�^)��lf�������Ĉi'$j�H'��Kް�@8ϙ�kS�iuS���e�cс'ⳙ����*6T�X>k�/�y�CP�ݕ[�P��/O{z/�k��^���ű!���hy�������d�6V�`���Kp������@T��V�[F���t'v�k.?)*����y�јأ�aq �H�`ަ�d�X�3D 1�fONs�s)I'�M�W��LK)���6|A����-��y+�P��X~�6�����î礠j�:�e��V�	�\ey�Vya&��u���{����aH��HRϒ��9!U�}����T��.�W�<��U�4v7��q+b��O�I���(�_���!�f�����BLp$�Ix4D�,��S[��	���xG,sԃo[�9��3PYD33��\��/N�\5VZU@����:�j�dD���qG��c����4�W�B��}��R��h��U�8�F��5�=�XX&�.,��FW(b�6Z���0B��Q����θ�_�"����n�3��8jl�ǐnnV�R��/2�c^YD7���q�)�׺��ce��v�=?P��d�FGP���c�|7�PB8��w�T��V��r;���~n�2�̪|��Y')�c]�[�����z��Ag�:F_$���e�C��q����o���\�=�l�Wf���K7�H_�j��'Q+��q�[mK���r���T�	�<N��ǯW^�ڕ^+����E7X��d���ZK��ʺ��׊�����bK�EP8���Q&lP�����h��ā[�\
p�MЊ����-���e�|��ܧ��X�آ�ƥ����4��V�;$]f������2�_��Vh|���Xq��t��?Pّ[�� ]���zx�k�D�	F��3̇72�X�_�WneW����u�n��K9]S��yz_�v�KM=��E)��)B�4E��7V\AD����7�̒�iG*x�Q_y��\���9�G d�����?��
uuOR/γ�z�T��Y2G����Nn.ڮ�)-a�K��%®�d&㉟2��n���"�i��c��K�2O���)����?�H)����a�9d0C�e`Vr��0�>%`�\l����L//�_��%�kx8�r$GO|�kɘ �!�~G\���AW��� �J�ES�͢6��h�9�����P��u��Lw$X���<[N��_*B�1K�s�f���?ȍ��jf����]Q)��f�ꂃ1h:�i��T�k��J�x���=�ߡ�wC �3��`��H:�9�l�`�_8xE}u�o��_���H��'*Ə��>UN��qå�b��rû���`K�<�L(U}����O��쳄q�1�F�wc���V���\Ϭ��T�hf�u�710�E�@�����������;Y�:�e��@A��NZ9k������)koa������ܭ�0;0T�X�DZ�	�R��A��)�Bn�w;�������T�)vPY�z�h6���8���)5��`�V��H�9í;"֊|��C8ڒ�"���a�ڪ�*v��C���O�&ef]UW����A�!)RM�&�O�RA]g��{���Kz_W��;ـ�&��v��"�Sm�G��W����'ʔ���(�Q�\ʩ߃K��jT4�.��]��Qk�]����V	�s6v��x�2Fq����J=�z�jG���9&�m�9��ȹ�$�0�����CLR��<,��,���K�oT���6��{�������*%p��')����n��+tu�g���˷����!P�ʉ���(� h��E��Y���{��!!au՗��t$�{�;�J��)E�����T(s.�8%N8�<~�=�)�/��Т9�{c(�z����	��GgX�̈c
#F(�_��^�T�ҟ��=�M��{:�$�w����K��V�b� ��9&���$��%�[2N�)_�����T��2�Zz���R�HX�K���,���;	S��o7gUJ�$3P�ycڑk҆��l��X9r�GY[�p'���YaZ�	m�W#O�� z��� �Y�5�W��vъ&��H�\4bK���N���ӄ��	�[�����(Q�����Y@��6�D���>I��N���"_��{���$�L�*��� �����c��# ���C�-$|����ur����`���
�y�4�"�*������E<��Z�܂���p#�~�3dGK���+5�f�>�s�]Q�����z0.A������l�� ,z_��o���%j�Cݺ˝B��_�֯3��+�(�ߗE�U9�� ��;6!,�e��]�M.x!J��+� ���Q�r�,./w;7��k]qF�c�O��[3۶��`~C �qi\+kA������'�g<ڞ��4O�����D"C)�sCQYI���Ɠ&`Tz�PHznI�阹E�=��"��p�o�Aa-iM��d��J�bR����yRN&�"��'R@��~���qp�����6�?��x6s ӆ�����ha��V�Y�C�/RZx�+d�Ay��?��85=zi���,��?|����A��d�RE���q��i�<��t˙�א��^3,ռ>&܆>�� 诉��Et�m�UO׹�9����� ��7���!�.�� �mO����B�D���d�,�h*���A�<`�0��Xl��Xj�n�~�y�'@ ��U��FU��3��qg��8�;��-�.�A�¢bP(�P�@�Z�旱��[瀦c`�w�R�u��k�@��y����sg�fj,^B�L��_�~nI�ؽ6&y#��;_�9��Hf��~�k��X�]�y�7�aU�K�e���@���=�'�.7��ǋ���{�l9��D��xP��A�V�W�c{ۍ�ڦ�V�R0n�&j>��<a��r��(���ȯ�羧 b��`1C��?S�Z7��rM�\�mx����Y	;yH��m��H����%�g>��ΉoC�l�my�h�}S�3#�:!�j��i�Z������Ҳf;^^=ʧBVP��7�K|(�q�ݩb�6�;�?[�퉋��2����Tx�s�f�u?�_��諡��CS>�k/�9�5"����b��r�|/����������8ɻ���>F�~�e2,�|��9k�x��$��%�~w�05���;s�~��L[��(��.�(w��z�� l_+��|�Kt���7$P��KJk5��<�����
��Y>]0U�j?��t��S�X'^�3�㓷�����dy'8���[|����'>ܻm���ʀ�}*�Q�iZ��R���4Q+�
̺W.�K5Qw"m:�@�u�TLؿ�r�6+�H��-��̒9p��;?��*�Y�\��$�?>vrh=������o�'/2&��x%<?vFbi*�����ss 3gP}�W���i�iq������d��9?�{A�8�R�nX� Ih�;�E�p��)e�Z��mG���w	�} �jc�B��R� ,ӹ�k�ɹy8���F ���JU�F#߉�3�n$b]t
95��F�X�Qw-�v�V��)��~�p������);S	��8"QA�i�����E#���a�L&,j���?#&YGņ5��8�s��Mz�C�����%!B�
3���Α%�L����5�K����%:�=��2�[ !�����X�Lz�~8��� r<q�����(a�����M�c3R�';c��u�՘��F~C�)��x�5:����xH��P��W��~0ʲ�SfM ���S�y�C*�Ζm��h���4C���y�=
�@�����h�=���n�2	��~�Wb'����gu�G6�^���/O+L1��>O�n.�$�8֘������џ�V&��+eY��
� S ��<���ra*"'I,���w��S��..)�m���Aƻs��t?V��x����m�x�?��9%CΉkR�RC�mdڗ�5,j���X��sԎ���|�5�;%������Á@�jyX���Qh�|�����z�Z�5 �j��Ϥx�춱�5vd5�yP�VP��F;Z�Q�Qڟ�
�M��ߗj�^/L�KT��(��XJ#ؿm��e5�0��Q��Q7.w�˷��:8ľ�P���9��`c��24�k ���X�
�!4�|e���F�b��
����kwR6��]Y�
�����PJ�vI��agޞ�9�Ȟ6��/h�ã'��o ����� �1��yKK��=�RE1vغ�>��9�%��W
����c�Η�%���zZ�W��Z�ڿ���,hXi���B{��905�߽�h,�j�M�*�����\2??��jݠ��%�Q����dD{��s�V�r�q��}m{�����âV��/c>���/�(�v���s��xU���D9�F��L�If'������J������/�1`��@F-E�]�^�w�+���H����1��h��Px�� \^�$���o$�c��K�����ex����甴S)n�Xq>I���R��"-��� a�+߰a�EhJ*�ImͼN��!��J��}�"��1g�}�#��Ξp�)����1T.�3�����5W��;'��f����˓!�eX�-^��^��T|{�/i�������Ϊ�⿎-%��
^�����,��i!т
�0]9�sM�?���ќS�U���b7�1�̦������D�Գ°O�Z�rִn3O d$����U�iρ��Vf�7�r�<��揢6+4����Ye���L�<���|n~6?b]I|R]wS�N������i��:l:G�r��ԑ�VL��au���v�ӥ�B��V�����S��!�io鑒k\N��QW��ɫ$��V?�/��n�cDh2�C3!�=Z>ށ
�~�
��z=z���qYq�^����,퀌�L.�Д��P�$���Knu���6e}g�V���~�ң�d�Z�i�MС�vm���f��Q⟚�0�������=�S�J�H^���̓�u}��x�d��fA$��9�mc`��}֤F���������}�����U��	#���\`s�8<��W9v��!���;��V���J�D�L���3�� t ������F4��j��@������S�П��ԝ^���MB�Țb�n�GB��)N�gb��)���,D�p9&�Ƈ�x�.I�H���Sr�I#���95���{�f:K�-|2���آ�A$�+��G�$���jn��y�D��V�)��TL�d���Q�E	V&�LB�=�&��Ġj���i�op�G��{�$��$�5ze*��nW�>��B(��;8� -�U-(h���0O��V�Z[ۃ q܆�{�jиwƱ���5��̇,G'y�����V�/�Ӟ�߈h%���L�ӵ�̾��$6�k�ۚ�#���ɪ#�e��g���ԃ'.��(p~!o������7�b�5$/ 8�TK]ӆ����w̙��塚X���c���+nr�|2�v z��o���9˩�� ���]U q�L�A�	�2�=(Ǔ�q����g��ą������.�`T��^��̨ueO�����~Wvx�NX�[ۣv_�]����CW��'b�����<�F��-
�ԏ�0Ko9��٫I��B��яk���v�T�V�柭6!�&-]�JǨ���܃�T>�F�`*���~�r/����Z��{�N%��8e�οXh��ұ�!�J�o��$SA94�i�����e-�뎵�ο�a�}��b�Yc�\yu�n52C��k�eN�h>Xo˗���y�f1����2c��m����rfꭽ����1;���|[}�^����1�D�T.������0ӛ_��0D /�=�X�?��&��_M�a@���ʏ,c����@��I���05S�<DK���́���
g�U����L��"_�U`������G,,#����>*W�x1�ѡ��Udꅿ�d\��]��åd�jkL9`��;�j��%��wH?݉�L,�E��Z��:4���ǩξߪWԘO%B��C(�K�f�r�}~fK���Ϳz��*�f"tF�@/(#�V��i�O3�p�ot}t��4�Y@�t��Cf+_�S��k�o��s�V�ֆ�LI K��#	.��;O�r ���4�7Ǒ��:w�kZ�h�w��M;�O����-�C��F�1v�����2���\X�8R��v#�Qx�5 1�J"#I]�Ϟ��t���.��R"��d��*�+��w��BS!�^�B�x��w�/�����Ӆ���~�@}F�HW���c/���9��cK%�7�N�n�F���i����֐��,b�Rې5E�؛B'>@�U3��a�t\��r�,O
��ؙ�@�J�+���o��3�6r?4�c��i���?<����@�Zdڌ1��#�}��_Qc!��j��H,�ؽ]�~��(C'l0$�c+غr�Dx܃혴 H"�	���6P�i��H͈*0��S{�����4��t/�.��|F��pnu?���Ҷ}�+��_]Nf�myG/�b�	N���	hN�j:�,g��`�͍I�pM�{uK`r}$L|d�}R�r�4�˕�	��g���/
���"u`�3�V�n$�ۼ�Y�F�x"j��h�
J����R�VJ�-�s�
�e^Ö�G�:���r�1�Ͱ^f�p��GZ7�'��x��ro]�q�P'.�c;����w���`G�����i~�Z���m����sV^ʟ�U��m�����ꊼ��i����!ǐ������^�qm��sԚ��P`+��	��G[r���=�FIkq�ls���8��,�����(�6ޙW�[.�(���/k�<5��J�9j���������X��U�s��(E�h+Ѧ0�zƬC������ӱ#AC�O6em8�k��º@�G��nE6��x���(��o�? �̂J6)����%f�t6��N�$�3�����"[U�����Z�����]j���cͿ ?�)$D�{�G���x@d��n��uL�����}o��D� SowF�W��r��0���V}���L�g���#�:�Yev���j4�d����w27p'O^�z�/V%�"Ճ�O�x	ԇX�SO�������>΀��D�L�6_SuN{���'�Ǜ2��j���Z
'U������=�z���͞�*hf�h�;���OYBԺH/K���b���`0��9bO�pYpLBa�w�F�/�F74|&5yvd��
vs���Ύ�H9t��b<m�S;�Q�8[#l\��v.uV�6B]H��!���E��k��t�d�`����=���`G��dݥ��jj7.P8�0��k�đb�,+�z�׸X�9�s��a����%R��_tǞ�3��,�B�\�p���#��[�<5`�@9v���!*�� �a�e��Dc�Q��yz���F2���H�li?ux�WF����(zS�xܺ(��wN��l4ͷ�i���h��+*A�>���O��姌��|��ԖҲ�+�-)4:�pĆ��+�r�sA\���-�*��K�)�� ��?�/�E�,��b�('�I|�6;�VIp��k�B}oj�tjV�X|DQ�o�Պ�V����`H+���G&��*���R� &{@ݸ5�ִ�S�Ⴘn���gաQ�U��8
f�z�$чO�Ku�m��ݜ��Ǐr��r*\7�F3��׌����{S�ﻼ",;�o�ߧ��2���ަ�r��m �T�B��lޭЋ�m��+������@��0ϒY��:�赲Ȇ��0c�m5L3�ق5q~ȑ4"37?�.��\^% 4���O���/�'����*Lk*�"���?�^���͜�� ٌ �3�l��-6�	�iO��S�)���
�o���Űh�$D���O�:Ū��v7٨�vL���ᆥ&<�A�~�kyW�q❏�K��d�۝�l ڢWh;�f��t�/!�S�������u�ɬ����LH0����6��1�R#��Ӕ�#w�5��ֽ��V��2N������)bB�<X����)7k&Xу�b�t�"�ш����HP"-io�O��'�._�{�:��� * K��
�E�.�f���r���lDA����5m�Zn�|�2���ɽ�e����/5�����BёQ�F�������[#3�<�"�bga������^MU�����Y>�� J��͋ư��������Sӑ0m/���<��w���e�Px� B����&䌁���~�m\2מ�R*{}�5�X���d���ƃ��<�b���njbd�o�L}�Ҝ#����؄2Wk��].�Ք[�-��D�yc���oc�- q��S�B�E���:bi�K@�y]�aGp$p�	�}��-�������2��h6�
Ie�����F����,Y(�T>dX7R�3D��2����a�_��S��m���8)B��"	��؏����(.�t
j(��HM#��^�p_ƅ�$�$sm���m��Mr�GҰ��X�a٩�� ���U%A�X�>?�����v��<�f�O'����&��J����8�z�iD�ߐ �e��rz����N�k:�������Ң��h�%9���nN #��6��4 g&�Ķ���L����]'N���1�q�cVjڮNCג}&�yL���$n]?�H�����ިn�� ��Fa7�w�Ը|I|��J�r����',�[܏P&� ��X K���\��q5{Q��;�@6�=E�}� 
`�~)/^=�:�E�z
�_�ޔ��^��МL.`n�	�B@x�oyɥ8H�
���밴�Al�	nV�;�M�J"��
(�O�A�S��\���{�vl�K6Mp��cz�4%�5��hp�V^���Hqf�"SsɽU�c�\V�����iq�96�ɢ`h �"��K�n~.�o����/$���qю�\���,~a8EE#S��[�4;i���T
��L����w�T\nRݗ������n�ꆮ.�K|�㠔ҁ�)�k��B��_�x�lF��b��T�۱�
���i�N��JŭkY�o�y�?T��7�<1
�S���S��p�Wd�-:[��1H�q$(����&�.x��vܤ�0��Z?�a�0�t6����ݽ�xNE�K]b�K�~�̢:p#"���@�k�йf��7MD��RU���Z4���Wo'Z����N���NrNF�M����zڭNx�QgH x�"�Z��v-�7�γ�}v�Gq�B�`r����d"��H�]I��xx-�.S3�[x!l���>��-���&WU�����\I���s��?���6�
y�x���!i �@К�Y�5�k�-��d)!�*k���b�v���%���jA�L~	�z������q���lr����9PUΙ��ފ����X;�����g��͝LÔf"ӌ��^5�G�.X{g�3��/�,ݚgo�@䝃�ׇzq�]��[����E����ੰ�	����]S�HܺZV���F��/V�f�����)�f�3���I���T 1GP���+"0?[1�qD��G^裨�C������u��M�D�/�\��C�z��Nuy��9�8�3�s�����&/P+����7!+|��a�ɶ?1j*��l�.��W�l�� �� �$�)������g`�1�?Z�F�(�nτ�\m�<,�����f.]���zi��`pz��J�C��d�v ƪ\]C;�M܁����{\W:�ov������$fޘ�ޘ�МB��3J_�$���p�8Pt�y%�h�*w��t�Y�/���Os�� ���UʢX�9D0cA-H����vF�(��}��y6B�����`m]Y#�f���Ri*%��]�~n-�"@;yӂޗjf���Qx��+ ��Lv��'�))k� ��_R��_s(��f�N��.`��Q��4|둟�H&X�+%���/���t�#� ��)��=:�.�J�75�C:[bh��N_��7	�����5�3�D'~e��zA��.�+�$�t$�?�F�U�9,1��t��j�>�/��/�v}Tڃ�|�����2�.Cxd�ߊ(�]���d�?��U�����i<�#�WM��iC5�څ�3+¼<���h�)?c�C�|�̥����:B+��>��;T,�_I��X���( ��=��� ��1���o穩�J��MVQ��o��@s���E�����f�w��H�xg���j[BO<	��#�����VHѳAV�i��(��:w��M����ѿ~�R�iK'�q�f����9W_'N�>�Jj3��N|�г�e��-�ub����Y'XzԵ��r���.:N/3f{�Օ#���.�˫�5���۶76X
����Nz]ld%�����/����x"�!�`�H�zֈ�%������"������7:���,�$ꨥ�u��6!'^��}r]�d���J�8jρw���sNt)hւ�8~>�p���UF:u�L������
�Dy����
�# ����˒�h<z]���j�V�*~�n�(ǌ�hƢ�@BJ����|Fj���GL����1�1��m{��t���\����E> �D#�j1������1MR�Q����ъ$�BV���0�~q�����w߽����ZG�M��F��`xZ�/[dD�@���*7��E�+�~��}�'~ghވ<�-�H�I2n�%�!���<�y�13�?�9�HcCA t���yX�kj)�.,:��خ\�e�kO�ﺄ�G��(�
&0�k�)��y�I ��C�1}�?0'1�s	AU?�Z��m�w�bZ�����cR����e��O$��"Ðd���^��Ł{wЂ͕ex�� �UJ6�b "����6��#�NA_�Cs�D��ǆ��)����� �R�7�j��>;�l�O8����$7^�%֏Xb,@H��ոN�>��aN� �n������&�v������5"�����]QӋ ߗi���6�@d��'.y���z.�5� �s�jj.��=�����ʄ�D߸��Y�yI�s�+>�r!r���AK�;�� �V��f�� �P�NC|9Y-(��p��N��%�6��u<�S�g���z����H��4��G|������9���F���͓�sۇ��f���n
��ⲻp�F�k#����t1�KE����$E���Tl��c�������X́�dm��h~>��cM�^-i}�x�D�%��#��\t1�ŻDd����yW����z/[�t�Bx�:��Ed�Y��c7?��x;i��6�p�E��`��J�u�����uU
�o6�5��SO `���pr�Q�3s�Z���e��E�9����m���^5�^3ҁ�]�.���/�m/��3��gJ��H����-�[�"EH���z��B~�U�:y�����dm+E�%�`���H�̾�c�Vǲ��Q���{�����O�S�4�)��Y���8��
���=G�{Qx�9j6,2.Z�mg�ʖD�����H�Ѧ��ŵŬa&j5�|��H��������1�+Se�c�E�U�b�O����4�?#:�1�M�*����! 3�^����ؒE^�cZϑ,���k�	�~N��J�#�t�rRj��UG�H�Cm��q��b�(OS��g�fV
O����h{�tȨ�r{��97�����ՙ��>d��
��4d��������LXdק.zn��䡷Ae�bO�<Up���{���ZR#D=.<$�m%˨x�b����D�U�}A�t��*�:;�g&��8��c+ʋR�7���\���By
U�D��`&yo�������Y;�k־�:��.R�_Em�ۙ*9�"�L�"h2��@�J
��\�x��5	�G-�WJ�k�k��i���S�s�	U�&���Ҍ�ͩ,�WDBk~�̯�u\%]a���o\��=d�Tr���� �wI��SIu��aݮ0׆�����fh3�ۼڕT��F�7^c�8�3�Dn����	y�>����:ُ�mˉYxg��A��r/�cA,NA��Oxǽ�%o�ދ��Y�g��tl�c��{��l�؍��2�X[�m5�N�/e���N��6\�A�@Ef��}2 �ǐ���:O�>��G�?���Ślh�YA��,���oz:f~��Ǔ@z@��A�g��X��F81��S7�$9ct�k\o.H��h�b���ќo mnܔ
}��[GZ
g����<�
9��4CR������y�^�c �eRx��������v��k� � DTv�Ba=9X��s�Z��2Z��� ��m����U�͝�+��?lj)E��ا�
����e�O�#.ڡB�I�}z��T��1!��ce������DAWk[e�x&> �U��!���gq�{EZ�� G�X,}M=Tf��|�n)�JS)u�j�Ș+���;�q��ZTD%.DN�p�':�U4�����L[��$��GoIQ8;ii$�r[��T��ւS�L����+�ًb9����T�ZI��;�Y�o#wFZ��H���JN������91��Q�dp���G���N��yI��&WPP�rL�r�l�d=���  ��������cIV�B�;α���a��#y��ۍ�N��^'߱�Noat�Zi���D���K&�|Ɩ(ߗiKHxAT~�ѫ`�=@�Ҟ�=�����p$p[�51[�w���1�nAwH�TRw�x{��[
b�Vl[�o��g�q榸����_*a���k��bjce��
g�NY��)�12Bǥ��ǍĽ�KE��AC�V���'}��������g�=-���hTQ@�{�a�K���h�(jC<~�1�����jm ��4c\�l�3_�� p~P�	�Y^�b߂��Cw����R!���+��k�b�t� 	��~6�կX=�n1����!
l	ą�:m�r�9��Zq~��	�7�n�����ခg�r���bh�Vf�X|��
��j�[������e�b��2(����g@M��]֭��Y�J��v�,eJM��a������?Q���@a~�R�py�uX]���ԇt��?�ϴhѓ*�#���������Y��Щi�>�HY�T}�|�,9��V�p-5z;���'�X̂��h�N�Uz�9�l��X�u�.��qLo�P�;�W߁~��8�ekpgTo���"�S�䷗)O�4�E���R������gޫ�����t��+�ɨ���e���̓�{���>��ڂ?�?�+/�ʟ8/�I�ҠL���QʸPJ�39|�S��^b�"�OD��zA�%\Kv�1���U�Rm
�/ڨ�����ډ��sO��A�ꝯI!>��� �¶�T���eHj{��eq��e`���z�6��m���A��s��/2\��D�o�ׇ�y��u@<�h�~��s3$�ċ���Sa��\����qW,��"j$K� �e��xMż�X3bAM�ڪA6Ƣ����]N&(��@�r��GY�s.F[{��3h�y_����$BԫG�i��#��%�5���8��g�A^.KS���M�����^sS�ۻ+���<}�^�MQ}L
S�*�!��zD��67�6��i6�ɟĔ��k��4t�#�T�Ti��pD� I��; �2�MC2��)2�ɻ,+�)}��;�+�*�炵�o��6$-��<t��?H_~G��<��h��r"]�l(~B<�Y���# GD�s�pYoE� t���H������X���� �����G�ʸ�;�$�_����
5K����	����f?���!/3)��zUQ�M�"�rMv	���q�N;q�`E�Q���6f����^ֿt�L����x����`{?9�@�1}q�h������?-	 ��o~����sB���jS+f<�3���6!��K��u�o����Js��Me�ss��+n2VK	~�#��	⇋
Y� :�R�5���V�Ь���τ���9$��j:~�ŝ�'3Xh�<wS��ÑAE�;�;^jc����y�u&A	&v�Q\�PsP��?5� {��5�j3��g����
Pj�Jy�!M���j����)�<H��}9	c�'�U�1z@��gz�L���������`�"���uNM㮮�O �_J�1i�:*�]�40����7����B�x���I�WY�@����������%x%ˠ���4:��������>��Z�Z���@e�훪tU����V�c*��/5�_��d��0�m"mE���|{L�#J!T��F�S��iM�Kۣ�	��n�8��9����B����b���0��])�$��E#�e�D�ةs����إ30�h���]O���7f ^FBo�l��N"2%�QJxQUuN�<s|�HcQ���wP�e�^���fb�x����f� 3���� �Y����`æuIfq�&��f�(�L=:4��(�f+��#$ô��a+.D�m�&P8��0@8Oc��(�M'��-��cN'��� \9�6G�zf��pT��������4�L���^xד����ε3B���ŋ^�#I�G��5�^��,����N��z�,�7�erN��%���ʡ���O��̾�M�l�o�X�Щ��Y��|z`;\�/w��MwR摆{�@O�`˘lq9x�қ3�t?)��0K���9�E��&�P�,��`��i�ҡlQ-�/�6�D@����f[�H^x���|oF��ɾ��l���M�������H-�p��C�YBj�R��j�Jl���j�6�1׻�� ����yĵ�h d�.�?D+�&�d�J9Ѭɽ剄v�-� �e�i�>/�_9[X�l����6$X�Ym=Br筇	)��l�U�j�)@�����j�Ǆ�b���>�KO�LZf����¨b�]��+��X��/B
�0����"c6����XyM���x�'�a�,���iْu���H�D�����ʟP`z�uy�^�mN��>��k;o�h�D���+�q~~c}�(j���b���T�;�g��;�-��Z*y�O2	������M~F׾��Q����Rg�ū��¬���̩�}��/8��V��7�ݓ�o�q��F՛�����4�Go9�@�TӴ�z��`�+�&L�6�%��LR�'u�2�u���]1��H�P8$�iԅ����2Uј�,AW���l3�gFv��+T�߭k�uy��ٯ���`IyE�⪝�AS���	�^ɺ��I�n��m3v;�������N_�뗲�a�j�Ѵ�w�����:B�h �'����	/qF��A/D���`kG� � ����t$kڭLu���.�q����At9g!�	��M�~�a����A��"�G�B���
0��b3���~=ƮK��W�Y�P����b �r��Gȴ�mJ6vJa��"tt	��e�0�ʜ��xZ��h�H��2�%`"W�'H[��ջ:���P��Y�Ar�+k��)Bz���Z��p��.p��X3��t�B��n��Tn�TP������) G�O����Lm#U�ic�n��؈bk��\"����0��M�5�x?�����l�����c�����������Qg���a���`=�n�/~P��O�ebE�Ċr�* QЃ�9��}k��̨�^,�PmM���<��-�Q������ے�
-TJ	��U�A7+d@E0&�F��5"��I��VI`�A�<�]=`Ҧ���5|sdo�AZ���x�?+��PH�&Fv-��EM��Y�̛2B}qNE%��ae��:�V�-�	AE��+��l����^kЦ��6X�Ի&�� �q�8���$���O����!��Pc�F��.����f`��D�o4�fZ��>x_gEF`�=fg(+������GH���&�ni�;�$�޵�Z���?d����Ils���xV��Q���eX��k����Nu���z�	�?C��UT����b_�Up5X�=�yIM��E��<F�6�'�N��R�-;���9��۴�#�~��Զ}L�Җ�.e+�Y-���y���3�l�_�U�1sS�D�;S.��;yi�,��U��}D��o�G���Z�3m���@�r�~=���wcj۞t�����hC]���ϔ�Gx}=���F��E1HA�M��j�dBz@��xS��/t�4��â~}��BE�/�O�ĵ[��&Rmy[(� ��q2�Q�8�=}�/.J�9h��2�2�$��g �\J']�0��ȍ���&����,>!g��vXX�>k�75�M�9�)��6�mͲ~%N�ٸ
x�]�[�L�=�'���}h���'*)�8j5����zȖ�7;vu�4^<I@t��p��CE��A�o���\dy_� ���~�\�fc\����Ɠ���_�D�?�}$��o!ƃ+��Ӻ'�3<��ׁU�o��G�~�F\�ƳQ�U'#���2;	���F'y�Ǥ7Ų-� 2"m������-�mMl���gQ���
)��� oGt	B&�3e�=T?���h��gWɖq&�f)E�M#g4��**���(�jg∯�����8r��Q�6�����p�����s��j��R�7oM)P��0�zk
'��Ź�����f��7!6g�-�8o~�4��܂]�2Y�c����������8��t6-/���℡���t'���~o]>���F)���n���˼fL����<XZ���)u��Dm]P,z���(�vW��i�I��4�`��O�[y�ڦVWu5RX5��wLx�[Rݷ�Y]����`o�$�=z�6>#��L�1&�T�U���G�0�t�o,��z� p��֢�;EZ�Mgc�Y�r��2�ȡ����G�d��Q�pO@�+B���Y~%�9�+% �)�S�<��O�"6�{�ټ��ʍ_`���i��ɱoD1r7�9F$\�:OFh��E,;+�Jh�R%�O?%u���YkO?�(�g�}�\f*�aV�툛���X\�����Yϸ�t-ك9X>U�.�VD��V�n��ٷ�*�7[��NZ�_�|������ �*�'�S%�`�S�*^��RW-�#l�BjX�����F�l�^8�;�~�RdnF��^ܖ��{8�(pf�D�i���hW��8�(8�O�4,�Y��3�u�f�S�ӣ�Z�a%�$q����LLW���.H���/g&����(^��pH�3�x�49�R�3��ͨ��)�lf2�8�?�Zwk�'�~�# ���C���He �PH��>b׮=)��9`[[�o���_v�"TH�5}��n3��-�F/n>0�mH�
�T��uh�o�_n�NB�K����F�P8Gv������8K��Z#�����i?��9Q�;Mo���QR�J����\В[�˄+H�d#��Fl�/��,l�-��l�8Z�̮%%'���f8��U�97w'���&���pdL(+>�0@<��#HMs !9<�2:�w��燏�����ߐ<8|1O�O��T�����x.-4;5��yk�q�L9���v��/Q���D�� 牴;Н�2�Y�����:����RW�%�5�Ah�N��MFezI�\��F� ޱ��:M#R[�@}n��W�J��1��vV�C���Go"��]ja�miX�r�֐����/3D���Ap�#��Z#n�~�X`������Z0u$Ӣc0I���$��3���a�ѻ�#�N�@��ĺ ��� �h߽ty�K���lj�0�n:���ZY��1�/N-r��� �A��Ae������`�Zf�zD؎CY�Ǌ� �I�����E�+4��$��`O��C������yQ�:w9PD�-A*����Қq�y��#N6�����-h1��	ϑ]]YE�#����B��:��2<��9i�u�e��̥t-�vOz��k�ZhdN~gy��n�͵]i�
\.���Q �kcxK�:F�3FJ���R��\�-���ƭ���H߉�E�ߒ���dI$���#Zق(ld�h���H\vY'����n����;��Q�����F!��`���x�UaI��gܖ�)��b�3j�7y5�-U�i�H�g��?�������`V�'��H���|����v�b�.�^PS��\F0Yo�O>Q=��XwkKzo7A���˼!9g"�c܁F�o�խ���w�bR�Eҙ#׻��t�tV�7T.MK+���B4V���Ȓ@�I4%���N��#{~:o�������uwD�N
 sI�<�;�R��*y|hX�z�mԼ�(�������ԣ
K��v�M���ԉ�HL��2]�Q��j��G�3��2�ʆ�����+й�'�8������<�} s+DPg�}�O���n���
d�^��1P�_%d�j����Wk!_1��B$��o��R�y�SP�3]�/���l7c��Z3\�əy���(��dy��7�|�����"�XC�93������I�'�J~��!Tz����(���JO��h@x��,'ZA���ȸ�4�D�1!�M���t��A��dwcbM�O�[�-+��D��O	�(��9(h��7w�ǃ!K��ç�o�'�h߹��(kՇG�_�j�9<��7��R��,��Mu-�ݘgYb�`��˿'�=3"*禩�{8�a�'o/u^yL����~���E�x[�V��&s�K`��+�Ч�H��K"W]�k��Ÿ�Ls�$3�^u��{f���A?�;>/$y2�S]��RD!ܭf��:=6^��Ď>�Nm��Xd��%�V s���,�7��^域�_��'rt ��xV����أ���;�4Jߐb�|e ~�~��M06(�pk,�Rv׊��O5��F�_{��$�T����M�bN4,T�<A��$.`���76֞����Y��]-�A/2���
$��W_+m�HϱVsF��@��0uFC2�W��3����"5�9�X��M��������)	>MGT�ՄV�8L������i���E��ΥK�`��0�+��t�$;����yr��c;E]e�4ۍc�fI���~m�q��zn854��>�s�I鱡vZd�kld�b�W0�JQ�_^$J�3{Ԉ`ఱ�¿3��ҟZ"���@�����@�M��	?6�AKb������	����l���I�(܁t���y1m	Ю0+��{��u�PY�0��&��{�B�)��{�T8�BS�k���/b��f�10�J�g��Y��q�iD�h�@�D�V.�Ҹ�q �	��LX3!�(%�9Xk�{/U7 ��5|)�d�!��Ɯp���PZꠒa竑,��g-��m�r),�@��rU���ZøY�'ADי`K��0�٠z���A�������n���8.S����JM�˱�z�rp�ai�$���aL1�x�]�{@e��/-�C���9��u��ꙣ*���w�������-uJj����ݠ������{���m�.�G�Yo��|�*�*N&��G�S��� Kc�&��!9qA��8�-s�;޽���� t(�&��Q��+�	R}�
����5���7��SغՂ��W�i9�ԣ{a&�Km�I��!q>��1{�
b�v�8���/�߳���.�����8��j����پ�͢����"iz�ar|�JWz���dA��"�&)w���7rY�u���-���c;��q�I\����i	��j���3D�*�kF��L�XG�
.q�F�R�^�(h�3Ϫ�*�	�"<�X���ʝ�*��@�9�k�bK[�gn;��,�i�3�"���Q5 w�+���CJ�]��^�{��E3Yq��xD�-o���(���9��l����Yџi"��pҪ~��7]��m�j1	���xS`�~K�:����F@8~ +�w�CR�ø�{�0%ԁ	h0KG���F��KKS�@��L�]o$�r]m��9�/��-%_����i��R~�����j�!���rc�Q�᛻{X�'��IZU.j�!(9c�Y����m,�S+qŰ��1�HW|M&Kü5�im2��sV���6~�8Ł��t�����V�
��3w��Ýt�N����U&���&���f�.y!\z^^q_:`<�[�yqVb^ͫ���r���:EV�cu[F4�ދ�AY�n��77���'�
�����~UF������LeX�]��$ڜ*w�3|M��fL �~\�kK/��тm#���
�kOgi�q�Hb�5T�F �|��F��!쎝n�/�|����3��J|�Qb�s+�Yk)2����c�B�I���8�l� �p� ���ve�9o�_T�xm(O����Q�?��c�gR^�H ��,�"xOZ(,�/�ؖ�K�3 �o�2�G�j���}��9��,��k�q�Y��*gx)E���#�o�J�6@JmX��?l%N�zF�pLxv��n�b��P��
o�7�9�̷;�'��2컦X����=-lI��4����EO�M0�w3@��Z0ԧ�Z~�N <lF�i�VoK?����s��>�g�*�L�����s�zx-*ޑ�-G	��h��,;U���$��䓀T��J"�~�82�8�;�S��+�)
jF7%d�w���4�6�6�gefq"4�_�������R��α�{�O�� )�m�37�:���J,�EKH���W�g���0D6ˋr�+I+�����&Ea�
˱��~�� ���I ��Iu<��i1x���K�ڍN��7�~�BP����p���h�_���8�V��C�����p����{.}$��o[66��R�)�� �%�#nq�����T�V�3,:V&݈m��o�k��ԯN�]P,�O�Oش:�]]|���0Ώm�R��_�J���J z^T/ ��Uf�AH$��xx���zV�"Iy��w�g)�n��<K)�%;ʸ�ЖAE�#�cM��'��%|���ُ�d�O`)���#�2�5Jl��>*�#���������b#��)�}ypf�I��~���sT����s97�f-��"��H����S��:�+;q��3��Պ��\٧	к�fg0HۑbP�!/���G�ڔ5P�����P����.���Z��[��۱��ږ��c�֨�.��m� �3;�'�8<�M'�(�9����_[����MIq�v�!��gcl��Y��ܧ�!����@�˩���A��CYa�Mͪ�����d����3�
Je����F2�\���
��u/F��i�,f	���γ�Iw�Nc��F>A�t���H?h��x`��]�!����mt$+[��/������s���*8��&�ϨL��ŰV���$O��G�|���hY�"e7LԦJ��{���F9��)��'i�Ԫvs�h�{���{����4��:�S*�gt�&E���j*�N0��-+i���d� RL�-��������<�w鰺H�۾ھh͢�O�;N�RH�����)�r�.v�Lh�O)� ���F�t�P
�a���'�E��?�Gn�[<�|)�ΎdD��=
�q�c�'���D��g��i�N�����b�@�d{�����]YIha^3O�8:��",	�X�|(�z!�7�$Y� �<�^/��|�ƀf�#:%9�zk�������4����t��[�w�T	h`�<(�uw��K�*FTס�R�m�B���Su>��̵������Z��y��^b�����j'���"�{W��������lay�ݵ;Hǎ�r���I��ꚫ�z��!�h�SPp�Ծ��(%P�4u�"�eax-�0Y�e���};�}���aw��؍s�P�p7v/�)U?��� 4����(�� �KBhᛁ�}����kh�C��Y��b�Ȟ-��h�V���k��<1�F$�hZ��8�k�Eɹ���]����U�a�H��+�X�����Z�FGۅG3��_L찛����Mo[���=��*�[�]��_y�����|ljr->S��\���Y+�!�2�p�ج�⩻��k?9
p/\�MP硟wG�1
�ޓ��>d��R�&$N(�l8���{ߥ	-ӵq�ε47֋@/��y����OM��U�	i��S���7O�z�؈�����E����
U�.�BSr8�:�|f7E�'�ʩ�149J�=Y��rj�m�� �lE/n"<���T)z��/[(��fc�gn|Lf!���bH���{N���ν@[z�!Ꙫ^I+f��xI�x��ߤ�*|
G��wDCl��=7d�I�����(:�FX���T��42�{U�T+d�|N~M����g�~Æg;X<jI� �l��g��_H��l�^HI�&�\[8C⫔e�����pJ~؜�PŎ �LΥ8v�,��J��^����ܱ�6��9�|����b���� ?�M����wY�k-�O+�6���̗��T��(.��Y�_�%����.��/~I/��u[�}��o��m�Ąu��F�?�'/�JY]E���V�F�Bu�K{�=%̬�J��G[PoA�0���S�{���+�B~aSue�G���&�����+�G{�C���(��Ar���x��m4��\�̛ٗ�.����vG�e�mQ�{���%2>�B�&�*����n/��p�����eG����/
�<��D�����A4�"(�Rd\�|p���{��|K����1�b�
Hn%��BI�Cq~%r\����=��uI=:}�)�����e��ظ�@n9�6��LښJ��˼��+
�C��]��wu��#)��ɪl-I}(%�C|!�TԹ�N�a�oh��[�]�J���u_�JF�U����h�BDk��:9��ٌc-ѫAB=�n�>�GՂ-n�,�a��6��{c�:�=xn��[�)Uh��N0K�4A�19�6��ie*T���wv<���hq��E�VR�����D2�!l`8�ʪ���\ވI���GLہ��qv�	�������O<-d	wy�H����;P��1����zrˋ2��IkN8.���{o vFF��TSF�o
���yy)ƽƼD���+�T���� �Q��Մ����F���+�Z?�2-#�L��N�*髀9Yg��6�N����N^W	�i�N3%���f�8Vx��y]�J��	r� k�/~�zr:"�4f�����=���g��իۺ��{MK�>���~Ũ��ǟC��2"L��{�?C[�l�5���ƈu �7}i!�E9}�d�:����c-�V�?�2�`�X]�C�\��tD%�/�g��{e����Y��;�L�� ���w��z�����t�H���ƞ܋�d��N��n�T�X$s#tCx�/I������	ϝ3�M������t���\��O�����@J��A�*	�&���S���F�:�{�v�R�#�y.^e�
~~�x����&�/��y���6�Bs�=�]2ai9���W`���ܹ�ϙ���ۅ��9X����&�sdJF��S.
���)P%�2Ӽմ��}k���+�or7D��t�;�����B}L�u|��g!�B�#���[�$�c����Ƶ,�F�QY�H�9� ���{?ٚ�Y���������\w��;�%T9X�7Ygf{��+	�n[��.�$����~ִ|b����(	��9P��	'���-���Mf�(�KN�����Nރ��Z�������쉨q��fBy���٧�+e�ZV�,�����qE7��(L�4�x����F����})9�\�&�����Dq8��2�H��iɵ��^�n�Q�z &�P_��3*��S��1�I�ۣ�A�#�/��j�:a����׽�Jf�ְ){>���O�C��X��Bu1�(�A���	�DY�/�����k������.�<�T]Pe}���P�e�s�gRe���!O�-R�~k�l��ե��-�>tο���_�t��@�W���0=��"�W03�rK�_��[v�l���"1G�z�-n���_��g�:���8F��H�霪R�0\fН4	tB5�!uw�ˡ�5|f��S����=�D9��c�/\��S
1���Wt�o�*�E��ЕS=��?i�'f-�q��p�a(�@��C�����U��v�N�獯�Yޠf��o>���a��O�E�S�	b�d�[�:��e�&0��;^)�����Y�2���:��g!����;&����q�I����4ਘb�d�KxWB�r"���D6�e5N�;	ƣ��|�/?�MY��/}fy�w`�E��#�����vd��x���SDx�4���I]q�޶ݜ輛��i|Q4,�����ޡj���Ue=�ϭ�#Y��`��)$%
���Ե��r0�Ϋ�|��L�p	N��8ssjd�`�\����i����P4�1z��67��,��/S��r{/9fH8`�F���R��l��8��U��TՄ �	�=��IP����q���mݎn�&ҏ2��	R�EvZ=��)���׭|�B�<�)2aиU�)�U��'{�h�����W��R2!vJG%�fYE}�j���\ �c=҈�MM��� G����u�b�'t�X�%��KT5o"<��R��շ�R�j(�&��x����m�6���p�i��8�����B��-�O\T�%����t�
,�7��r��:�C�~c�
k׺��q���8[{^6{,���N��� 1��ܳ+m�Z�?O/sVgʭ��+/�������h}#�i�@�R����ՠ��g�I6曈jt�h�߀��
����]|opp��*��i	}�^~l��Է�t 4��w�Kqt��V���O���>�@�b��t�g �1W�-Ad���� ʾ�X.#I��Q�Q��N��;pp����v��&H .`�!�Ot#�m>��C�)J�xvǓ���*i.�� :��R��С[��#��x5�R5�����j?n)XhP)�A��D3�����ث/~`l�O�0��������sKd:k��2;�EyAY�b%J�\�+�Jx��Ug�6�@���i;�B�?#�z{?t�j���h�Χ~���K?|kBA}�@PP���Lξ�=��~	ӗpm��_�h�n�>��#���dF@n���H���/���d	��
��T������@���m��e?V��y�}���\�0��E"l���]�0�*��W!��R_ޏ,�N���V��[��@�� Ho���b��:�zҹP�Xv����=vƖ	����Η.ø�s�������Zjԕ��9�bj���#ƙ}�DN<����X�
.�c?T�9@��9��;ɵ��v-��ҫ�ݚ���=TG��_��uŮ�9�I<�n2��f��' !F�tf����_\�j�It_�fp��M���՘��|�l�U���� u���%�QV����|S�[�)�Q�W�
uX���D��;���hު��Ɗ��곕�a���ʔ!R�9feL [�< ʊ����xHP�Q�Mj����E~�.�l4��-3:���/�s`�q D;�_S�&H_�Zs�j�~�~����Ȓ�4Q*p�;�s�$�XKB>�S"g��r���S�f�Km�ϝ�X!6f�N�?�LV���ofg��T�v?�֜iA+�H���|��LfJ�<G<B
ӊ?H&��Mƶ
��w�:��n>�4�<�0ۭ�2�"-�T��]�YjP���������=}
��H#z��~���)yGp��Fr~�ܹIUV����pW�ѝU���:�nQ�L����k�w(�)ȭ:=7����Ibk4�C�,w���_�)C��W:�(IEL���	�R�*c\����!w���X��M���WEÓ���g�'x[\V���3�� ��,s�B���]�JKyα�.�m9�nZQ�u=������a
NJ�`m�)��,5�Ws0=�8�j@왓�q^�s%K.��/�V^��|^�
 ��`�yc�۞ �qQC�/�l�-�\�dqr�%8�1�e`�,��,���b.{̮E�׆�W�yr�<@�B��9S�%ˈT��H�=&�)���W<8��,_A;:���G�DuoٹV��nU��kj��ߺ�Z�DNW�X���T��rI��ݩxb��/�&Q_�@��t�8��vm������<��iGF���k�4��y��]DM^륑��h��J�@����Rk:cSz�3L�P�!�;A)r������߽�d�Ql	ˡeg��193~��΋|����"��e����
�*�j� -
"�0�y+m6}���F.\����4<����r�#/��J���wN�r��cR���Gp���<�1��r�k�����w�f�`�zM9�,��u�o���:'D��~X���p�kh08$)�ԴkVD� ���� 5P��Xg��Q"���̾����Q�u�F�v)�-��+q�m� 4�1k�0��k�W��}7���5���������Y���rF�2H�(t����Y��{ @���
��p��ziѣO�ո�Ht
�S�Zd��,�
{uN�����)I����0�to;�L4 ��w�6�j][;Sq1�� ��^���#
�/����9B���\͐sDL1yZa���-����@��ł�R�W�=UCÁ�{��B�����o�YJ�S6��Q_���z���4랓���P}�X��4��j�N�R��rT bH�b��2�`0�b��(�w�F�U|np�'���1}$�zl>��{��~����4:�rȝ��)@�G`��o����8�-���秪ңH��i��C-�654�}v��=k�K���A���re�IC~��O:Qj�ߕ������(�@>���ҿ-l`��VnE+���5�$/������FK��/��E����KKӫ�ۜ'��r{��iW;@��黭o0�;��cѐq��S��ｹ�";����s��W�8��_7�K�&��U��0�h������d��v_�M��2k��{�{9|c����d<�4��Kf�4x�$Z������b���������YFQHm��i�a�<�mۆw�o`�I�.�,�q�O|u��5�]�J��&H�P�l����n�I�]b�<��l��_3��!d
�8�� ���
�B9��^����}x�_0�o������fϖѧ/�j�O9 0M4����;D�E\W͊�%@��\��N�\6���$�5N���uQ�h⴫=��n�{9�`��X�b�,O�T��taLlƃ����cܚ�,��}�լ���"c�<�ܘ�e�n~e�E;p)�9W�+�O�Z�����-c��_�9�O��j]��<��x�qm�CZ�9J&�;P0x`�`�Z���/��TUg/�#:Pl��P{k�!�[��Sτm���JF�{�)]�Ԗ�D��3k�}	�E�>I���琸n���ޤA�S��XB�H&:(Z��zΙK2Z�q�ꞡ"l0G��қ�f,�rɸ` �����|
�e���0�д{|Xu��P�P�gצ�ާ�����яf?�u�W6�m��
ߒL.G�������ڛ6
�����8�nx1P��A�ꃷԠPB	,:��;�֚;����A�������V�v{�B.��,��$ը���:(h�{�c��4+��٘�� ��� V�J�Kv-�\{(�g�`,�<n%?����h���<�o�;�Y�5A���WXs ���rVR;A ��Ӯ��(���E>�.sC��o�9~��ɽ	�����uD��DA���᧧���W����LÄ��zz��21�@o2�.��E��S�����-��$dtI�H��I��pϳ:����N���R~>�oˢt�����]ﴞ�ŵ�K	x�%��=��Nx��7�k���o$��ĭLj���B���e�VO�*�2�W�%��I������D۵�Шߘ<M#��c��I1d��Y����?��A�؛�3jx���8��\��� =�=Ť�x^j
������̩�.�-������q�A�HU=|�FY]zǶ�#��ૠ1X��7�N��r";��5����3��e(v&\��	�0@z�Iz��7��~;������Ց�+ ܨiH��&:���c���E6�ɡE!x���s�� \��46���~� G�É˱���BYqr�:zlF?�������������9��I�@={6�2Z+'e�ؔ�v;��3ƴ�Q^ ���A��I����	�c�D	iޔ�Y�y��,.~A�%����:������<�5���o�&m��/���\�Aǌ"ף�?�n6�r�!�~�6��ד=0�c����E��p�Cb�Fw�����ʲ����_�.�я�{�h�p��AÓ>*���:VR\D�m��H��َK�cxE� �<�#������=���R���D��9B2Z���RK7B	�;o�Gr���n̐�f���)��3�R`f����E@J���XGz�ߟ�n�8p/ӱ�u��I4���������vI��5���� ���@�ɕ�� Mr#��y�_`2���%�f��(��G���n���rҒ���%����;J�q�qi�((��a"ؑ*�]o,F�[)��|�ҊU�V-���<fPQ;�ɖ������|��=�v7XE�e	�����O�ۉ����g�?;���'����+����!_��1�ܬ۩n�ioxa8�&ɸ�.�� ���cj�8;�r�7��f/��U��S�Z���I����Ur�G��Dh�t���[j504�&���K��*�pJ��:8wGWy�M��֭X�n��E�:At�½e��ģ�'ݏ�K<�f=�>��躗q5��bW�[Ք�u����(wT�E���a���Ѥw���|�����k ���~ʅ�^?s���r�)1�
����k���]0��J����2���b������������g3�T��ǽA�6>cv�D����n� ��㽎rV~'�"�HjG�%�Y�6�O�ƥfiv�����)h��YܺX����(V9i�ψA�1�[�<�\�ں)� �#WH^��}<�2���k~�-0�/R`8(4����9>j�Ԛ?n'��O���N#h��Ӗr�+����<i������F9��&�=Z��"�g=d��GX�U;��}�ڜH��|���(��H^[\��I�Be��I;�`��o�z�:��N�q����m��S�Zؖ'�-�4gYS���n��[RH��f��5��9�����Ѹi>���1�-(\%z2y���_���*�H��	�����CE+4�i��u��h����:Hث7[��r�N��������u�a��j�JU4���P��lH''������X5X�M�g�Scle��'1>���5F�F\��l����ZYl�7�C� V���X��v ��:#��&�K�-q}��b�zͦ�_EL�f:�����
<X�]��ѣ%�������$q�yK�e
0�f��φ����	���3�{G�E�JD|;���RĐ~R�;���L��Y*Ϟ�̜��S���.)�t�p��0?Wv6%��+J�;2 ��@�¦�g�!Lpƌ�R4p`�Ld�{��T4sU�ͮ�)nC�B��m`�  Ce�T½�V��-��% ��='N<w�d�4A��)@icS�Dh�wA�K�!����$�g+Xɫ�!?�8�9>��02�[	�C 	�ߊ��36]Q��M?	�mL-�"��`�Ap������D�'���B�k,���Sg��ODA�����R��=կ8�d����3��[2߭-�-6��a3e�;Q��]iK���h��f��TV����(�u :�-G]3��T�.�ęXq�w� ��)�{��i�ng�[ߏ��*��:w�@뷃�͟���O\H�ڔ�!g^���>����"L��Ǜt�f�5� �K����#�fe�ؔ�֩%��/v�Z!ԅ ��o;��1'�ъ�:���h4�~�X��v ��P|�{[������u�^���7�Xէˣ������/���X�#V��q�H]l�^�"�و�40+7���A}�g�1�(��L���j����K��J�S��8S(D94o(�.���K�S��bS�!��V� ڪ�������d����&xڏv��t����Ry���<G:��D5I��G�0]}�I6Ӣ�W��tL�jm��J�`�S����g�@1U+�ԋ�*z���5vD�PDc`��*=��2�2�&�`�T����@�0j��r=�����棧~��lW��{���w)o���Q�{���c����^��3O���p�> �(��]AXC�QΈ��b��*��̨P˰̋m�F d�l��j�_t=�o�\b`�e�����u���Csd��+��5��3T\����w\��wE�^6��=m]F7�Y��Z5�뷝Q����1�i=��&RT��-ԕ�$�8V|�0�ɐQ����Y��'}�$5D��ӾE��S��]�py�4UL���Qc��	f�E��+�P8�eZ�G�?n�G�Zp0Y�P��+m-M,�f�2�g޻p����
)f��\�>1�>kbɳ�?��V8��	�N�@
���s�Ż%#�-���f���ԑ�-C��H8�/
�6��s �fK��Ђ��q}�5,_r ��P8`�׹��2r~����&�+W���t�5�KBBˤ2�#F�a	�
������B;����V)r�a�'��w�t�3X18�f27��X��U���_̋p�����4��,u�<=�-��z���D�R#;�6w�̈́�ݝ��	�G���e���8|�d�Q�B���E�^����K��Ԇ�6��s�U�vո��K<x���︯2g3�d}��2� QƗ�8Ψ������A��5���G���J�c#��tߟ��R;&�ţ�W��i]�Epv�c�w��H����4�OէPC*w����#��|���H��_�y�
��ȕw/��jq�a�E@�[�j<di}:�i��E]W��^�t��	U�^��2��}��O��αV�Z��[�f�?/�w� H��O�|�5zTu���8Y��*����fX�)=ÑX�RE�G�F?\M�K��^X��- ��D<�6z�i��NX��r��A��+�s��GҸ7D[D�Ϗ�Ò��:3u��buĎfqơ�P�H�M���)��H��>;�PR���wC�*�ޙ�K�t���{��ۍ���$�m@֓�_��f鉩���_������ƴ���09�}g}�wg��E=m]�}���$LV4Dv5�b*D}�J*�Y�����_+�Bt%�Q��J.=팬ZF��W�CXV~��"P��Pu* ����� #�Y��%SJ�0�?K<�-�y���{M�����oJ�0�ʁ�����t+���S*�l��S�]�ټ	젚T�7G��6��9�ڮ%�(�ܿMS����DB��^X�]?�o�̳��T'ѴOq���Er��`^������3�U�r��-UyK��4�]��>���� b�i/�(���m�-��-�VM��|t+�z��4��G\�j!�Zx��� 	�E4�)z��0y3|'���"[���=�@��%Yr�	
�g��dV�Y�U@x"�� Ļ�"�o�˰7 �`i�w�4ے�98e4{I��b�%�iH��'e��L;�#�m/�2��
E�--�̝v�]��IB�M�}AZ_�-m�u��PM�Ԓ+d՟h?;��{D�u�X�E�"�w<h{�������̤�n+�ڑc���-��^���� I�^��*U"�I�ٕ�{ÁB�"�3p2%i!ߒ�J:1�L;�Ք������{'p�^	U��B�78M�&�x�3�ۦ�uNg�ݘ�ʊ�T�R%_��5��P��)EB�X�M�%�)1��}/y�F��q��Tu��e��5�tn�9��VZ�N�#JP��؜�g��$ؒ6��iq��P_\����\`ʅ@�}B�̝��$x��l�sZ�Ĥ.,���؀���b��i4��0��}h�v*L|���Z# 5��x�
�#�yMV�~�qۘ�e2(���T6~F0������97&�0	fڋ��	�Bז޹����y���P�:�Rq��ë�����iKK4$\D���EU��Ü��F?�1�ab��/zvR�"��f���l�$Vz��O[V�+��p.�Z�+�u�=�sMi�<Qf�;v{r�N���nCƸ����b��������'�X�����c���w�76ů��Q��P����� {�;Q�
<P�ìW�ǒ����4Z�":�?��"y��X[�vh��\�^�t����a�Ї���"����E9��ՠt�k�x�SE1����!	9��-F�7S������-��	=O�\�_���r�Ti9�)c�̌���=+��W胾��_Qщh�}�'���P��)$�;��ZV{3Zy�j��y������S�$������h�3<l��77���V~.ϡ)��,��(�� �|gˈ_2QrA�Ia�D�/��-��M�՚VPux1�wf�A���qu)̯wF�`~�	x<��͡Bu���=A��^G�rT��N�$;Oh�83D�y� W�I:ˆ��\s�����c#G6a��	���Gf��6LyB��1sq��R�[�XZ��Z�ʪ`�|�s�O�������5J�(��Ǿe���hb��F'AS�͆f�ۇ\2�<���w�	��������<�mw_ۡ�,䉥�hu<�t&8�
L��Gi�L5'�<������]kC�2�(�|V�U�`�ڻcS<.hZ9��Z7��9)��E
{Ç�kD�R����2)�"��V�W�W�yP��p(����;��je���`w!�t;�񢛊���U���(���-Ѿ�[�)Z��%)�f� �G�z�ǂ��%T�+	���1?������-߭�ߴbV�- I+��d�,1MxS�'��/eའ:3�y)oLz$�WS#1��#x#l�1e�+���n�9K����0T�җ�k+u�"���$����p���b�XE)3M�H�wCs�v��d�}v=,�u���Q���e�a	o=�.�I"�1��fj�Gٲ�+j|���^�!�bN�)�=��9N��xF������)Ձ̧��u������^��sU��x�Oߔ����_K0�8��� ̩ÇA�W��g�ٗ�l�e�géS�z�g ��%C��!�^��mr�?�M���2#�9�%�Ҕ����޵ެ=���0�_2,$A]�l�j/b�&sJzV�M�rOn<�8����8��95��o��N����3O�������7_Q�hz�u(I蚡���
����>݀�L����I�2&Ƕ4�͎*��36����Qo&r�ؒ��a9,B���"�8s~5�>E����p�g�S4{���M�w޶�#[�*o���ixD�jo��t0Z`�i޿O;�OSrDOx2h?�ݴ*�����}i���K�����40�Ϻ��v�^t�)>��|�T;��6N	�]K�s�5�obr����
?�(�ˊv�e������b�)��╊�F���uA�Ma���R_��dA?0c�����ٴ�θӯ�ڱ�=�pf�?ITq�
���SDI峩��ҡfh���w�il^a#�MZ���cWO��K���Ĭo-#������@���$պ����wx�2c֋���t�����f�w�1�kT�zZpm���QCH?كg�T���,)�-.� w~�ٌ�n�w����Ԏd��l��seL�H�O�D�B��< M7H��{+�ѩ�
L>��@�7�Rޝ���*�_����/^U�ɂ�|�����؆u�����ۧ�e
��m� P�+׌Ot��c�D�R>t��L;�#{A�'��F�y�����2Ƽ�t̚��֒�j�4tQ�6�E�&���R�#��RxkT�Jt������N����u@��"
���FH�<j���+N0�KA8}6uz��<�1�`$�v(Y!K들��Ez)eYG��@d��5e�7_M�$D���,p���@���Ū	!d�˻:?����K��7}��|E�-��$�rA��k*'�u���i'`�@>j��B�Q���CPE��d��`x���$�P��U�ӊ�ua���Ν���T�S!^ �����{�W�·�Cٗ�F]!*k�Ȝ�%�W�Y�<��y�HS��)�.��=��6�B5����L?y��f��?{�C5�HqC6�հɆ�T� F���3�K�a6Qq�b�Oe�]A�$n��6���ס���~ϵW�~N��;?t��o�U��
����,��y8d�і�BrZ��%r7uĳ��*{��v�M��ٳ刐!���ojy6āAΧ��������\�i���%�Sq�U��M�]�$?��O�/�4�؍Z;b���Ke+3�x�H��f{>B C���~��:�ي���,n�	���~\h����(�`���1K������Xu)4Uo3g��P~��*���(��1�N�W��ݭ\�"�M����N�&2�s��lEe�nӵ�BB�����Bk��F�"�
�q��t��,k�+�v�(��B:$�<��e�	iq~Ch�L,��IR��,�]L֙|�5�[R����r.{߸�E����}�߾	�#�����yi*�zn�-�xa-Ϝ
FQ��y2�3�nZ��	mnli��'ԁ�&T)�{���hT΂TƼ$
�U�>|y���h,mO}�J�z�~ݏg�H�W\#�Ψ��1�;	_bV�uOH�����ӗ�=M���S�v�\�?v]���$�dM1��)�D;`������� {���@b�qe�C��d6&rW"�M�f�p����$����n�1�@��"1�ֳ��u��8C%nP&��oԸm����dP�
6�GE��-|�\X�
`mƕ�4�д�D�v�{�i�Mx�`J�)e�=����3\0ՂN�
|F�#3�;	)�A��5�Ծz��p�t����ۇvP���G��㡘��Ƀ�8�"�ru����O��ʂN"��7WQ#`��K:�# ��t��7���I�4inJ�Bq1bÉ��UW���d͓�F���2iM�WRUJ~���obh ���3tH��ʜ{�S�dO�#��6�=>O{�͠.������a��G��?3��}����&�Y��z�̆&���ƪ��O�BT�>�ǉ��ɹ��%�bO?���$9]�ˤB�!exRg��m9\�!̴����e,	�3C��4���^����ZCP�3�"�a�ɏ�*R��8�
�|}�o�����w
�VX�r��!l�p��dV�$�qL�r��i�F��)�F/���+�i���E���Ԕ+GL�uT��OR�!3�8����a\ihFL�R�w���AݰR(oJ�8��,�AK`*U�:ꮞ�z�b{����M����A/��q#��1� ��ܙ�Nf��'m����ԡ:��v�W�$x�zW��⼶�n�<��%��)���<�W�*
SK�&M�ۍ�GƆ߀�f��g�\'�����^���H#{K#PO���g?��tYf�bM� �_m����T�:0�<6!�+�
c�´d]v�� eg�RM%3^�#r�<�$��@S�;!�V*�ܤ�GO;X��Ұ�?� �C��Y%H\��l?u��Oˇ<a鮌����De�X�C���Dvh��9!�;�ZS��X�! �Bs�O*��20��*ߑn�ߎց�	�[1�8c�����K��V��RP���wUX�w
���7���W�T_���%wD䓒�j~(�څ��� -��G�5̄�l��YA����#�ɋ�.��貸���e�����C3��$����j�p~�oL,��6\l ���Q�o��%gM�4�Vf�!��:�HE^��ఝ�������D	�&c�����n�Ǉ�H:�^!*�E߯� �I�E�L����I�~��e�|Q\�ൻ���$��Y�VN�;'sԙe�� �6%�j��:f��-_j~
ȩa�=�u-��4���/��|�:S�Q��poԖc��A�#�����>�]|��l/E��߀�e�v-.˪��ҡ�õ����|`���i4�dfzS��r��7�t���Q�JC�Aվ����8͍0�s/ڱ����F�����8&��i�rB����>8��i,;��rr%a�j?�ߨ F��r�<Ps�:���c�WO����sF�+yN-.�%p	��-�6�j2ľ�g=
�!�����ҮTc��>l�и?L���3t��	��C8���a|����'�]?�/�Nt�ץ+NA��ic�W�Aa�.	f4 V�H�2f��2�ג ��X�r��yP�#����-l��e�|w�6HѢ܄4���YFp��
~�p��$�T�����������VyW�g-	�m�I�0� :u�;ˤC��5V����6�'D�
~$֟X�]�d̰`T-b�7��{oZ#o�+��<]$5	Tˣi��G02^���nW�7��3�0��M���段i�3ϣ$�|���_Ͻ�� �4�#ͣY��gp> ��;�[r����hb��{����bh@?��&p�N��ˌ�P�,Pn��k��`J���[�Ȣ�[�O������.�p�[�ձ	 �p�eL��r�,�S0�(��wy���*=��i�jp���̇E��GH>GCO�A�,�/�v�<�rF�Q�.g�[T-�/U$<�g���.J��޼<vxނ�k���*��=۲ƌ���oخ�ל�Rz���{$@<���|9�bO���ʙyA�Ke+]LgT<ս|��u��S�d��U�m2}zv�Y���
��dYO  �T2T׎����Ǔ��o����S=�C"a�Y(�+6�f�T��q�l�}0�*�����Vյ�&�Y����Rɀ��g�h}p�Y��uĲ�j�B��*��s��p�C��MKꪝ�ã}���"
�<U�[��6<�.����$9������-)`�cmM��Է��;mg���#\~4���RBKMգ)a�<�����Z�_D"A���2�7<��kݠ���B�[�L>g�^&}�8���~*�M�{}~�Y���Q_�B��Hm�����uNJh0O�ڿ�W<�n�,U��5H%|�u�^��Amy�����Ի��_�����7	n�{�\t�`��V�޿����F,������}Ry_����� ���W�;cXߴr��CAB���E��?�4�͚'���!���UhN���$�9+d�(�m�k�k	��G��x�'�%`������4�07�Q��e��b%�ދ��x�1�-����\U.˹�X��q��N��p���D�5S3{[B��Q��%����ҫ�YdT �������`cXH�JpK�o��� 5Q-�%"G
X~SZ�I``(Y�� ��6oy����D)@�!���6!�~L]���4�ꃠ�|~(L��F�B�<�N"dXܡ�ߨ�5��.� eHF<���8A�F7u㢿&ìh��κX��t������åQG�wőy�nG[Ne��h��}*�*�����fA��;�N3H Iz~���#2"���vTCL�����ϱ�-��wR�<R�n� �:Jh��_Rt��EG��u �P�d�=��&��	0|�-�HꞖ �n�H-�N�B��O8��)�{��q�����-�9��O�=�Le�����^���_�=���34�������S���vInBe0D��G]ls���ӕ (���ݳ�ɸ��j�4����'�ZTӱ ;��'�f`�:�.����Θ8�gc�)��>(D���'ؐ�}�:{~$g��
�dIp��TH�� [�6�XY�]Ul\����QP��J��t�&<���?����T'q�MgT,e���{j  �����B������dL4܇��<���^�a��I�F�V0Z�Y���#�@�Y"��T�)a|��X����$��B|A�aV�=-���8��SH�m��h�zXȥD?����e�^���>m���u�*1��x���(��ᶯ�6 U���]Q��&"+c׻�Q�ُѷ��a��H��	"-4¼�J��o���`�jslbj��2>��/�I���Z�J���ĺ$�����%,D�"7������ɨ��xm��Ҳ�c���v�"�'�!Ȁ�uWLh�D���>�q�m�ĩ�E���m��{H����S�]�q�:ǼO`BgV����1s�~/*��c,�9'�r�y\Āv�B�/@�"�֚ �-�1��v7���K+�Р�9����,� a�R���1C���ttSfĦPde9�DT��� ��v׉�|�#���,�]Ld�j��뻒E�i�(J�N������7���I����o�F˜|��EYa�4m�1�����[������O��
�ɬD��n%]���S\awm�����kc ӫ��z�����"�19��\���xgD�������1�4f�?t)�~�&�v�o���Z�"c���~���;p�T���y0�^��p)��A?+}N�M$5��!�\��K@~��!������:�d�,�~�Zh�F��)
��,�DJ޸�����;����(�\����Y�A�[����3/�(���m��m���4�&&L����g�N~��{�P�TJ�l�,��2�_&^�V��>�-妮��ږyh3s_X����O�W�������c*P�l��\�jZ�k�Ȥ��Oqn��&�wSO�4���W��ٷ>VP���!�%�U?����9O����	��Pz��Ȑ���V���垼�TlJ���a���i�* �dD��\�'�(B��k����+(� �����'������[�Tj9��h?�X܍���V�q.d�㆓��ٸ��$a�Y���v��i�b����~z[4=^�b|DIӼ>ӱA��{^���[�^�����+g���:��c�n=���}���������c2����`�x�V�n�H�ZJk�Q���8�� �r�b���S��"�S|m�����J�Wۿu5;��LN�Y7uI�ǖI����n�SI��醙Q.D�}lj��ڄc���-����uAV�n�8�u�T�n��S�Բ���tw%L�{"�{����r���%k��.8o���PP���}�|��H����n��^Z0�� ���~��9�����<W�e�d#����d�S����ӎ�J�]ޖq%����ۻpd��l9A��u]����I�5'�$l)�/��;�5��3q+�-�}�P��eLև���ͳ�Q80"�GlD
�xn�WT���"���c��üs�t���w$�-e$��?͔K�#��_0T���<�倝0���Hʢ�l[��$��Nh5�3�Ѕ������Է[N��,j񊺩��e`�;�Or��B[��D/�E��_U�;�3�goj�ؑ[�及On�t~89��9�E���ÓD�3�|g�*.���bt�����ڠ(t�ҚjP3�Co�gS�0�R���J���cM����:�p@t�~����¿f����]n�W��!�F��O��L�9�)@������Z�;VĔ�ݴ�v�0�+���hVA8;��oQ��'�V�<��T���!�Y�q��i�ia�˱����V���Ɯz�68X6.�����p�8�	r����Mj'|�/^ӆ�oDԦ��:ϝP��b���V�1:+M�Q����"�|�ܞD>u�͉œAV�>jT(~����Y다��B�3T�R�D�����8h��bX����6���� á�E�SB�D�'�|o�Y�q����ݟ�G�w��!&��R-<>G������pE��D�BV�F�&��P�A�H�n�-�=��݂ �B}T{0��o���T��A�?gٝs�L뷗�{x]����S'P�F�f����,�~���� ii|���L�5O�Kb��������W|�o��������8�X]���|���g��{�[ ?6�����y��h^��>��.��H������Vj�|��-?���D#怨�g��4�N��?��j��l�)�[��F8�/���~�p�wD�@�H�%�K��	���uH>N���?�Q<~qi�����*M��t��ӊ�h�����DȀ{�#���%~�?@Q9�S8��Ϛ��p���{�x�ToO���9��O˅�a�9�l�47��� 6�R[����s��G�+r|G���2�[Zg^�X��ˋ�.&{϶!O���#:y�*�����������Id�Px��4��nU�����:t�w-��0Su�v� ��rЙ�T|F ��
���|22M��]��?����:$dv{o?����ONe��.�e�u�I�����u�$?G�4�,A������b�'�{v�8ݡ�rd��G9�M��ﱟ�ZOTn���9�����k�?�^e��g�éϪ��>G&A��(������z�aZ���V5�[/#�ˇ����P�����XFF��~p۠OGc	���+�p1�v[�D!��K��� ����� �)�Zvip����9zdC���~i�W+oݠ�o7a]j9�+t��%�I�l�K�_D��ǵ_z9�4�w��9�t���bVzs����U�s�y�X��E`��l�=vz�ޟ��p��[.#�[A/��7�e=�%��KO�����`�iY=�27���$<iw��35�0�����!����p�]��ŗ�&f�!4N=�h焸������EY��H����5֩:~��H*M(_�AӮ!���rp�o���F^M�̛9BA$��09�ܙB{�t=��D���S��NPP��<svn��6�аA㇍�Uȫ�х�*N��%TZ����������LT[89ao�5�o�#�zx"(~�?�O˴26�X�5l�B���+�8z�ڰTc'��yC{�d���ToXB�8#Nb�����T�it{x����~��v��La�b��-j}j�P����,�&��ީ�*o�>�3^}�=��;�lT�M��km��i�����
q��PM�ORۃ�ץ�lV@����U��n�%�2iC𷗛`�R�N�A�L�AbK�V�wz�uL��@�^d"E��C��'�(�[���W�H���	d�\鈴�1�o��{qk�2��ζ.Վɱנb���o��j��v�����6ɘ)�5����Z{c��e�Lg����[��Sf�n�x�]l�d}pLr���(��2My��X�&�v���Z�[�Xt,^��s��8N�ab8mP9�8���S�j�|��8��_̗ ����Y��X��������5
+.�� ��y��O�%5�ʜ鲑a��������-���pph�_(F��A�n��qW��i	J�d����(Q��iA)8ў7��9ɯ���AG��α���GV&f9��q���H�H�L�[xA�c����$7Y��7y/i��lC��C�?s����m��Fղ���L�_�c� ������ ļ��/��x��]�)X:�߁�E�q�&����.+����0;Sl��� �	͙�mv�ƋU@���f������Q��J�i��'���c��?��s�~z�ʚ! i���J�xY����7��|��A�"F9
�mq#9��@_�{�dYZJ�0�b��o5 g�>���}�Mؘg�i&�	O�����v��y�)��p�+?=��p��|�}*F��F��B����1ƛkh|�$��z&��W����%���X� t�(+��Á�~����/2�I�\D��[y�\C �u�	�]�2��^�
mݲ'J{`G|�6��ɳ�D���h%;q�Y��rVws3��%��������T��1O��Ր�Կ(��Hvi�A�C���%���5.ͬ���Kb��s��P>��Y̡��P9��O�;��j]��[�u�y_����{��aYF7�ήjh�����UKnȊI\��T���i�OM��*{*Y�k&���Pv]�&TD'mm��f�����j�(�D�}������Rn������U�u+�H(��g����F( {0�˲�Şzl������:E������Os��ܵ'�=����Fԯ��M䖿�5Y�/��q���#���'BtDT)�mH�U$�K��c+��%�Hi�;�h���P�>94�r��N��)O=�7ԁ_��ڦ:/�O�dFQVOn� #tU�\d0,|=�������87�Ʌ��@'�7b5�zR8�dg"Z�X�Yȫl޸����/�W��G����\�_DΦ.��Y�_�9�V���k��)]hl,4���͞��9P�'\���{�.9�����k< �R�ۓzC+A�^pO�r̐_��H�Z`��,�D���JW��Ƌ�A��s74��#`Y��dmţ��{c��#C�Q��#��5����ߝ��kއ_/���`�Bg�>_����J�21���i�&��H.����9��O��K�/��։ۑ2�А�� �'�j0ZnͲ'�nO�@�)�sN�	c�'�J�
�4��БR糸�AXʬ"��"`�T�����U<�]>a:V;���ܾ�`�S����+�'��C.���3��ָ���E�)�L�b�2��L'�LTO����C�6w��	�Pt"���I0>�	ێUp'�� �~�Q�u��s�F���&3ѥ��&�
%%�,uq d�;@�r�*i���%��%��wO��/Q��J�X�M�R�G��5�&�~F�ʦ�7�Lb*��7���l���dN�a����)ѿ�Zv��e �,}&����ts����Kpj4�cx�_և3�E⻴���f�P>n�W5&�%�AGڥ�:f⢲�I�������}�0�N
��y��q���p2�A�۹7q�N�}�Ĩuc���'!J�u��$������s������2�������6~��*8^�2�/t;.웺�!rh/�w��B���y�)�\��S�n�D\��%�D4�ß�j�]XYK�P`Im����G&�q\���v���$��� -@\N���x��E���/H�e���ʁcf�A�;�{�c\wH��)�̒�!Ёǒ�
�i�;���BQfN̅;7�͠��g)զK����>z;�<Y�Ǯ1i�[Y� �<�3b�\{MR�c�AVF��0h��Xqal"'�*`)%��R�`�(�j|[�����l�-��5�=X��
�N�&[ΐ����	?(����YQ�x
�1��w���1Clve�,���F�0���Jf�'s��8��F~�O	��,3IB� &qcf�uq�>
/l�`O�*4K�Ek%���Z�H,g^�PFi��s�ٗ���å�9�8�E��6S��;`����)d�;�z���>�@T�����@:Xma�u�Vv�<JN�f=�۱��2ܣI諡ɱ��','5v3hf�V�
� �x���(2��3A^�RGi�a������ze�`fDO��O탕�q�=�8S�򞒃'��/�UQgR���v��Cc��V��s�S�ް��1m��r�Z]\�;��k�������|ИTeN��w=Iwdlm��x��<�g���趱�ߒ���:��1W`����xUΤO3�{3'��A.�M���?�-ks�_`"�%�|��2�m�m��18�vK9���k
�Q����z�@f?�n�����D�� ����>q�u�� �� '�� �{aL#ڡg��Q�z0_B����V�..b�Ƿ�[�(m�r�$�tw'R�O��*��c����A�h����z��Ռ���^hLn�O�]��spuE6ѹ��e���8��-�Y��?U��`X܋�nN��u� N19�c'��������+��,C\��2R�]q���ďo����ꆪtJJr��yn�x���w݄�jY�RH��aK���Z �2���Z�	�Z��@� 吶���K��J��*���D�,d6ڊ��Jĕ}��A=:�T� ��w�nONZ�����K��𬒽�2�&Y��lY۔��a.B�mz���j�6;�R������qw�'@�Xߕ���CQ OMT:M�S���Ʉ���Hl���׌ʕ�JX��)q�	�w��=OeE�<Y�*�G���(o��Ts�Q<��^Z�1�������0#�:���E�q��F�
*}ŷ��?�g���30�W��Ą̏�<.Sád�H϶\��n�s���x�"v��F��j��K$�1Z�a�Z�}��'��&��L�vCȥ\ �wGĻ�+So��.��l�6a�
�U�����MK��%"��V�	���7�N�V3x�gÍ�b\���?=M��7��)�c��6q$�LU�Ov���{���#�|�v��+�&k ���VV/�(�\[�[�<��p���J8�!J��~���5��GS8��*��ER�0	���;���\��N>�h"Ay6᧹.ɋ ' `L���B�f�2J;A�|q��:#��GˤGL{4�U�A��d��T�W�xʶ�4K}+z_ޑ�ɍ��Q�B��e@C����H�L�ع���?I�7�NNB���?fd�2�cGa�K�R�7j[���[Q��)VX��Լ�ȉ�r�0�
��� 1�c�=�D�[�GV؂����T���x�	�|]�!�Μͽ�ގ��7� ��k�(n�'�����X6B�1�"�tH�5T�����a�X�3ڧ�k�a
+T1��\kam2�oQs�H�C��@��"} +�b�\�@�l'�[�7%�!Q�ܷ��$\�')%T݉j�<�`*Lh���ç?Ee�N��ӤNjM���ضevO�R�6�V�S��j���Ek��\馰�4��D%W5��vby��\�1�����f�Ȱ �x�K�х`g4�cP��ǳ_�5�0˄{�UAB��g����r��P�v&ܠX��!V	����k�n����S��F9�@���R�ykp�>[�oDq2+�D��E;�B��0�K���JV�Sl��t.�ok�ȶ5�UA�0������c�����&�V���f�b�wRѽ�B�nu���xp�����@�X�@H�~��1�7G	<��j \��]���1�m_�/�8��֖Ar���C���G��m�Cr�D2�ZZ�������cX��4(�!�SK���x����}+��I�s̄��P��v��[��}ڻ�v�Gʴ�ߢ���;~Fm%k��'h�Eo�7F�d�3��d�#&��Y]���5�(ߥ8�뺀��|�����Gp���+����N��%6�I�U�r��%hk*n����}p���R�<��!��t�z�U�S]�K�6�*�&�W�$��j�h�MG�m���&*���]Bw����.9dŕ�G�\;���J��b�}W.��}+0X�r���I��<)W:�#N����pT�j���� �F*dܦ��ޢ�k�q�`bvʿ��*pt��=����8I�E���g��ǻڦH'�,Z�bb���=F��l��zp�LB1��}�=�l�7'#Wx�f���C�F{��o��Oe��"�U7���-V�����x2��=���i(�4+@�����P���aa�H�h�{c�E4���!��?Bm[�6�A�N��ߤ�m-�\$Q�����������f�Ļ�	�Yنu�O�U�|�e�.�@L!d*��(�j����tS�MT
6Uq��,V��'��ړ֤�X�_<B����PH����s�p{�z�P֡K������0�G� ��i�R:֦|{˪<�1cjʵ��J��t~����NL8VR��!>YyՓ5���6j��2�D�vl`a6���,*��z-$�kSF0ޜ���H٦���kGO,� �@i���P��=��g�8J�@�NX�[Ɋ�zir8�y��5�I,�����=��K�C�
�+}޹jQ�v�8|�������H4L�[K���m'����"5��C�R--�IO�R�vZ=BxÕ�r�jK��=��>������?��b�@\RsF��E�5���b7?����M#
v}�,��4J�$V��\9Lڛ\znq��?���寲K�S� 3K�6����s�w,�1 ����h�)H�c��d��3���Yהh(ZGADDN�S�h6\zt��B���2��E77K�q����w�4XZ���oǫ�=��A,�8�·�c�S1�p�JW����E�/s�J�sSkf#����ߕ;���b�Z]P�����a����UL�{�;���� ��0*���֨�5弳~�)b�n����{(�MP`6�KtXWM�E|ן��LBpD�Zqxj������ˍ������~N���7����^d�B�]�1�<��ٰ~&��g��$��c������{`x\g����i06�4�_IQm�V��B�J����H.��wU����M'uVPd�вz�l?������/-Z�}�*���x���Q<N60|�7�e�L1ی�m�d�j�"�{d��A��*�����͜@�=�ݣ4�ft�5B5B<��dͩ����u�r�d���2�R���wئ?�S�/�-���$"�b �������Nq�#�q��:�-�H�ѥ�{�m�K׀��:% �p�C<��Y��M�V0��I�3�9���br�S�w�e)C�9�
<�3�zq�nï�A�2�t��L�/ـ�Ջk�v�v�³Ⱦ��I*2���@������Jެp�e�6��ܡQ�"�Kz��)C�-�d�W+�D�Ң�y|.Ov2��x�J�J�w�u[��s���ĨwX�8e"�8�3v<�J\�y��\�R1���g�����sEf�nò�\-�/��]e�`��.���+VY�-,�?X��<��_X� ����L���Z��(�r&��,Vr�0Ew:�)H�\N�׏�~L3�o�9OBԈ��fn� ����&��¡*�d%���"袬������#�qw���K�������Gt:t�O��mR��zX���V�}H4�n��.	�.~��X�w۩K
%�\���t�a�̢i�a����.���k1R�n��P���+Z�_1���c��!-�(�_,��_A���@��l�F���th!�;�U�z^c0`�F�1AI��d^I+ƽg�q�#v���U���ȇ����C#�幽bl���p�♀G6��;�k��*�X~_u�g�.�zO2�����cn���D4��!�����DB���Й��1,�7PiB�!U�R�ښ]��C���f���3�,R�jxA&�G
1��S��Bz:n���<̖;��x*hό�%ë�[�-���x�5uh�L%.dp�پ.'5xI5��0T-%�g�������)�Id �uGf��D9ȝ�����z��uy�#g3�wD1�0��ԧ��m%��3k�X�D�6y�f��N,�\��wM���2�.ԁ�	.(�;��[�]Z�~��x��-t�F1�3S�}k�ҧ�A(cr�t�"ƭ����N�[�8�kܴ��h�#V�'_�l���v5����S�AY)f�$���U�-�e
J�E�=��6$��ت�U����(*
�V��U���.�G(���n�#۸5��vj���hlk��I-��4���"��@��E�ˀ����8�=6>Y���%�y2��gq��{�?j�>��ѡ�e N�j�=�р� �M��x�QX�-�~���q{�>�`�T~u��f>�!*��~O�р�s���>�u�MK0c�t8.}	���g�V��u���,����<��-�"b?�	�d�[�E�
�s�[��:�j�g�W�� ��|ů@fI���� p�vSR�,��s�,O�U`��-�󌛐�}���p[���4S����CJ�祂�t����	�XmsV!�tb�]�CL����<��)���Gu[�G5Wr��̲>��މ��G�l��*�8 =합�ej�?�*������yؐ�9����E��O��G�Js��oɨ:��@���tһ����T�C���0t��GR؊<t�̓�|Z(t?�7f>��e���_6��u!�l��z8'[�'!ci����F�g���\�B��?�i&[��0w�r3����\ޯ�&�)�iBpy>�!x:"Uj�&�ط����=�͍�в�K����J��,T��憫�f�-��M�RݤkA}����Ge*���ffX%�8Z�C�G6�.� M�����@�E=�-�Z��f�d��|���՗^{�1�� �6�[~�R�v���ޝ�Ҿ��F�v��J 8�����d��M]T^�ۘF�G;��b�t��ں�.�R��F�!`Nj��7q�J}=*���9�	͢P�+�v�����X�t�Q���*n�����=�~����U�՚vj����}��t�n�ު�
�5F�����.@�����ƭm���C����r%�MR0�0�*.pJ�!d�O�L����C��3l�cc|��n�I����\)W�\}H�	�k�}V�?�!ʓj�R�n"]4�#� ���Z6�x��r������I�o�n�LJw�NW���Z-�s�'?YBa�.����<E$��Y��M����DfL:���:bq;�#e��Í�C�G��xc��1���f>�Jߓ;�W�M�~�ء� 7���}�^�ظ�5���&�q�1��ul�Hi�(���EGC���KaMOJ�L���.h�	E˪��H
ī�a�E�3�6	���.�0 �79У"���6�(1h^0 M�N93�Q��6�t{/(V^����%���G����麢�i�5Ӈ+�t�(��� i�K22^�;[��}�B�8'�Q�=�5�K�1�JH�X�)o�"Hџ-zK<�g��V������ l�MD)w���t6�{D�H����7����=�~^(�`�<��<��8B��K�3K���D�tN���y����%�0dt&�u��d��l����+ͯ�԰@��Y�6�}"���,fv���J�����[X,�s}č�x��*����n��#�Ժ�e}p?����sZ�-/5E��b��jD�d7H���$;h�@�^@��#�����fy�哶d�pf�����V�X�t���Fa�H�����ryx�I�gm%�	O�%䔱;�l&j�Mq~=�W>�x"X��`f8�+����.nNTmP��.l�3��N��zZ��bޜ�v��.u��\<�� ��I��?oN'����
[1\\��?�R,ɸ-��b���JC0��U^���S�|��a�]g�ip�<�gs�e}���[9#j2�Ӳ�X}%��~�%�����6�J�-7�_��2�͉�X�
��톩G
hVq����xD�jx<.V1>̉�`���k�S�p��!���Iň�(���x�"g\��T�6>��)��Ťr�����h	�p�)����x���[�w��7��&���5yV�e��/$볇��N��ї�<O��^�����]!w��!Hҏ��:w?����$��%be0�.?�.`n����8��o%Ǒ���N���Si�E]�����e���?t������tZ�m��z����'�ሎ�I�3�deS� �a\��Ҥ���g�q��q} sC�� rW�x�*/��~p�x��X�j�9_UWh��ؓz�U\Q��Ѫ�sF8��YJ�(����f�������*�X�%%����e�6.{�)��Qt�sh�l�X�V��V����s�����4�u���;@0YOb��W��fkQa��� {\^�'SN�}EĎ�k�_�A��z�������"Ļ��3�_ b)���]滅��fE��r��gx��S�%��0��':*�+,ڳa�5��#Y�jRIn3N; ����	kSA8�|n�D&7yIr\zT߹0�6��gF|�U��9�ܢw��~1G�^��5�J.U��b�r�W��#TRNQ�'��W����`�����I8 3 ����GhR�x�ak]���Ƶز��I����$4\{�J�䘕ۢ�|e��R i5ϳ$ҟ��4��q�5V*����/�u����`�@DN�U�&�c�p���q�(�3���#x�ˡ=�}��u�`4�Cf�"�6��k��p.�9���m�x����Ӻi�G
8��K`;���ghUI��T{$2�.�u9k�m�e����+`5D��l%�N����2I�tO���xG�~,ͤh�5�U���6���O��fcsFy"@��������|yw,���~�R���-4Rh�gUp!�V��W���zƈ3�M��Z;�Z<�_���凙�)�X�w�9�� ������[1�����c'Pc~PY:�C�I�
/�D��h�-���~Kl9o<5�+41�R���fƔ�x�n�n��2e�S���˩pʳ��3�+��Y bn@4|m{�����㲾Fo�5�'7��e�/"^���t)�EW�-]�g+�{�*���W��F��㡪T6���G�sqe׿:�?RY#{9yR7��f�*��q9*��.�fe =��E�H�q���Y�Q�ż�Ř,�{�lÆN�>Jz4-��)u%���P+�E�)
Fb�˙Kf�s�4�I���듂i�*�3�!yc=ž%0�����؇�4���z���n��TF�1|�sX�������Z;�$�˘�����~I�%��WC��`���\O���.��=#t���-̑x��}���ӫ@�����t�v6%L/VT���ίƂa�?���wYEM[d8�W%琕B�P����vTA>[J�$m�k�� ��f$Tt &�J����=y���>�����!*��	����P`f�)鰛.�F��N�[KRE1�R�L�f���~�_2q��;Z<^�3/nz��Tcͩ�b��l
��5�iW�q"zh�q�d͝�޸�p��ԏX�W�p�i?-�7Em,Q'AT�~�Z5;� ��f�6��:�bcn4TqL�3<�ai��ƅk;��ߎ�����".�1���ϡ���:�)���Ƽ���g��/�qX�zg���X��������Ħ�� 2�s^��)6�U:���������FDڪ�iq8�l��=r�c3J%a������i�l�n0�!��_���t]m�GIg�
!�C�צ��sҌpEE���R�]a�t�����]���uC'�"���)�2�������`�\�-`��m�ϰA���c��7$��� /���`fR-ԉښ�B�w����K/��qK��a:

)���w['զ6b�B�B<�M������"���<Gj	P5,)Ru/��4}a�	��˸B�cŦ3��tV��%��f�I���)#k�=��yP]K�l����s1�P�Yઉ0�`��J-;!tPhJ˵��O��2%�7�T�����+�
���2�:|~���&�<��C�7�_��ŐG�Mq�r���4��m�F��@�������y�
���)��Tu��u�Q-�0!�;�ħ�J0I��+�s�J�c=<�	�Gx�:m#�\���;%Q�U/�������EL1=�:�^>��,M�tFC�F��Q�/SɌݻ��8�	V��څ��.����-�m�`��E����S�d/_lv��K���_V֢)�6��b�w�<6�iJ-��Jpv�_�i��l2%13]��W�N�q�ʇ��͕�J���|mH}�qJ��J���5����?�y����� �D�9���Dn>�c�pa�wS13�l�4�CD�����3��v�:���@��C����nC�����%���Z����\�<n�����O�'|�SE���6��"���M�ǩ�pj�������
�I�)�#�a
�q	��11�m �o��h���j���L:�H̢�U��FT%�J�����!��2O��	��V�Յ��Hگ$\�C���!5����~��|>-ZZ��$��HB+I�������,��z?���r��9(E��7���4����=���S˥h�6/��Z�Q��'�ʅ�O�!f� ou��#>�5ٟ�e�By����C�N9� �CrD|b�	�хJj۟oB�_3�˴�58wL�Sn5�յ��[���B���+�/PfGHƯ����zn/.ue$��/�9yq��XηJ���X��A�iN�Z������)������?�C�5*���>e��Hz�|d �kC�}!V2Oj���V?�7{
lG�Qf��b2�5v�v��P��r<��������j�0�36G^�q�>��y&�g6|��)oesBŏD^� �e�nMrHf���H�6�%;\����W��qWِ�� �U�p�D���T̗P�o$�Fxz�������`��kf�"r{�&$�- �Gz����;�GIGJ�8�C�aD;4ܙ��F�CiW�q���H�9�D/�g6�Ĺ�~�z���q+$� i��h��2��J�O����Ǒ�On��,�blD��;1���qk%���BQ�&�.������E�y�s�1�1L��c Qb�=B+P�
dK#�$M�j�Z������~e�*�cBh���XU�I>6:rO�:¢Ow��F���E5�_��I�㆓.+���o�vl<�p�A�a��sp���(�!��r=�*iv��cڬ�W?��5HdӮ�"���Cv����5:�ʶ�97i�.�j����_��z�Pܧ�|{54\0|z�٧�p�j�R��#/��X3r&`rv��R���'m1��[�W�=���Q+���>��Buq"w��kj��b����y��1���qØ�>��̾��J��Q�N��=����g2i[�=7�2W�a�9�^�F~DV�|C=������T��\z��i����h�:55�S+���.�q����ܑ3�8n0^�׮GC�;c��u�q�Ԫ*#N>V�s�3G��7)Z�(���wIK9'l;��br2��/Ȳ���K�FÏ�˻w����<LsM��wEI�;M�9��ё��X�@0��ӭ���jT����1A����b���Z����R*�ȝ�w������Q��j��*�o��']R�qw�j��F����`͸42($��O���4�Q+�׸H|����p�'6���� ^�z��@gd��H��b.��}D�i=�^���;�س<n�*�e�yƲ��=t�G~_HfB�O�3l�����U�?�h�`` ��^�rT:�0�t�'���Ō���wW<{�b7~m��P�&ư�g��G5�f�/�2���U�F�ì�ԕ`h�>@P�y�r���:1�S6v9h�1Znɣ�J,�?`v��|�b�}�Nөdkx!�Y�f�:��_|��J�GmUo�;��`*�Ĭ N>g�sJ�w�`:��%K�l��ȩ	Zab�Dhْ2�HJ����Ҩ[���]B=�Vl.�O�N(
�����&�n�ޚ��Q+��8XV��$��A��mE�Z���3]�ƴ�n�T�y$6
W�&�c�[�H�?롘@a�����`�H�ߤʓ�,?"�)}��}?E�F{�o�E�g`[6��Pq�Z+�#�RN��8,��hΒI�P�?���I�>wB�ר�)���U��X��@���K	#=����Ek?lm�Fq��m4����% K�|�2�����P�s�b���ru�� S��X���h�s�g��*������D<���e�Vz�ي�:U7�*{K���po�-',+R�����7���ta�|g�t��!���W����`z��(]v �
��w��U|�'SL�o`c;&\��j.���ߝ���;ikƮ}4K�u#���sZcٶ/7о�%��d~��$i4(j�6��D���|@�'j+��#��5�wHN�L�H��8�/,���!�r�!p: ��o��<7�/fQ_�O	�vK��s���Q�}�>��U���������0{��<����pS��㞬�b	�M^T�{��ak�*�P o��j����%�g+=���^�`5q��y�Ea�!���جƬ�� �^Z�0�C�����N��q),�h\��	�#���n7��l97\���B$�7 샨�t��]��K[����W�gbL-���3��K��l4+�gk�e��Ce�da�~�n�&1��_c}z5�.7���$Ѩ���Q��_1���J=pju���g�w�`-b�ϼ¬[)�ZA�k��Ⲭ��=�ɘ['$W���Ι<4ksE�>�����+�5&�1�ݨ9�F�.���l�)�M�J��NB_�)������:����!8��*f�5*CP���lσ�+��QM�l�NF�L^N
��&
��7͉Iio�,�I��c�5z9X�Kl!�����8����T�Y۪��"5����,��0��r��	˩�����ݒ�h�ta�����o�ޱ*��.T��)u6���|�Ҟf/�P����,	�f�Տ�(z��N�qѡ��¦�R�г���n�qY4^���4���-�s>�� IT^��j�d�3�煩O��+�o�?,W�P��|�g�p�T���U�ʇb���v��>et�"N$H[�;�5��gCXUu���f�٢��ۋ.0��rCg�Pxd)�q�p�w<��ǒ�~LhC�:�U���P���Z¯����W�xoP�0�$mZU{�^��d˰��3���h�s	b4u��$i�a�}Cq�Fkߢ��{`��������?<w�9~���dX�%ý-���>�N�7�0f�O�?�X�W��9��dP�cuה�sJ�76雍@��]x[_�FWk���f\��[u�*���H�O9Z��� �t��Wǹ鈁t�[�$�}�������j���N�)�k���ab�,B�$���
W��CEu1��`E�+2zql���[/;KÐ��;d�IP��ݐN$�Q��H|��4DC�1~ϸ�	>�T0 �Ӥ��p��#��܈����+m1-BY�l��ӮiD��ɓ�0�p�xX��3ӷC>��]����c�:6�"5Դ��[ �RG0`�5m:�e�!����M��1�0	E������Ϣ�2����'8�"��M�%���|��e*ֵ��O�&���<p(�Yi~'Qy4r�� ��-�[�(���B8� ��\=�o�j�AP�$P��u�]���mn%�����|��R>"��} ��!R�c9���󔗧�l�LdqZ�8��=&8�;�L��6��?�u�zuK���X�$�}蟷BO�e����E���y��q�2��QD3	-svQԻ��p�Fy��s�MH�Il�?���ee������N���;q�L�q�{q��u����I�f5|#i_��ͩ)����� AI%a�I`��H� ��諿�.	K�'�>��<��;v5��
Z�f���#�����nR��{ާ��ql%5J�%� ����?zUC���{-���m��kQK��Nz(�U�I�	!�`��F��FP�&CC[U:.W��f%.ȴ
�M3�J��������d��0��˒,�+}��c�?�9�Q������K�ۙ��?�e�<�Ԏេ�_E�KXk�|Sob���^$��T*{Nn/����:�'e��z`r3Dz7P��!�=��9���Bz��EwT�\�Y�Q�X.|�$o�
Rx�
�1�ђ�"���0uT�Q�K�έ`��6�*��'\8���� CQN��dZ)Q�<H���d��,�dH�;:�͙�_9;�^�@�u�'�~jh$D��󎔺g5$�Wx'���	^�'i��)�('eҽ.s�3�[A�I����n�@��CP���g��n���$����m�mU��W㔾9P�[eHR�'��@3!�?h�\v�ڢ߶gv���ҿ��i��g(��k2�����7����D�y���\r[N�֊��@�:��]���X
�Q�tR�L� �WW�>� �Ѧ��}���S,��9�*�:�$�;w�����g5��Y yv.�E���	��R�S9ڂOQ��O<M�������{�����"�~)�b��˵<#��xhij!o��G�,f4=Pݲ��#����Esi̾��(^0�#��x�$�]W���Ln=�*}���FOH3E��X�-�>wy,�6���5/���@����R-���#W�{��K��}8W��a��\(<�����V�_�W2{pp���\	�T�ry�R%V��w��xH�#�8�b�y�0��؀�=���
0:�D���}�=(j���[*�C�'�d���&�:��aZ�=�?XQ;�\�?��&�-���:�����
�,���9��2З+�\.�G�==�����T�j,y\:��+��􎋷�� ܍m�K�'�@"��Rͪ;ը��X�A����޵�!]�IKQ�]Fރ�
�_��t� ���4I�Q��E�ghDr�̏u-b��,���;����"��Cʼ+�˫NU溃��+}�K�eo�ȍ���r�&a����+(�_�kL+�ʕO:�W�H۸�>݂�L}^�p�����@�?B��9��"p#j�'x�^�4�"�昩�5�#�<����-]6?��Ё�2mإc�q ��D�ކ�g�xڥF�?����K�8���� �2�*FM�]���'s�m���+��kz`��3��!/W��z��;%�:�8�Y�#ݯ~1UO��5T�~d :Q�A�R��z�S�d$㴁.k�y�.����,�̗��o��%.��5V���U�	�KNv_���{0�.������!
g��Q���g�2/�Ɖ��Al���C��6֩*��+���B��ԇ���l��S<+�e��D�MC�P�b�[{�Y������Y إ�
�F\t��S��y��kU�c�1�YI�v�X��G�?|n��.K#PZ9g&�;a;Z�T���9s�Z s�8J�X c(4U\�����s���K_;>}�l������-��놴�A;�%����۪�D��z�w�I��Y�Z�F��;"��>kn'��e&l.0�\>�"H�c���/Ef>df&)3޼	/ݞ��=@� o��<@q"�]��H��7Q( ���?VnI��uĜ6?
L�M9�#Ǚ$��c^�C�7g�!`dV��n�]F��|AL�DQ�Ѥ�:B�4@�Q����pBeW� ���A�n��_�*@GΤH�����v��f�#>Ӏ��Ҽ��,N!�~xs�B§s�eb�ۨ#���118�4��Z���)a�!O|�N��u�@P���K�^-h�y����ʓ�Mz��9o���Z}�T��^��=�QSk_�sl����8)�>\�FT�h� �eSO���Ug���X�x'M{��f��e
��b����m$�X��sKG�aMU��Ӑ	]���g�� )�-���*��[�_(C�S#�q�	�S$��Y7��E� i��lDmH��"��#LɘK�S��o�W���] ,����N��[W-<����jxu�s����+\�n��N/�ޥa�	�h U���)�����J@~txu��_7�����'��JlQzd��(�h�2Q�Z>���(	RJ��ۢ���8���4��$�GY-+�8HB�g�p2qq���;���]��\�AG�1�S�˃����j�S�{i�r�]>~�9�+$ʾ5�v���Q�,J��g< �Ӫ_?J�c�ɬ�W�+��/���O�U��VH��3�mxv_D(}�LC�Gp���K�nK8c5{�Jq�1t=ѧAՎ����b/��+$�������L���s��ⱼ���Hеv�@��[�vpz�;�U"']�w�æ~�/��E[�},	�6��< M��0��ī5��K))���(\r�k��,8�O�-�Zl9��Q�ˢ�m\���H�� d�H��|B ���eh����F������A�@�����FN� ���z�j�������a�A�u"�AT�/�i�����.�~�stm<�~X3K� Ĉ�UXb���pZ5��=�ۘ���������*���E=W=��/���%~���W��?hf{�x��d�M���E���m��F����4y*��� v҅9ğ�1W�X���8�3�ޫ0��y�1�; 6̂���Z5��{��H�K���`gPi�������&a��L"��^�펴I��jnҀ�?S_�1�y̲�z�N���U���+� ���j��8ڋ�?w�o��+m�L�X�"���=T�`^;��?(�n=�4Xນ�cg�&���ɓY����DEs3`Zɳ1�/�>���y������n�s&˞��a'V%˒�-{�A"f���<G��[Iy��(�l���3Y�� @��R}r�=D�*?[��;������G�7������c�.^3��>el�?��w�]\<HX��z�����T}�c_��3���!�r�S,R�Ð_?������P��Cg�)l37���}-RO�9�~<�5���
(��,C����@��r��6�˖�p2w��Pi&��ܨ��G�1�$�>|H��o�F u�k�o���	I��o�,�I��'�\?��0J2�M�a�_�����w�p'�Uמ޷������ǭ9��{�mJ!�qa��Lyo��9�i�?1l�ݤ�;sN���=����%'�ma0v�Md���M=	�W �q�(j��ֿRٚ?��̻��9D&O�'B�x+�3��1S����Ș�������󺄶�:�����O�����܅�]|�����OM)�xd�"���xP���9�����} �^��H�,'��t�����\��q�!�|u��Mr��'���Y�]@�s�"L$ǉ��#�:�s�x�iI6��Y[�)��\d�Y*����Y��c��`&H6��4#��j��<:u9��e���J��y#8�)�R�P��&m�o�)|Z��#H}�`:�,�{���Ϣ��Ѡ�d�`��ξ�|����܂��[q^��Q9�5l�4���Jl��PX�3�nM��������Q��jWUhKw���R�G�h�	!P�k��4�W_`�Y.��Ѐ�{()��]���u�F�D�c���TU����@r9�fTS���V�]|kV)��/��X�I���p��~-5v���L)�b�׋ ���5�8X6pl��
#\O:kM���1H�l��BD�Бp�>*K��G;�bqm�'Y�`_����r��A���[�XY�� �(�^������1~"qp�W�H.�|Ѹ���}�N�$.�>ů�]��Yٶ�$�yv���R8}یm`$z��B ����<A��=�F�=��VN�vU�3�U�
��_�������kϣ���j�m�����ov���`�<r��;�4��/��t��8]>�HCʸ=��	U�\�$�n�G�k��L�����R�B�
E��Y����\��}�E�1���?����6b5t*����P���1��ɾ�le|�g�����O�C��/��T���&[��5�U-��*�U�I3(G��SA���^ro�GC�����G��(�o�2W.n��5����)�ă��PQ�LN7x�x��L6w�m�ɻ �ݦ�`�x��`� �����i�n�C2� �1v$Μ�X�h�5F�%m�ujN�+���;��<j�D�&��`Ql��Z	5 ��}T�� �`��%�ވ�9�|
	T�a@�{O�z��R�! �Z#����� ���f��+��Ұ�M�(�Α8{��DNb]zu�Q�-�4����[��S	��"M0�A����;H�g{��!���M��@
xi�hH�/�x@
��
���qȇ�~q�h�Xb���5�wi��,Nf��,O#6X|���2��rI��,��~�BP)+�o1�H��(1\ ��������bڵ�?�]r��0lx�WiTS}S�\�7�Fǐ"��=����4�͍UT�4WG,�(�7�����CvN���`�8V���Ǖ��#����ا"v����%L:�u�R ���ee�a;�·�L	�6ߝM��}(����+���l�}ɻ���wNG=qSy������MYA���ʑ�U��/�ݚ��Իߊ=d��[|8�T£�$>��zpD������t�*���8���0^�.��hD(m3�uL�+���@U�L2�uzo;m����V�K-�ᕡ��OX�$�fz���2��%�2��֋22R���r�?���~_�C�~�bKA(��^B�z��;ۯPA�\�4�H6��N��tq�nt�=ˑ�2�Z2U�����N6��<6"��g��j�o�5ʵ����7O���fB9�j�u(���wo�/��ш~�oL&0!RQ1&f}��v��'WI��+^5���3���}���)�.e��#Y!���p ?!K�FuW��$��
	T��R��E�s�B:=�u���r,��>�;��}����W!�2@ύ�@��-z�;V網`�)�� ����=�B<��{��:��W����c���$u��j�H��_�6�B �E�L����wu���E�&�jIί�":I����r����^�,��w7�:,ѻ m9�e�DZ�I?0+]$�=��u� �
;�+����3��=x�Ռ�D>��I����ls5��tRQ#5SW"{�F��r���,.Dw���+�Q��>����dC�������Q��C�֕���n;lO���z� �YY������c\�&('���!��.pA��{��x{3i&q?��o�L�p�6�ڋ��#��M�����F\���w'��5���]I�y����Jt5�)�����a��,]6��Ϸ��E�\d�k��dt�S������jG*3e-�{�떲@��E>,I$P��"��n�/B#4]�&a _�*��z{/�l���b�!)��u�mƞ�H�	�M�?��[$�^��"|j��6�����O"��.Ӄ_��a�±l���Vnԟ�/Q�\6̈́�4Ɩ���f����.	��b �!����{?���9�)8��|�p6�
�KC��2 +GVħ�L~�3g��]�2_��vM�v�h!�V)#O���/�������1�����ׅ�=��jm����lGŐb#�b�	��Pt|�,��ˎ`>O�q��'�X?���o�J#�-�+��W��2�r��?���ς���"�'�P�
-��S�͜ԢԻ>J��A�Q�>J��"�4j�/v�|�8�����P�!�s �_�8uSB��E
��L�&��oi��<]���� �/���1y�N��6/@���}�Hu��9�204?�b(�����YX�#����cu���t��f�GZ $�Z�vi�#+�`���� .����͉솺�ة��:��~��yc����Om[�nrH8�![;���GM��Jg�Lфii�?�d[��&*H��|�a���=M����
|Br�;�(���(k�����<������Pc�%h�>���8<"�5�J{"9��5.$��Fvp���V�Y,7"�oX0zIvo	:�1S]v��C|(5��C����M9�	ak�����/�1W� H������;q�
�/\�}s�ciJ��T�yi���NL�D�@�͊��Kw���@���[��7F��k�CS��Z��<��v��.BY�bKn6�	j��Ճc�2���rz�n-f�KɁ�^�1�<�x`��h�u��ZW��xk�͂V�XY�ⴖY�t��̛M���C�8�8Ӻ`+�\��a�����e%�����}�[�JuS�G#g+ε1ԌeK�N{!Ҋe0��R����&�,A���~H;�����4�"�T+{9�|�aPУ*ĺ�����t�טVs0�df�U[����n��r��R�2j��O(�6X?h,k�&���'A�*��P�l�^'S�`�������is7�z%��oqNG(��B��������7x�5q�Eo��T��x�X�j�"^�zr��Rrl�{�5͒����Px�(������um)b�Jóo����L��/e�b�5(-�G���h��B֒�����W�w�ܳ+��� �x��ħ�V�_:�����+t�ɧ���
3���[�#��^+H�;����@��mݹ��;����enZ���@�'I��E�R������H.���-=B�vuIn��˽g�vJy�a�!���׸C�O�4����(�d4�]��P�#1�_$��զ& !�x��a�<r���ƽ�t�4y���QU�nh���Dn >�s�t�j9��r9}�'�L�e��i��0�=�y�P�zhmE��B�V�a�L�W��qL���g�8��$VI�/-���:�o��ƣ�7~�3�����.�	��85G�ߨ�޶�a�vw�]�Ԣ���{����#p��g�S���q��4V�w�AX��P��k��c�\0��y�/�{&%ϓ��2q<T��8GT�b�>�u-a�$.�q�?Ë
�Q<V.RR��̩��`oz�xB�J{�SD��6����fU��F!�u4������˰��)�X�Xs�	3���%y�k�eނ�m�q������Տ���*�~�Z�;��o�`��/�}��%5�	�`�8�yl�!�g�;[���{K�W`�$H���'&�ӉvZ���.���J3��<�
��x���� t��2|�j�R���ătJ/���vT/"��>4hWA�jJ�rd'x���A	� �J8��f.�n�&�ejBKl5�V�,��u��v��BT���n����1a�����-�����g��,
Q�����m:�Y	�)s�����7R�����xU�N"C��&�#y;݃l���v~��Y ���|a>�z�E?�h��E�F[��u/hN�k��q{^���?�83a�E�W�i�����`��M��1�O'F.=�{2��{�����U�װ��,<�����^�u/���@
�|D#UhA�����h@[�s�J���kwf$������:E%����Oc�0}�^{4H��|i�q:'�3@�*�|F
�zk�u�ui��
�2�ả���k_���4��F��)_;6�j�3����2���}k�K3���eV/��H-l��>A���_5#��0�Z�k�D���]C�P)֘'�>�*>>�,VH�	#���h�֋J?��J}݂U��e���3�T����F7� "}�"�����g�q�LG�-����f��jK�5�z�J��9H)��Ӂ�>Rs��y�(}�Q��&q�kv��.�)�~3��A�;EN^���0�l���j����m)�����d��JJq}��=Εz��gvny��)��j�f\�`�L��2X�a(�DP�����L�_�Yc�ى�w�V�8�Q8������Z��{�R�p�f׈�������E	V5A�eQi���,�vK�<�DY��� ��3.3��L�)H����K�h�E�b��?Eb:���oz �YAȌ��U���𶖵�qV�A����wy��6�S�����1���A��w��с��*�<OF;p.h�Ҫ�Ԉ9��Q^~�!}R�f��Ue>����.o�15�=�37Z�ǻ�S����T(w���~l�� ���$�l��6E۠��z�Cҝ�8��X&���W*��Q��H��؍m��w��t���4p��<�1�ڻ�	�إOcR��P#N	hs�N�|.���� �`(
��F�:��>#=��E���-tJn������kPV̝0Km�,�&���؇�}<��,O C��,9�_6���D������W��BO%G&@��o h�p3�6u�k�q8��[.>�0#ۦ��BV��f��4݄����^x��Ru���:Ǣ&����n�7��ߠ�~Ȑ�<�qLRV��q�;�:t�d�y+���Z��P�c�?ܪ�����v��-%��Ш��P���h�,��sX01LЌ��}����4���J�1���70 0��2�Y�}��ۀ�:���{ěm�?�z��ר�(�,�h����4ؚA�'����ML�V�5Fo~Lq�E"#L=t�\��\����
%EK�/ٚ88P6���ڌ��+w��Ǹ%�^���d���������&����� J�:=� ҅ �����T�^�"EJ��V�PM��Q�f6�u�,�b6����.N�	��_c����k��T*8[$�Vҭ��ʩ�l����	�H tA���wR��7cי5˫��#�6�/�������p�S7���=�~�f�<gL�Sl@��(�/�[X�,�k�.�Cz��psYuq�?�$����'�4=�)	��Z�J�$T����ˑ��&�-�J�o��sJ�hZ��^*�yhա�F�Ӥ�p� �k�@7w�x�$r��v'�;��D��$-d�J]>ZԼQ��=�W��h3g��Y%j�0�aٻ�R���Dq�J�5]`�b=4UW�bv��^ء[z�ᗙ���1")�]- J�|?�7��$����WQ��ib��j}	U�����&U�=�W6d��su̟	z�Ba���fgI&z�Tniس��=e�nU���8�ݿ��-y��'�@��ݩE�7�x
6��>�PQ�z �����6��S�B��/����E��뾢|í������G�톢)�D���N�A���̞�TX��c����(ш��1&��B�ӂԹ�؀��_;��2	�-@��-f5�4��tjD�򛒀C��+��c�Ϳ½ c+�3
������9k�٨�1є��e��/�t�U�l�'4C��1�^ƥ��OpۧGYk($��H��97��[�{8���-��6�cה�pI���y{�G���-�;Q��}+j�}w�j��&��P�
&��Ãi��F��g���T��aw�$�w�QL9�s�;���%]_���������)D �]�|g܌v�t���$�wX�V�l,�����+j�L
�}��(���]�>��c#��$@�"����c�Ǔ�y�*N\4Xu��xA��SP��6y��*�T�!.n���/S��$y>�x���bq�C�2ei?�>��j�.�4Y>�{�S��p��d%��*���� �7`d�U�܆�E3ӆ��߬� �����6ϥ�n�6�2�r���Rl؋�*���K��VT�A�U�))oX���2�I����J�IpR55{R�ت��(Ǜ8��I9�>S� �E����p/l}�"�B I�ٜ��Z�E��S?���ȺQ�ܩ�9v��!�Ogؒ?D�J֏ؔ�﷎W���P���&�������4�Ig��3����Y�ٛ�h��+#j��������=�!r����Y�BԽ�1(Ws^.�Uҋ�k6p%��~��z�宨��l���w�m��Ω��C0mʐD;E���X�v��b��w��I7����j�:�"ȗ�&�}^6�@�%A,�򣺉-M������Sk*�E���n�x��!
���j�B���!�~૿�E#��QS4&c+�*��?)�}���	��"�n�'xh�׋T.�Yã���+�n�Y&���+\��k��m	��ݝu�U������N�?�!2�'.�檼[�Q�b�x�,�u!xY��t[9�ʣGjи'�g�ӭ A���b?�ʸy��n�����%��/���Z�뜕]a(	¼��Ƶ�q���=~,���.U��)�h����X\�YX��
YR&��:/9��@z�<z�~k��
~���w��ީ�GĨZ���`���3�����ħ,vW�Y��o�0Y��JDTv@�eןO��@U$7�D����u'bf�
�#�M�u&���+�O*l����~oǂ:�Q9]㿡�I!b�&�#�.g a�ףtI�|	��F��~D`�
9n8�~3��ڒ6���&�4��c����9�$VJhY��vm@�o88��q�af_%�(�4$>�/"{wՍ�C[��6�֪S-��x���ig��=���8c1��1I���0�p�
nQ�-/��ۤ��G�0����;��M�'g�Y���a8��t;��b��f|�0�n
�\jڅmO��uA�|-�S�&�"��R��.�����&[�Q�m�J��R��&"�/y
�FWo.a��ۀ\�g�YY&�s!u��u�/(��X�%:M��]l�(n�K�N{Ɖ6��S}��=s�� J�1K�N�f���`�c��f�1�j�R<�!�{���,��P�����?9V��Homz�����(e͒��r,�ȅ����! O@��<?N�|Q�X4�s�r)3ྌ&�W!��&<T*��5+&@�6�0� �;K`�ů�1	.DC�ST���(uFmv���>��(�6����#U��.�רd�>�%L��҂;�=������ދfh�U�~�����ZM�Ӏ^3��G3�I:#�x�;��+�Y�� ^��ST� N&>⑲bI�VrMM��.!$i�B�=��Qh&��`\4q�?�����/�	ɪJ�:>�A,)�����JH%��J+'q�������ͫ�s:�q �%�d�bb{hT��ձ�M��Q?>4��;�<*x�eP���1�U���Un���H��"�i9$.?�xSU�l5	�ϖJ#�ɥϹ���m}(�B�`���)�������!��FiI�{�mǬ��a!��T���**yu���AS�);�]��?P/�bK�U%Q����+GR��f���_�R5�~����
�X�s��F�m�b�=�e��>��`6��Y?�y�{�͂�qm�����.��`�BU1ǌ�́����f@[���nK����.��3���������er
6Ѷ��	��1W;� 8��cS�*��-����?�
Ҭn�#T����N��'.�8��9�#����7:h\IO	v
�m٧��3WP��̽�6f���г�F����Y�f^���IM�Ĥ�?<Ӭ���=�Vq"���^���2`~&�s8��Z		�y],03��|%���Q2YW�Z���T���>�a�4�q;(�v� �N�����{�TnC_R�D�4+xQ�]��B�,��b%n��#u��-6�~���Fzn�=6��Yg=��R���w�CV���U6�\���{诓����.�����a�r�yL��OK�v�G����ΰ�},��nҢ� 4𪃾|��� ���IT���s�y8�2K4�ߏ!sc�E�{�gڬG��% ���+�XHZ[�	M;���u͚q�)>'l��=��)�IP����oF�8vڒ��#5�V�ꎤ��rt��T��%��dp��g�"�N)�d���{fh���ϳ�����
�?by� ]�da����o]��y�b�gTZ׼I?zSvbۨ�+G��nK�SOsÞ�S>���ٶ9���^�D������J�^s�ȎG�+���?�>�J �y�QǍ�.�0�x�u*�q��ȹ�t�N^�� �YFC�!��;獉�T&�PH������%�?��+^�F����0~�ѧq�w3�"ZD��A��h�"�2�8���r%A�'������+�w��f�H�%�ݫN\2{�Т^���+���j�+F�_�\���
��"�٭i�
�R6otN`R7��Ƴ�?�/�?���gC���B����6�D���Gni����è����u�I&��:����VE��c�AMɎ��슉�E&�����Z����w1����Ċ�
��`�B�|�)��O���%�ɲ.:�c'��5�L�5�Ih~4��V��R���[�1�c�b�WQ��gsk"O�šwW�'Ta�J�%�c��� �btk�������iΑ��i;!��֓<2���i.��G?ƛ���3���8Zw�#K:��:`j��:�� ���&�U��`yT��_hXr�����t��R�xH��ގe)g�@Tkf�j�C�|Nb!��_b ��O��g)L�����I6��^���oN�������ޜ�·	�x�VA������:��`:9��+Q��֍n1�	t�K,x ����h0�Zd8���W�+�4�Ŷ_��Z��uT�w()\NrY�N羦m�4ڢֱ������
e�yPK��2�BY�U|��KË���H/}Ӥ��1ȩH��P~��cl�WtA�*�@i@�iL]�$I�3S`~�[7]�-�W/�;T6|��q�Q���p���� �����c		��5�_�+�n�H�P�:�R�	T��H9}�vb��N&�����S�xU#Yvo�����SR�mT�m���Y���:|ǡ����+�"Ԫ�E���Q�nU�D�P�swM��r�z���Q!V_��b��,e��%��@�T���hX��U!�BE�{��E���ڙ�e����˛p�V���yN���5+RA��CK��P>� Hב�J���KQ�G�������o4�(�0�{K��5��0�t�^�<b*�m��&��6��w{��q��҉�}9�y��y�}�T|6���+dF�� )���f�+�[���!����{�0��A�B�hB;<�(��Q��h�H�)��=# 0D;�O�����<f����n8P�f�]�v;%�����_৬�q���2t~�*����/�?�#,k����p(��w�u]�,�-N%E-%U��f�m���\�ʖFN�ΐ���w�f�)�.~��H��^1��aA��h�N��h�g#��,����ncm>�$��F�#z� ��;�[�jh,;�1xtN����<.Ӏ����<�=g�nR߼d��n��&�	�7��!�a����v��}U�X)=]�Xg�M��zi՘�g�^|(�&�M��2`���x!����:. ����G4�J�]�o�.gޯ���:�|��Tb˭��T3���YMY�T��ߐ~�d�	&��_������#�W�������+�v���R�+*��75I�H�rt���=��x�kVl����x�x*)�+��b��q9{>��E��7cêvHzwI�F�SKCRc�y4�\�|�Oڗ�T�UD�yx|���(���)32w�J�OmNP��fȩV��s_gÕ"���"T��]Y:�*9}�(�
�[#�_����"�e�\D<�N�O;;>��]K{g�F�FUn??�.L<��cq��5n��ԥį��q����PTï8.�
��3��aߓ2��{R�6��g�X�\�-qFu(�����s��噛N���K�{��fLiW6��=�T�R��X�/��%TXS�4xNH�t��7$�6�i;�Tc6�����Z���m�
�B������Y߽宍+��o���(*��Ϋ�L�Qu�?�G��dTYf#YkOR�H	�f�2��\ 1�%�oj�d1�!;/}Φ�]�Q{�w Ǭղ�ЩHđ�K4�q�E��Q���wo�VQ0 j۾J%�����*,f��o7鑑i�mդ�	Iӏ���b�/Y���g�G�IQ��_'G3���*�z��@)��>�����B?�'���!G�JENI�ɸ��!Et�G��6�'#D��*���"��c��VE�YT��M���݃����ʆL�|�S�C} z�М�ra;�g�T�)���p@�s����v�V���wL���4�L(&�{��l��BJQ��gQ�^6�f�d �o_�ՂUE������ן�Ӹ�9�IiJ�<
�1ߩ�	.bq�i~�h�}1���՟��C-�<��Oŧ��s�U�;�Ar�F�q��j]ɸ��5��=�n��>EaP�:�@#������S���	<h�[�+�S\e-L���������Iʶ��HT.�4ggt���E��N"���h�؆����J�|�`�R彑����3
"Z��w�n�؊�)m*0�$a-V��CR3|�>W9��E�eɁ3L	w,�O|�WrU@?���<��Lq���f�B�FaH�E���n�t S�#KRcW����T�<�d���:z��]��>����x�������O1�!]D�� 95%X�u����z�q4�O�M:�)������7��w�$evP�&��CS��)I��E���+Hq��=gb�G�p��H��)(����fo�|�e�`Yl�D\�˕z{޼ق"��y|��X�f$rf2�����Yi	�P)w��
d7	�7y�87����A[>&8Y�8�J��77�xe���&���''ժ�Pz�VPW�Ɗ�kڍ��{���JXE ���A�#:)���<�]f
8�g��3�is�
7oS���Y���e�����kE�J�ѹ2������a
Og,�EMF��������'�9���P��Jś�d��b��1�_U�5��l�����D1�����"	������!K�c;ōӡ�z�<'�.��6J���me�-Ѓ��Ɇ7hV$���^@��w�p_)ey�Gֳ�p2�sRf����>��^��e��)�Ő�wǹm����� ���$Od�U!��i�Y���qU�Q��!p|3�?b����z��+��P�0w	�m��ʗ I�4��!�H��ރ���$���p�.���q�$��� �~
F�����("�_vs�ّ�/�,�ʝj#Q�K��H��F��t�m���HC�/&|����l���bL���*���Ȧ�VM�N,��Cg>��r4���)�TA��s��A��8���	>}

���kZ�C�� -�o��e��ǋ���%w��g31T��_���8sc���TX���G��/��Tw�,z0!���H"2��Mz����jL�o����]a�&)]�rN���Cx�d&�Z�q��T1%��暠E,a�Oֆ�7�	'�_T���"�͆�w�C�~�>�b���ծ��yuC�J�S���B���>�^V嫾ZO�@M_����^��T�TY�n4]}r�8 ���~G�O��G/3�Ƨ���������l'��@;�A�|���c���/cR��|�;AO��gm���x�X������ۊd9u�#�C§��}��'�뗨���8��H�?%��:=�\�;Z�_��T�)�j��,m����>��z����P�-8b��Q#*�{'�&u#����I��L�z|-ػ���0'xF_FaK���v�4R�{��X#=2�Iѐ�s ��Zs!=h��|��5TQWз�#�)�����~j�9���ӿ���9|�᯸póѽ���0d��ǄO��i��.����sI�ia��R��XX�$ֲ�7��_	��Sqb��_�]O����$��L��8�~����Ğ�Z�X{�ѥl���F���!���ǃ8s�_��}�p"aʈ�Gz���/����A��_�(����1���w�'F�Ҵ���%��rUfR��r�5����[��DO<��/[�A>	�,3Cp���X?7��jk9���`�M�i����K�4�3���TO�#�v�D��U�j~-`�����*ч��¶�sq�����5bq{�d��
G��U�+���~��ﱞc��t[z���P((�]�����[n��m��Ig�E�u2�lb�@1%/����7��9^��b��*��MzE9r�yxְR3�A��m\B�������Kڇ}��a`�5/�18׊��c8{�_p�{q�P�HN�])7Y8{`�#���0(�qS�<��7���GjiZ@:Z�u����39�\r�&�F%@��ֿB�佁2���o)�߆�w`�^�}����l;�*�:8�o����f	�9�$�$ ���3*���/2q����;��;_ (
�_���#����]J'�����&��p�"�E�K����T:�p��wP?A\u̓�2���G�c
�@�Ǹ�SY�:��A�� .���kD��zŮ�ھzj+����]��u�Q`#��`�';���!��{�G�3�Y� ѕ�="�����t>���x�-�CV0���Ԛ�~�"Uxu��}6ԟ�t��f�L0���*R���Zw߿W���p�e�����O��~�z�Cp��hO�����*n|�������\�#c2y��b��S��B)�#m�h0ߘB������N��W�����l��^]G�_Uw����)��	��_>7���j���&�{���T�z�纁䢕��ە[����7����0��~�"N��-y���脾� -Σ���z���v‵�w��#Ld��^s�+�+-��<� �����J 9ż�j�!��&8FD(�}��#���1�쮇Paee��kWVsqF5�xe�?p��j��Ũ@�L�fU��1Q��N-9WY)nN��bz 4��"��u-�%���=$��NV�>SNM�I��`�l�"��s��&�}$�8/��3R���Z ���`���k��貶�a�]��E <Q�5U�m���k��X63T�A!�=�>��J�=3>m�Ҭ�1>����vv�2@&?m�pA��F"%}�!�<��}3�N�إ,'}�T}=�W����]�ssY�Q�a��6�g%6��be�݋�yx�D����t��9,��q��x�DEv��:!%�c|��m>��Y�T���sd��Y�3I�%���5�ĘX�t�������G�'�,2���ޟ7=�2����=D��F�"w����ee�~۷��%�&7M㘺���ǃ_T?wƽ��`��=��`�ǣQ~��%k  �h5&3-�/����.�4�q��G�RQ�l'<��JV�=�����=�T{�ת o~smL���M��:8,^˻����=.���_����o�wdƜ����]Κ�xXuy���g�@��g=-�
�����l�j�Fh;���H�Z�0�"���9���1�ꏕ� !���Âu$�K�q�KL���#�/(��ۃ�X�W3-l�#�2ܘ�,��wΥD��	~5�S�Cg�ۺg�Ke�R�(ě�I	d�����&/ ,D�A�b�O��m���C��%�H�)��+����Ź^����{�S��D@i�jfG9��XC&�N���)�WūP�U&I�&���$�25&/�8�!�U��'p#�Ocr�R2������i�xи�a�8'A�g-#�8v1/zd#8
ԁ7���Q�V)���ِ\�b{W���h�M �4�n��E��Vj$��]^9�*� g�r���J�P}˺׬c��dq��e��D���:+�?B�������E F��W2kP+��w�EIl���"E� ����x,ǇkЇ+�џ�p,c�FNٶ��+�-�8v �xԧ�v��S�u��U͖���j�������6Z���8СU�/=��;���M��j��W=�����J�a�A|�o�A*�p�P���ƞ��/�ʭ(洢�,D�&Οh���i�c����� 6x�����6�ij$��cӾ�A�o@�V���Q��:�Oאv	9�v�m��3xN����:���x�F�+��N��b�e$Yυ9�vt���?j�O�����@�Ku�cP���0EՀ�n$+��#��w�Ŏy�f�3&L����@�lZ�a�I'K8Z�^��5{�r�O�cF!1��r��;[�cs�>��nR�I��y���U�[XQ ��G�%��dr���K7��7|+�i ��_��A�.�r8\z�[�&��]U�f�'�p��l���Ȅ�;�DC���f�\�Gs� [�9R�����A�����1s�k��@ʞ���֩W��>�7��s���n"��$�[�
�-u��̴�@��\�f�2���Q�ܿM�� �$��L�A Ea��]��(O3�Z����|-K�+Q �r��)T�*���D�"a�s9�hU��Sء؛���/~A�j�u0�Qi��U�8IA�*
�[�uA$-�9�ϓ2�9��@<`n�߾����m9�ߢX}�nan^Jt@)�LQˡ�L}�b��8^E3K�Z��^�;���j���[m9������%��=�.�i��y�Th8Sc��#�/ȑ�ʗ��D���G�Z)|e�/܊�>��/����5�r��9Vȋ��jde���ܜ1��;�}{1e��ס�V��ڬ���ečf���:�ӿ��9qUS}^��p �����Ӭ�&+����*MT �-��A��R̉}�g(ZN��ď�:78B�n��l�]�T\L6Y^ݣ4���ث�s���J{2p�0=#,.I�c�%޲o���(�ɛ�U�E9J����@ڃO�\������ۻ)-@�6F�MF3;�W�`0���օ��x)3:�Lue�g��qv�v�+j�N���9��H��\�k�1����\��.���{(ԅ"$cq�[�T�<u/����wh�J�Ҕn��g5ڗZ�I�y+)��-����DFv���[T�U�lM=\a#�v��u.�i�ɕ�ov���jz9��M�r⚪����\*�$� f��W�j�u�Q'Fa(^�&�ӻ��E�E=ژDNHE�B��f����.� >��q(è�!A�x��A�Q�|cd"�>
���^i|v��~�2��>�*m�f�#^�X���4?�qs�S��ٹH��j9obR�Ƿ�kc8����J�-��J�S}Z�WU�N��6�9���װʄY҉)�s���'���MK�\�5�Y�t����&���C�4Pu�Ǵ���
W���TҌk�$�s� �а/ߛqZ�ϩ����@o����-=�}gu3�~�i#OO��rA|h=����d?���m���n�]^a��"͟��#~5F�Îqe��w4%�@G�#�Ù�ʄRK&��&&~qNՖ���uŌ�]j�i\h|Qn�)�5���`����P�����T�7���W�Ш�]&�S��q40X �_/�2G��D��!C��"玫����@�
�f,�(�l�.����yRRd̋�	�*��<���aH������A���^2�r��(
]�Zy�K��������"��I?S=щ�� �R?����=�|4�|��]]�y��O�Vf�0E*�u�(!�|`n�
S��(\�\V��J�^����K����� ���m�B=$��.�cc��N'H|������0C�m�߄ +q���\��<�>�h���,$y��3�� �OD��e	�r�[�5�g�2��fOl�g��*��[\�E]-C��a�E��-p�>��3���՚QFc�8v&�)�dqRf������Qڔ�R��J[Y��U-Gos$�X�àrBOm��WP3�m�׋�37�Q%&��X�L�R\o�@!�<�g�V��v��~Dƙ�Cvg𤹤�����%����g{�k���6�����}N��VhH�
7�j��������s�#�27�����Vi�'V�����~ũ=:�H�>�B��j��!u ��&i�&����b&�vs�4�g3�IR�a����;6�c҇˻��/�'����wޔ���)��wQ� ���ϥ��m"P�G`{��v�'��`� �<w|�/����M�&(���K�6���L�	���l�3D�!� ���E���C���
��}�L�Uw����Ɏ�j,�Q���w���t=֗�:Q�θ�u�o� �S�R �$D;D�}Y~�}�(*	�� b�g�5Ȕ8��]W8	 �i�8�sb�:k=�f�������Je@(mʊ���I�'�U�.���?�OΖ?�D�o����7kf,��g����N���6�Pe��0��i�=_��y�%��p��Qe����͜L�5U3��z/OaO�`��/��^K�hA~~_^��wE�
JYF\�Hq����6�ջ��K��@d=����b��ke�w��G�� W;����e�z��i�G�;]����ilڪtY�w�CAax�Sǘ#���H�|q�8��$8 y}��ʑ��M�|�{��.r�۬m<�R�W�Po�����tִ���mo.��vٰ����C���*m��7�<����Q&�N,9��1A��/38���?����W�]��O�6O3BZ�Ȍ�ؤ~Y�y=NU�V��Tz�A�;3r'?X-�	���SX�h�3~�C���G���sRt��.��St8W�)��1k����!�VVcE�ىN�$Xh)�M�۱w���R��U5ﭦ�d��8P�E�{lO��b��pt:̖�G�ɳw�)v�ìݞo��m@c��t�B����o�����e�]]U���1���a[��h�Qs;An-I�z_8��_�n�E�@sTm͞��_���-���ӛ�M���w�R�ʤX&�?>��J�E���8A�L,
ig�}��>���Km��m��q;�`��������4����]հ",���`pH�ú��c�q�c��89��O;����؂�A8�t��@8�Q�٨ Mc/�d�iF�5���b�!�#:ӤI��o�w���^-���1�H��G�ZK�	��c*%�&��!ֺ~
q��׍�+���	�v4K|T�j^G2]��'��#Z'�z�)ߛ�n���`����<3�z,2M�90�6)���s��!�M��p��F�Mh�.�0��qnr�����ک�Ί����m�ٽ_�N�^�c7�!�f:�c`�r��з�51Q�EfoQ~KB1T��S�N�`�8��[����t/�����1��b{A�\TxJ]��;qˋ2X�_�?��"Jhz�]�e��s� �q�1��x�uŗ�w��ɤ�v�.��g��z]DKw�__���O3J��>D�����.��ը	��0aR���P��\���������OL�f1!�L��8e�ƕe�=Vq�0�	ª��ZL�Ъ�n;�ևȐr~��!�ϖ�a�]��/~a�'�ݝo�r�?�&�7׆���6����G���/�J�z���$������AB��(�00�q�Z��[[ }5���?�����3Y�A���?`��S�6V�|��r9���%���y���f�Qh�9d7�4?!�s�@�B����Ka&�6�n�-����6�D�[�UK��t�dy���yN��þR�Ca��/ӥh��7,+�0 s����ˠE�^��=�����GT�:>m
6��B�m�����mQ�t��c�C6<���)m��C�Տ�%L)k���Fq`X�����Z�b�j �<Э�z�'P��	R��:�쥣5��ނ*b��a�dY�a�d��Z���W���B����0+��햣���_�{�5H�gZ�5����?f��~	��q�|��n��w:�)~v ։�vK��q��ec�%as}q�����)�YDf=���NE;�۳��<�f�E�Ɖ�x���r�^.��_�4D��$I�u~R�~R����g�+c��n k>�h�T�j,S)e˒��%?������l�=FI�2�>'�e����M���%��TR�gO˔fT8'��{I�����N�a�ouA��l�Fd��%���Gz���=����Q��;�����y6ء��I���-;���~'�<��]��6(@[.�i{�ũm ��~m	v��V��;�e2i������	$W*hx	�Z�N��9o�JB$Y�=;14dD�$�Z���h��;TI{B��*�`��X�;s��K��m�!�^�ܘg�@�>�9���邊Dd�E�lI�^ٝכ�5qP�9Y���3�,k��/���sz!���N�f�LDB� k���^~�=`��ܳ�ʫ��n �����H�;�$�����nd�t
��g�����G�7�Ҕ�>y���v�=�=�,ǟ�mVO����̧�5����;��2�я��!\|��
A�ҋ�˞�����Kg����,08Fƪ�ދS��R8ͭ��8�]�?D
�x�x0��j�j@�s�I0V#UCq$�o�h����%Ǯ�.�e8MbF�)6�C$Zj	����F��ҾJ{�m�� �@j5R�r�5�떟��-��_qז3�����B�1�ۻ��y�}ь,%�2�{��cҳIQ�X���.f9Ö��թƣ�g?���M#5U/���;ʺ�@�����\7�S�AElۃ�G$���
�5�Z����y�U|����7��!���L)$�X�L����7,t�����"�c5v�iV�B�nqZ�-�%C����]�'ڋH�4�>���Mx'���֝��q�̳G�L��1 �o�`�?h\J�Rp��FћW"e��i��
��r�ÎeWP����d4�&(�`G��T�;�@��~^�5�}zq�8TM]jך�����[�ᡮrD���Z�H(��n��3ҫք}���T�5)�d���q���H����*�?���g1EV��Uȭ~�@�u��W��U��v�E�T(٥T�Yk?d��š��g��wgʼ�c���XўN�].y[B��7�L�ɛ+R���=Z!��k���m&kV0��u��K�]�k�7I|�ߣ
6q�Ĳ���,[Nmd�"rXw����'�6��r	/��݆M�a��݂M.9�E�=h�[�U���Č48��p�p��{�W� �O.Qt+s���Th=�	�u��9ǧ�)���Z���p�Z�jb�]5��qh�a�B�BGaX5p��� ������:x��*��g�������oZ@�A���iC����AVo;W���} �=�/�i,��C�Z(�J�Ie�n���>�����3��}h�jWPw2�s�#��샧���8�'��l�8���#�1�2���&x���a&W�:�Gܕ����Q���85�:u]�%�>&>�� "o$!�d��R�Ø|�M��*s�����̀�A���-�&�b�����M�p q�ӇT;��Ud��>q���y�tn��M�������/���v�ʭ��	qrp�9eV!E:v�BOj?Ɠ�7׶��d��\5��h�j�OnɄ�"�RX��+h������]/R���pkQo[Z���a�=0�ò1FPy��ጁ^;�� uY����e���Z����8�����?�j��9�����<>��x�G�I޳� 7�%	�q��������>��?~o�U�w	�$��E�u	?�Sȣ�����
�nVׅ��� N
��LQ�鋁��G� �:���z�Sm8��#��2��a
��/�%,iY7�Q�t+/Ɗ;4���TCKڣ��z�|An[���$���L�5������hɣvC{��,P%�W��~{����s"TGl�˿Oh��9�-�=��m�y�q:Ӂ�Q ��7�f\zQ>
L���T�%WH�8J�������5��RXf�Ky=T�ܙ������K\�qq6�����tL�5[�q�����/�~t�����Bbp5�3$0�9�u���������)t����4(�\M[�8�����1qD����jDQ����+�Ձ���ͨ���*�ŗ�|�48�NZ�i�����]G�p��Tq[,�3	��4��h7����h�ѤO�Z^`�LV$#o)���� n�?�4_}��mB];���*���@�WA����oV�.M2�8}���D� ��F{��#V��S%5L�����}����LJhS�0����š\����E��:��rc�t�4b_2��ϙ�C�B]a��&�X��'cU{�d�a�O��π,EF��w���m��)k�8l@s��x�,��H�Ѧ��+i	�X���F����`}D���N	:	��	ֹ��Ci���;�F��;�Mމ�<(m¼�#��6g/!k�`zsay�.EY��V���v���ȸk�dYɝ.�}PFw5ͷru��뷯�qz�)�������+�c�VIAZ�p���7�'X$��^�ذ&#��l�Y}C~�}a��^�ot=��,�E§qg�)��v�����Snk���:R-,7�	|C2����s.qV#y9��z�N±��^+ߥ�qjf"A�Y
�{��f��5@�,3���̿���0:`a�Lai��'ڿ5��m�r�?�o7ֲ ��|*B��J��K/�.u����`	�n�w�����m�����i怨� ���eJȹbXQ�/�#�bgXBcZ5t�8����R��u_���Ult��S�dcg�st8ic^f�䫝�i�f��3�����ƅ� 
��*��f��=D<0�H͏%�:��÷�^�(	�tZ��1�l^�>���~{|0SM�
�ۛq�-y'���1�2�V�(�9Qљ:3� 5�[W�Z�r(�*Ef���D���d]J|ʯ �H��i���I�7djb���x�I�}�b�ǂ�s0Ǚ.��/r�.�7���[&|�� ��X��[��_�ŗ�A�V�˽ X�C�b�П��<��7eqoѡ�b�϶sJ<�1
�}B�#�U��ta��u�BC�+��^�����J�5��g�;�)D����y;����f=1L��@/X�b��H �*�0(�#�����2�+���N7W�=���>^�A�$z�;.�=Fq�:�f��vܘ>ׁ����^�(��N���c��9I����n�j�����<��%Q��=�R�$��;���楶6|��s&7B�*��/�~�_�B 8Kn�U����j�S�X��_��x��`S+�W�_����,t��Y*��c��u�Xh2|j{�[f"�Ѻ�K��=�������Y�`��ʋrZ��9͒LY��0�T|F�i��B�&5KP�уe
��@����;���!��]�|�DO�Ѡ��~�?l{����{���� �j���	��<]�N���Gѝ�+���+��1�'ؕ���j����5�}l�*��?F��L�����S��7$au����3��<��\�����Q㔦}P�\T�}��O�����ϥu�L��ɉ��!��^�]�e���z��]Wl�<��r��G9eVE��9�ɺ�(ioH��e 7�O�)u�P+���0a��`eR�`�J�Z�M,:�(ć��\`���J��]/QQ�kupDѼ�O]��'��� ���LL�O�Bb|�!Q��[.[�)'w� _v�SE�8���ǌV��Oy�{�t�b��GǊnegB�w%�:ݩ"UJ������E��=�\!���4��m�q6�.XfzxtUikqG~Gޝ#�t=�P�@���הּp��쨜�#�!p�N�b�$��
N���x]D�T�'�Pt"ܙ`�b�0��b󔢁S�;#߰&��d�K��l�Ќ���J�B{w�x�Sq�f�d��(T�6?mL6N��Ǉ9��>���)��ɷ��8/o�M�Nǿ�:d�Uj�������?Q+(�\�o�;mt~J1M>O�"�����VebO��� |�͂�닁f��×C L)'�՝V`nT���s�Gl��/�#%p7��O��n�o�{��7{��xff��rp9�����$���!W�o�a�My/��|�C/��jϵ��n��_���|� ���oOd�����H����s(�Q�����E�������v}��"����fL�+��Jw�6
	!����>����pa~����N�Q  *z_�y (���݆W�V�gC���'�t���J��û`��-5-4�SJ2�t��m��k��*d|�<����h��%��Ol�T� ���s@	n�	��kQ����UeK*	� L�3��=�e�K(i���6B}�V���[	܀�����]��('3��(�;�0�v$x�x���ֽB&-�/1�覉��Kv�N)B�^�Dշ��p=���.�2�oHs��nk��MrqQ�(�?L�0�:BfJ�r��%*�)���B������Mvd���ط�iv:�
�� �eC�y �&s2�*D{�-g���n9��N龧�4g=�Sl��"sM�û�ھ9�M�yY���tΫ��"���c+�a*ΚF���VF����%�1RWu:�� ��	�������m��DV<���Ě�;2h��,�I�}������$_���	<<�"`�7a�� u��KU����9C���e��a�jۣ8�\�#�w�����T&*�G_{��<&�t���K�Hsp�����N²-Y�[��l�,D�a��R��eU���h��2s�BI���U����?#���e��AN �@O��K�V�
p2�nD��f�ݴ��a�[�-̏�ַWZ�4~����W݌d�,աd�rӡq�^34��{��/&�
�j׊��̶ˊ������yJ<1;�eE�-��;��q�:؅�>���ٗ�x��W�b���S#J��7͹#dQ�&ӜѸ-n�B��W��!��a��ķ=�o��E[,�1��1.Q����ge-�+濩^%Z���B�8T�~����+�]�n������^����,������+rz �4�)���Cu��"��K���Ր����t��ۈ��?/P�#ŷJX¤1I��{�<�b8�]��(35�+4[��P�(lOW)���#[̖���f�n5��b�m�C�r�6�UqAw�Ժ��_�tAf�?ֲ��� i�.ԧ`��ׁ�wqC��P\>@yl�b$��3��,¼���)�/i5J�dde_�|�z���׋֢��W��Jt�N�2�H.���N����.�nF�;���&���������X��u��̗l8z�>G�@O���"̹��$'������k0Nե�x���]��V�j]2�����W���iL���iC��K��d����N�;y��H�ٿQV���p��$e�������k��;��Pf}܃u��	;�ֿ�l�&b�[�%��ۢ�-���Ψ����jf��x�a�Z>�Q��H����K��|���������S��U�Nt�����>�m0:�s�Z�#�<��:��ǶZ΄��:~�^��\�_�c�W�_�[Μ���u�g�TeE�?5<f����?�-p 3y�$�#��˜���d��-LO�n��M���e��+ő�v�j�0u����}*�|b\¡N4��E��%0 C���e]	pq24~����:�)��h
�P���ïq�/��tEAo�աvA��;
�8�MZD�<���{���S�<4�P�r���l�!P���K0��oΣ�A�[y>�Z�-� �4�5Ȕ\�Wg�qF説{�`��ң�Դ��dT�)=�q�\�J�F�ث�\�ŀ=��)y�(_���Ff��9�eG�ٯ��n�J�%t��G�����夙#�5�JUHw�r2��ƀ��fR�!H���4a��I��R*�{�l��m�$��*~M���Xfa�ԫ���+M
���if���)v(<�����Z�JK�LD5�7���`��;c+}T�w�M����g�1�
oR6�"��=^Ƈ�9yѸ����~DI�K�K��n2�+�9P/Ol��2rX�ߪ�Fs����6���xGM�|3M�+��eo8�d��g�HI��`�|�4��]���[{����_QE��E?կ���m��'�q�`�W��%S����F�VÌ��`aq�~+���i21 �_]�����Y�Ϯj��Z7'�rz�d�KY:đV�_4;�r�z�x��p�^�f�n�	+*	�^d���Պ��	�Xkj�֦���@U:P�r�
y���n�~�Io6�22iuY;�do�]z~��m��s�q"U�tM̋�����T!jW5挖&ёϏ�<�[Y(�+���<�G��x'V��}�7�|���$�:*��l�	�#��<�A�����6"�&���J/$/y�P6�W�@I"Ή�%uJ]4Џ*����	JsZ���ۯ��b��x]�R���J8E#��Q��B�� RCQ��E����w}��/�MKƒ���Dy�F�Oɭ�<���u��H�4�5�h��k�\���Wq��F򥯌�%/� �!���hE�9ÄC���M��3?9�^�y�T*:)���`>�hQ+�qY�_C�o_-�:�/ �{A���_����˷�y�x���X�P|2T�s��tG���u
6���4�#�'�ٟh�db�p����v*.a�eB[�Ƙ��ݦ�۟/Π��NK�X�ʠ��y`W\J��aY��1`���G5or��҉�&��k�@fzaW ���'am���b�J�S~uL�I��j�bsd���[��f�E���{/H����	�%�0��U��xq��Hr����`�b�p]ô?��f
3xv��AA�>������]�f���>W� �a"~�0��g��I�$��C�`~����SzjZ�UF�Oҙ�?�Z���� �M��m��PQ��c���<�}�wY�ż��%�[jKE�%����Ce2Q��^r"�]�L��܎�6c��!� Z"[�cJ���U`|);���������T��W�d�E]I:��! y;j���QE�O'H}�G(B��+��� Z�pv
Y�
�f���4�;.A�pg�t��������cuEr)��Qp�0�n2�tί�3{�,�ic'9�0���%�/�f]�5D(�6wcª�h���0�*YB�	V���^g-Y�5���W[s���P���X�@A�Ҭ>��Q�*�0�I1�0�S8���a�v*��W�9��/�yt?Se�3�,x��ϰ��'T����熔0�{���`�N�W���^9��cA@.��۵jy�:n�@.aEh��D�?{Mʯ��<ujm���b��c��J�Y>i�v�m��,8�$*Ja�p���"����$�4�/���JƖ�c_��p� �F�/�[�����RBS ����
�*���~��(�{����w�Z�Q��ðڑϪtmrN���R��+qQ��C0�W����@�c$i�7�ّ�EQ�a:8��|\�vnIv�&�E�'��{�	Y ��5I�f3v�5\��mA��	"�m��3%XЍOl*�q�N���y4E���6Q�R��G0��RM��d�M-XEh�#��֪DW`���e�}�������1w[Y-�FagU�U�'�8�[V��[;��g�]����JY�@%��Y�=6	�UɅ$ ���U9:'3���䟀�����f�4&���Y#|�%�UUSqI�E�)�r�f͔$[>4d�e6Ž�Z��D�n=B���Z�ث����D�@�IZ�8��.o��F�90�)�a��l�%� �4�2�%��>�^�V���
�W��ե�W�$��M�����ۿ�k�:���91#뾈��1Dr]nI�?�s젦�k�� c-� ��*U��\h��2�亘O���J4~��X�r'w3|S��",���9�j�)o�(&x�Ǧ�pR�lI�񰡐4>u�R�m|��']�V��k^�P�$���ʹP�0���+�
�!�g�YV���A��4�r�J��wEq�*�%Q�[�"�*HP0��>� {@�׿���+��?~@$�@�b�S��Ji��Z�M^�=�T�ү�֧�
���J������`��rH�)�[��G�!cY�#��doӧ�w�����?�b�р��6���$������r�ԏ���5ǝlM���d���ݽ�0����QD����t�$*���)�a�"!��.�+`�S �m����/@�_C�	єik�az�&��m��4��G��t�#�Y��Ӑ�)��Tۦ)�zF,��P�D�t��j���5�*;^ڐ��X������v��E��a�&���	{��;{�,�j�v��і���I��1���jQ�K�~��T:�q��}�F4&pNA�c)�1��2��xnV�\�eEp�n?j8��m�·5H=�P*��@L�f~� �f�X��x�W�	�����۟��-!~�V
u\F?���R���d��'h�w��m��h��W9�����w���HV�Ҩ��^��M���W�i����1�W�#k��@�2������Tȶ�Bd���$�ZY���EQh����X�r� QM�3�鯡lC����c��ș����u�=�l��+o(��W����74�޲]�38 MFsTU��$��KՃ��I�
�8%��vɒ�����a�*�y��
:v�������+8ApW�f�F�ݠKU$�����R�K��"�Ҡ6��1긅���K��;
��!��,�`��e��]����C�k���{�"���tG*h���7S�;��%�'i9uh@�00pT��� �G��%ISZcp���G��3����n���eP۾7��b��B�M�$��Ϊ�]�J֞��_�Ҳ�QEk#�$�+����6x
U���x�kztz�a�<وIқ�3z���! A����n\Lv���o����\.�a�.!7�a/�Л.��u�i������c`
���X�=n]���X�������L�o)=�;��~u�2� �n�X��z�ڡ���wC/gAYpD�C����k����kHANR�3��}��@����;T@�=��t9�m5���Mc6	�6mY���S����[���)(��A%�nV�U�+y���\���r4����[;EGؔ�e۾�c���N�s����M�D���Jt����%t	JZ�@�q�G�U2��q�i�M�S`������9��!PVp��\1�F�?��ӧ}���D1A��R@cv�����@��MsP��rUT����2�� <�x�ר��3��1���tL��?/�%<�t.�7X�dA�o�0�Mq�(�L�þ��rՃ|�ƶE#���T��%�{R�>�lm��F20Y����n��Yr�[�;<g4�aQ:�?^_���r	|v� ����&.�*�l����M�
J����5$��ŪSq���X(~�#3���tN�?@d��ە�f`�$(�y�w��f�[4�dO�N��$�I��O����g��T(�썋��_i]�"��F��,����*7("4�m1�O�����T�"~c��yڨ�ͅHr�=!Z�uИ@�PR?�)��'
a [�eg������������뀺��H�-�w3Y� ���ŭ*:l���/d	����e�ON/�Oއ��4�o]����N�Q��@a�i/�?M�ѵ�H���Y�/��d��)	�+p�9\4�f&��f�;��!3�_�pn1\�eOF<a�M1�Ғ���N��nu�Y�(�I�m�j�ɬht����4��������;?kԕ`pZ�� ��qߥV���Z�u΅Hv�;轆8�t;s��8_�_��L&���T��<�6�;�S��������U^|������5�D�tB�Ʃ"��*��"Hs�-+F1B �8��!�7����� �ᤡ}s���e�Ƅ1��s9\�o�]5�@�9��:���X�i%��qo���g�l��Hz��v"|@L����qKC�׈�,�KMx���  ׿� �#�����uᑫO0�'��#��bǯDb�%WmJ��cmx�`���ΓӰ����	�`��I�e�v��#�P�e�<̘���|y|p�P])���b��ޫ�[B�P�M�|a����ܱA�R�x<;�[��G.�<Ve(NJp��N��l�xb���?D�a�a2��`�]�wʗ�Κ�J@!W�&�%79��}�sy��o�z�V�@GVB6���2�NS]�d��1k�e�
G��W�夘�<��IW��9�d���M��`�7|ʵ(6q���cRN���k�gRl��8��a�n.���R*)} ���˂9�+���������0�ތv7�R�����#�R��=Tf�}�w3uג��Z�|Yh/�/$���@��?�
�ܛ�Y@3�/j%�ܤ�5Tȴb4���� ����e��~�E�5�'ڐ����r�36S)-�c�|f�����n�f��H�#��]��๙7��G�B���葋ʴ[,�g�Έ0t�O�Ц���d���NT���75�\A�8���\O��� �"��V�)�z��B�Aj�bI�"ɾ�qj�s�{�뼞d(����>���H̓�讂�y4j��%t�쭩��p����޲v
�+o�^ AQ�0F�LI
-W_-���Q��ܴ��a��|��f�o�p_�3�pu���e.F��;$S^���	�9jLʝ0:<@���V�ڃ��ӑ "��=ɼr8}SQRAF	�M�����ѝ�O��Y�W�v#oU[�>���/��kL�>b�J/��r8����_ps��C{-O�|r�7�Jng@�^L���9O>��>�}#?Yϩ}�?�S�\�u��]��S�����R�A��|�%��	�$r�X�m\ta*��$�MN{8Y;ڊ��WF)��8d����c�x�Ɛ<ٓ�y��uhG�~3���KlO��7`��Ѧ��K��I����j��Q�6�qB�����q��ՙ'v�O8%X�,�0��;�D�F�%�y0��!5!z1���5�ϙ�ڐ���`�QB�I�s�O'��	 lE�j)����}��N{j0S�7p���N�9I��*��>����uRm����@�]g���{��
N�ònnn��]�Ѧ�Mo��p�	��׿  �5tdT�.tR=�w�90�[�ą�I���m�r���+�N��ȿ:̉Gǒ٫�ry��{CW�Nw��]�a�<V���Znx�ע��7~��,�n�����E$�?��c.0�h[�=f��̧��M�e�{��W8��`���@�(0PcqP⻨GD�,�M�O����\~����������I��􎟩)����3�G���fL�㫲�ZT<Ea|��&�
n]��k�5p�p�� "7-G�}��Ј`�2�ѱ%�=����!�Wƺ�w(Z���?�mug2��q_�=jԡ�����7*+�U�4436c�8m�l��5g��C�?�Na��h��(���F�g��I�>�U���+����uB�l��%�k���:l�K�݆*�|u	� ^Z9�	�E(>�őn'yU�d�P��[R���?x�q�o>$�D�)}�7%S{����,*H��_g��Q������b:s �@M�W&
�OY>f�{���Y��A��$J�}��8������XN�>t����iٟl�M���e������Z�u}a�)}��,7y��8�
��WX�p��ڛX�4�-(�LS���� AnjK�(�����Wp׎Y �Ӓ2�>j,��0�.� S�A��pl����٩������ӽ����cV��5����"���	=������Z��cD�`�t2�i]ב���~��@�>,0k�||ˎ���T��w���`����"��8�d�o�%��<:	��D�H�}�!����d�'���(�ԃ���� ��-h�`CK��w/�c��:����7򊭇V'8S!n�"1a��<Y�Tp%"�k�̰K�`MtB6:zrWn xtz�&��L8.�������ʜ������E�+����LO�E	�I4\���fr�!�\��_�x���YD�i$�l:La�VCU=�8T^�VJq� �Q��N��t&d�v��S}�5.ٰ��/��O�����Wp�w�/.���Zqj�%o�w)\:�Ѱ��ܞ�tCx��ِf��}�\p��]���V�Ǻ��|�O��XZ��~����m�q��='���y�4���x�Tn�.v�}�l��Ԑ������`�K�w�+��R�&�?3}�L}�$9ۮ�
��l��@���i��YI7^5�|�vَ��9�FR��q�<k -�^3*�jk1�kjP�C!
�gy��gmI ��@f��:��K�1�\cC,q�5�h�ao�������x?�bPw� %,[SyrԂ�F���S4m�u��[��0Q}�=<B��΢�C���ö��*`8_Pb���O�q��\��G���u{b��Ύ2��&�K�?�2����h�gbS%qE�Oa�zx�BB�R�v��H�>�6+S$�y�"��c��u��9�ixie�'�(S��a��m�@�6O��G���l��%��3lQ�Yoͧ�vAyO��"}�_95ݥ��ә�!I����)��,��w㊚项r �}y;��J�/�,'� Rm���L)"	��_j"}��Һr�7\�:J��i�(�[���F=�4�d��������aٱ��~�ޘߺ]�)�M�Mu(��_�T$��lNdm��YU�ZU/�~�s!s�kGQ*:d-���כ�7��֍����N-�Ъ��(Q*����~��mɠiŰZ�(�.�
�
��y:�@8�؆�����s�X�u�+��	�W�ǣz���U�k���l=>�69_�	o�:�8����s���sqR�^t����a���V{w"&Y6�U T5�>�'��f��x�ǿ����S���@�������^�ڍh�L���bn� �Y%^f���r�q-,=H\�Z�QcU<�À�j��lw�:�T���SsWd�D��M��nb�B�=ď�S�ڳ�΍���V����G���Ų])1�~nw��s��1g���D�d�WR�ˏL��^Z�((��k҅����Xo)��C�ww�?59f5/��D���9��G���P;M�d�:"懙Ӵ?�`o��8��ԅc%�:�1�.�L(��l�<����A�@_�t��jR��Ŀ��V~ћ ����N�/�=;�~Lw�FQ˓��uw�J���+�|%�,�ڄ���JW����������H9���t�T$^����p%�,�Dص�1��.����������#�,Ih  z�['�	ne=۩�e^#CY�Fr�Atړ��ܙ}x�!{͢�Q ����;��2��
�!U\5"������o(�7w�u!��ڬ�Ȉ
SD~t'x���FCF'�t0Ljs\���y)S�Do [�$���&\z,k
��X�Z1���� l9�ԌM	���t�QF;.V�rS���qЅL�#p/B���2d�Fn����)J������T&�I�h�>�7J���<�2RG/ݘA
>��:�w\A�M@Zm�󧬆Ј�ux�L�:�[[J�V��� mPG;��ȅ��+��e�˩�Z^y��V4*2ޭ>�C���0J����U��4x�f�� b,��F8��+E���8H�<F|�c&��@d�W�W�"�~1(���A%� ,�f܆Z}qRC;��|Z=����M�n��)��*�:ڈ���A�t��X�9��Pـ�,�{�,��-Aj�N��l0�������FvA�|�u9�k*?jM?�IZ���9Y��{v�'����R�8%i��ь��<g���3+W�%5��^���� a&{��V�f$`ߢQ�TʏVE�/kO,�P�j^���)�d�q�!+E���6��A���C�6��gmdu@��kX^=�\҆�j��h�=6����[�X]����8]��$V�4`U�H~��������G����$syQ�`%�ϸ8v�	b���Ī��E^H�;�_�%b���0�s�箭����=�Ƶ��8��k�µ2.��~A�t��U� �Z��η'F��)}���@-}�����7!_��I9��N|������4�(C��0D+)-땯M۞��&s��7D~O�E�S�g瑩O9l}�eѠ!��:�$��r�7�׍=���'4�M��E�P�a'�"�y���B���<��Hs�ܸJ:\<'$���gP���ت��[����ivـ����gͻLIhP��X��T�7��Q���J�)���+]�w��A�Gي5�L�n�� հ"�|�/�q~�h�B[�5�ZO�:��fQ?�z�PF�ڍ����4�{�;��5G�[Uf��v|��W^�k�#L����,Q���z�U���Dд`�SY�xHSP1�՟u����S��[�����U%��*�����t���W�^'N�J"㼴z�-5x |e�>��Ū�JR�(M�ɝ�i�^�])G=6���uȚ"��UH���x�I�����:x,���&�w�#���Q�����6����M�2�,[�� (T���;+���8q�l��W���qu��~2}qE��5��q��K�d-���]������P�!���/�C�q�w��B�-g ��d�j�?��I$i�,����'Zw�0�"@PE*ڧ  O(@3�k_ŀ�j;"P���F�.[(r����X�us]�Iu,���2y�n@LM w\�\v#��CD��+�	?QM� Ó��
��ߓ����/�� kB�満��9��%��:� bN/���u�]tL�;m@��f�Ke\%���S��NgT������$��id���Q":=�x2�����a'����1�����*��m��uˢ���A�;��>-��4n����j��)8�=���ظS�
��^�R_�[�MCw�讻4���^{��
^9<���w/ҟ����+�W���i�[�u�<�Ah)�.�NօC���1Ac��J�X�]���V&�ˀjW�]x��>1��ۇ]�5D?�d�X��>Lz�5i�ZxH46��om_�ck�t9}��v�3�s�v*ks�����
xKy������(O��5	���#� ��G�v�=bSg�ZʆX�E]#�z�K\�����ǜQ�*�y�V�y�W�!BN�i7����N.��*X9�����v3��u�W:��S�0��Ƥ'Y���������u�ԳI
�^�a<� Ɋ5�=	�ijC��v���p	˫�|�>>w�БP��T�^�Q�w�
��x�
���H�}�@�L:%���}�mQ�vM�f��4�I��8ؓ�hd�oA��|������%���t��W�Ħ�Y˂T�p�^���s�:���Eq��b����I��>������na�q;�S�o����[�&���^���ŏ�+�� (Vd&?���&�K`�f��U�L(�������Ì{hj�e]9�@&������Ijh&�S��:q%Af�) ��>�5���5�:&��fӔI���S݆1j������6��UI{>�h8�F=H"쟋���A�+�	��f:eAbT%�2"����,���357����;�W��$ړj��HDA�q��8���p�X���aP-�k��}Q� �f���'���_r�5`��iz���V��T"�Q�hkHڙ_�0V��'� ϛ�cⴱgH���cI�$�,ii(��h�Mo������%�/�a��z���A/F���1Q�bh�|K�_B�D�V�9�C��HV�� 9���NWz�Ӫ�t���CR�7�3]��I��(	j�~?	��,Q�	��6�u�*U:��Z0��^�Gh?���) ��\��O�e��y�`�(�
�\/��:�X9�;��>e�&�B�<(aW�Bc>����W��|���%[n}J�	����<H�w�"���4���*��}⚄�#Õ`p�Pnj�I= V4�sZ�us������b]7�6eH<�B/��m�� ��#C-��x�R��D�h�.���>��Q�!霓B�K�C������0�./�~�8s��W� R�!���-�PFl7O��A�G�֙�Etc{�`�"�ܐ
��L��Θ��ɩ�������� �b�&MǽK����MS �7��C��	F�!�+�t
>x9��_�����mF���Xx�,үA����4c4�{�vGI$�f��xT��b��Ñ����*�ߓ&c�^�(��`o���/:%+٠�7^u�isq�r*Zjs+�Zx.�#4 ��7C�������C	r6���,��|ߩe����	�ׇë�:��~�h�p��x�D[�Inr�>A���O� �=�sY���%W�P�%��72��{���+�nJh��e��,|C�c�,�a��m��v��9�?�^#��=C�+>�foSn.��)!0�2�ɳ�#@�|y��@�N��<�;(ܑ��+=�/���x�J[e�>ul{M�X,�	
<���<'�k@��[6[2	�����<gHZ�bf�'�ONO�iH�i���բ7���6?qj.|��Q�;x���Xj��0� {��)F�|Y8��Ĺ���>m̋H-�j����fK��ԒSA�	�m�;8DE���H�t?��؜Iݭ�5�S�#�ԅ���Ԣޛ2 �R��㝿�(�T��V�<Q������:h+)��<Y;��d6;�Ǆ�l_gLS�#~����J�Q��M=�~�\�y�O�_7)�3������l�����~T|��u�8��:�4�Y9�=ҩu���uJ�V ��g��Ӑ�b��� ��vCɗp�W��`�1Gb�;���J���Y��3���F_��q�Y�Ȼk0�dHEA+�w혉x>�
�^��%�$Ȫ��xn�A����p���ʥ���v���zU�e������E1^���7�t�m�����	{��RD�s��b6�D��j�w�"�:��[Jw�m���L�^Lfnm�*��,�NY#D�W�҅M6�	�p�}��n�-�3dO8ALF<�q@0Z��DZ�m8���k�g�q�����R��`X�< è���Q�Sz�zڳ�l�"� ����D)Tm�s]�x{�X��e�������D:�c���z��YJ�7}�cW�d����ɭ̽�b*�[k#���W;RQn9��:d�p�������4��h��
�x���CbEo81���C��X�0r�ڔ�V\�=�p�P@�M*�P$�Rwc�u?|���B v�f��Ď��XQ����e��(�f3��$j������W6P�}.U���2��[_v�rH���m��yP����q�Ȓm��6�kH#�F��1��v%&����D|� ǸIS�{�}0E�H�rGX��'C�	_�VӯM���h�i�i^3Bꩩ��_��P���m���$D��%OyχT8.SBViQ=Uu	�!`������9�w�3����t����I�y�)�w4�:q��s.�g�����~,e-{08j"FO[�o0ITaN�5e�6tv�~M�����O6�{���Q�#Z������ �]�"r[�\��b�2���$G��X�D���^/ w3lg�^]a��!�/~����3'����~'D�B�2�f� |��CS��}��{��/Uoo��	 �����)-�f�V���q��:��T���Ə���"[X8��s��6:���4	�Q-U��3ذ������55�1��S�z���-b�|s�֞�\��53N����6Sk~���im��L�?���1�)��b+��y��9��UО� b�,�pM]��9XS[.;�m�� �j�����d�z��8��"X��$۞�_��R�n\�l���2#À�Ct�0��x� B(r��>�}�/x�l���4�哨�h�tq����#��m����f��JϾ9	D�����qҿ�4�G��*���{<�nE٘]�D���,�P}P!5����:�>���"��5��I큄�֬�E5�H��l��͆�K��J
�� ��GԤ��_2\[�1ʂI����[��~�5�O�"t�~�=��O~>���=�����T#V�#�~{���Z�v�����M�e�؝��2�`��_�����tMA�n�nQh�H�R�n��Fk�E������'�ͥ���̚�7^��d����pÍ��kH�_�i�:�
����u�^?RZHA��o����zb�IY�oQ����/k��@�R�j�ѥ���s+����׶yv�/�Ǖ��c;�����|5�O0��L����������2 y�]�HW1	�;�r�L =�,�+��eO�����:��d�-�I Q1@�C��$E-XƙDP(�^�H���2~��D���%W[��H��#	�PV��X2V�|_5�q���l�ā��>Z���.�籡�ğ�e_����u��۞��Kx	�e�4J=ਬ�:/zCX�\h�F�Ђ��-8LS��ʴ�(��+o@����_m�ð�n�0PB��?jF���N�¯��C���"��9�N.�qw+�*|)�ʫ[�U� �=�%�\���	ޱ�/���HÌK�/��*w�G⒢��(�< �!�N�PV�յ|�de�|��U���� ����H���`&>q~�F(�ïp���uv$YC� 5,lQ�%_3�]��"�T3u��w���s�-޾N1SQ�gm;�N�CdG1���t'�������Y�]��\:�",���}�̄��tN���M�|�ߖ��4�y��g���ɹe5���㉷�m��3� ��sL�ċ�v\��EU��K�\��@�c�xA�_�/N��m��X�p�w��@�ңy��(�[�#J!�����ɕW֍��}��s8M�=p������/��R���0��m�=Xٶ]�_%�=�"����ر&zԏI�?9U�`��5Xh<D��5J�7`��ݣ����KH�F�ϭаyWY���1��y��I��_{22&��Y+�����
������B���eK��@ҷ�N��w��5�_�����������D�g�����g�=�6}Lc�y.�Y4��x�}�j�4g�qhc�E��蝋!�٣fۚ�K��}� SQ���
q�l]m��K�',A�"Q��!��3�2mmJe��=��ȧ����)�2g�D���ݍ�P�E���ͦ`�i!b5�}A:\#��s5��ك�70J��Z�c�@)-좗I��X��JxV�N���V��q����9"��d7�^D��w�S�GP����ym�;p"3��D$$@?���?d���qv���}�A������j$�a?�X�Qh̛�Q�%��y-��o�p�)�s�r�8�a��v��!���j �8��d�oY���MY��.C�C��D	S(w��+��BN�Ϗ)����Q!���]N6i�<��#'���}��m}p��#K(�Tg;	��O���j$m�{�P��
�S�M��P����7%�l����Z�[�����b��}�P�nӷ{�-��z�[U�^]��(R9v{��B��R_��q�3����� c��HTA�Kڛ̕�^_���.;dkdl��o�W�D�R�j�B7+�T|���}'�	������	�?Cٓęn�=��t����6�0t���d��{_0_?|�e���v!�3Ƞ��R��ߤLi�*�S����mE��P���؟N�8�J1�!��1M�K��&'֛M� ���k����A}anz��j-ծPv眒��}�Fu�r6s�E�b3ߥ�3�ʺ�V�ÇK�5��o�>��u��J���G����Hd���Ҝb�7�񯅐�+�(ov'�>g�o���܂��嚸?�����ɸOJBAu�J��2h�Ȅ���.vah�,TB�����r��e<��o�
���<��s(2��5�'ĝ8`�nj^��3>��6���7.'��*
lD_y�-�Y��/$��Q�s3S��;��9�����p��;m=���I�(��q2��ȷu���A���F���M���Ob)f�ɭj3ɺ��^���^s�<�&����d 1w[����:�J�u5L��4�3cA��.<��~ϴwv�֦r�@�9��CU��̌8��M/1qG�|�u�`��Ƞ[uJe]����q�5!��RH����\�Q&�L���;�o����SS�څ��*k�K-{�LV�q���G��4�g���j�+@���^Y� "8W�h�����]]�^ͺbIOs,-J��Px�����ێ������R�I}D4j�ȥ�ۘ=Y�o�2�͋�ξ�j�dk�]5�8����Tՠ�N��,��=�F��@ȿz�f�=��QK��l�A�_��U$zɸ���xC* �x�T���
�,��-�wRĄΖ�� 0�Y���LP}���'�-ߪ���9P�)��95ُ�v�U��MA�����x51� Q��,����� \�c����o��Y2�A��-9�L���4&[�B�e 4�ߏ� ���5<�	�m/�(y�q񚬠K#�Ɋ���x�L�ᙥ�� ۧ�4��L�7�\�- ]�86�0���w�0
-�<�SKU�a�;�6��p�XܰI96R\:Nv����R�����>���:7��B�����qJ�'���X���Q�l%�t(7U�D�2)�ӹ�
	��/+~7�Qz?1樷m�:�]/B
�����P�/	������kC��������J�sF�1cb2#��}o ���u�Bg3���t���0ݠr��1�V¦}y����uOȈ	�9�O���#c���w�TLR֒� ]Ai�`)
Q�i����є�zBD9\)#P��������E�w�c3�;t��/XM+	l븮�&�����.B��!#�b�}�~P���h�8Ա��Z=F[�F��a<x���m,Ƚ������0A�|)�tT�*�f��98�м�$J�f��m���st���f��k��.�.��D��Z3����)��+�����_e��I��Ņ~V���q�����Td��������w�y���w��5Q��{W�g���|a��y�ˁ
ɉf�@�A�1����������"NПIQ�E�@g��u�"�{�Y�}"��"�ĽВ5��ks̮���� ��z���e��cV߂�_�	Jh�V�G��>XPNp��N�;9��&�G�b��]ܤ���2x�6���
�[���D;��hK�O�X��o7B�@�;iS�l��T��A��"�U���i�|���1�y�u�Oa����nⳬ�n�s�R��ҝ��I��T�Z7'uj�� f���am��⫄J(��/C�M*w񐥮:X%/=v�KM�@�껈�e8����h���Ֆ�}�nS�Vj�|�o�M-H���N�)�icER>B��XΟ���v.h�����3�r!Z�'A��U���}
�s��'K�d�K��&�P禵f�A����r��(�D�Y!D��Jc�g���K�d:d�,v�L�������\�a�`���w23T��xa������+,���cp�m
��Y��n�NG8�A�$���L=��.�9�.-��ZD�����xkE��~Џ�F�v�J���Ɓ�b9�Y����FJk46�*��^���+�NΧ��z [��<oI&���}2�ڴ�v׬YN+Q�MY��.g}Q��
~��	&��_�O������{2N�*,���pp�.n;I�8�']��ít�4�W�w�\�K�I(�����h�3�
�X�s3�c����%.��ѩWQw4]G�<���\߀�?_����1Η����	����GV��u����Ƚ��U}X+eīZA �~|Ηڛ�� �`kB`�6��L/�]f+�>X.ԇR������K��1��ȃG3
�o�(\�7��0=�Ճ�`|:f�r ��*�ͳ��u�5{�>��Lf���A�ؘ[���e��r�ZU��@�=��Q��g�V�pM�����.��\�#����y�H��n��݇nrD��ٖ.�!���6r3���u��g�GvL��_t=�D�H�#c7y�V��.e+�r���W{�y����C)�TX�,�9����-�C'z#n�#y�8��#Q�/e+����4�?i�|�� ��<Έ����'1����p�{14�a!�@���?�Ϋ��Տ��^�ޒ�z�#�~($&�j66��-j��h#�5�O�J�Ӥ��PBHT�*|x��l@�޳.����_&nK���P*�)@F[`iwX����4�5X�|s�� �ȳԑ9AɁ�H�Jm����Ԅ������8��? �␔=�2�^[8~p|M�/�.��Bsp�<�X�
�.��}t�CcL��q���<V���aF�~���4�j�rO��XE�Z\���Epg#k�E��>���d]�BDW}�6��m�4Ʉ�y���$����*a�l�����0���v��@*t����9�=�zV�o����BP�3ÿ-�"��`:�RL�b���Ԗ�>EmS_�b�XW�Ǳ�O��O�(��Ν2w�z����!�n��6�գ����im0p�WJJ�~=����@�����	y�q�ޏ�� �x�6�����B��w��H�ux��!T���}2�A
{O��������Fcå�^4�ؚ$x%��F�G):5}*U��� Oگ
V���i�b�4-��a��)xz[ҟ��[n��dGͥ~*oP���&�?a�Hk*�j���;Ǐ4���Å��֝~-#_�9�����N
F2K7��1�|0��P�$�����uWmM[�$8���~.��m�%�Y����Y"Hf<�� 6�H�,��ٔNUSkB�4`H�U�ѭO�[��B�Cy��%�]d���hq�]�E����7�S5����	��=��%�:ؖ@��!�B���9�	��9��!]�m�-�Cb��6*8�m�U���ؼy�K~e�ܾ��B;=Xw]�q��F������W����lګ���O���>BgGxw���֔(��9"��쎖��ul����a3Y�h�����ȣ�}�F�� �UT�ՙ��5$hrC{�?zu�X�����jm�R��T�ʛ��`2��ae�'Ő�?Ʃ�
�h:d��έ���l�j��T	8�P�
��}�{hx8�/�籭����#9��E����6?H��l�\5�B�/�[���X4�/�#z�~��N��%}��YA�ߥ�8��hMX���^}�pnH�H"�3�1(D�Ve�6����mM�(<�oO}%���1�G����O�"H�y�%�֨	UӁr!�i��{h���f��;�Gͳ
����⤳��o
����D�ܴ:�oG�Qu,�Lj��Ǖ��]���zܭ��9��>{szH���h��6�(�{�Ѱ�wsr���զJ��A���M	H��*K����x�6��*��:9-n^̶�XU+#΃�/�A:��T|94��Ŧ�$�ql?�T(!�O��MO�^�bq���m�_j�p�i]#�X�\WbqU��ĳ�5Es�K}aG���r���>�^x[�	�I���z���g����D0 �C�劣jV�M\db�ncO����~�Ʊ��z_��� �U�dn��R��)bK����Nm����&�u�����Vj�6�O��JI��DR�����_�4妌����I��Dy����.z���G	d�Ҋ�N��Penư
����deAr3�E������M��H4�͟�i�8��T@VE����7���ko����(���R�	k�ޡ�?w����E���/G,�f��b���-uF>�F=of�-`�E���)灐��@C�I��oQ7�� ��{�s�_R�#7���!�(��q��"V}�-�]�B�V[y
vY�����vT	t�� ]�J~0GD�ov\2�@�@��9l�5�1�Z-ytߚ܊gJ3H�N����������f���P�q�6��q�Q����3
h_��|$n�i�e8�������k�@TG�=�CԹ� ���(	1�Ap�U1d����~��U@���G7����/c��%dm�R6Gg^xz7�5�#l ��������S����&�$�UԌ�kI@��?��H.�氤����ϐ�r;GM�3�9�K���u#���W�4s�P�w]�a�z<�!��t��끈r0�㐭�jJ �v�?���f����v��/�Z�2d�r;g�\>���M�:����[�����K�^a�̢YkP��9.�y,\��Eaz��q/�3S�2�;��A>?���}�!�}թ	[y.v���/�����2�M���WL��\�΍s%�[b�8�r����bPJ~mXr�5zqM�>r��t��RI�ZH&��e	B�<5�����^#��Uv�Y=�8���*,r�N�f��~�-�<D�F�Nshc��9U���Cr�0K}Xa��IP��I�~�_���I��c�C�h�IՏ���}Q���f���e��-��*7>"u��#��e<��W�I�Ԗ�(�&l����������>�6�x4ű�S2��H�_�z67b����;��$h��F쵃ʘ���L��J�Ud��%^-�1�oL�N�|��Y�"Ʌg��Ű�:;���y�V�l
HрX�촞4�S,����MH���}j}jB�t%���P���	:&��˃®�9%��d�&8<5��� 7~K�>aפ�����GJ2�%|sM5���r?ۘ�:h2��^��&�����qbf�?_{#Ψ�Qsw��i��o�l�1 ���f�����L������O	�lBbT*�^,�z~�vw X��\�]֙�2/~X��&G�	�w�Q�ħ���40q9����9H�d]O��o�2|㗠����9z?�d��8����Zz0�8�h�`�PĬ�ǘcWw��鰓��";4��nۭN%�t9u;���,>~qf9h۰�M}�{�����f*�I�����T1�{�яL��6,�x���:x�=�ƍ@�ٙE@�݃�.���x=I�w4�Wׇ��t�PB=�/���T���z9�T}��Ⱦd B)c/e�^�twjvJv����L�� 9���K���:7�(�}�k!6�j��@�K4��Ճ�p���A]ȑ�hq��'�aK���3Ѿb͜���`�;dÅ��I���PYP�Whrlu	r ����u��z_O�~)��
����{\�=h�6�r�`���Z�������ck��
Ag\^�<Yd`_���@B9``vmXR�Y�r�Qp���I������#I�4��v��}0Ѕ�|�H�bH��`�;�lN,��qB�Q��$��s��ꦓ�(�]�z|R} ��Bhb�TUϑE��\��-��-��{�3�JK'���&)�'�[M�*M~,�91�<g��o�]�󭅓����ޯ�X�t�(S�A����*�'\H'#��B�1 ����M4E���8�Q��6<�,��nwd���L��2��41a���Rv�}վ��:�,�ĉ� �׼��5F�1���E�*�2]6�ɉ=�@I*�GK���2��b`̴�:��8I���:�y���Კ�լ��a狮���1P��\�#�o�M��G*O{j�g�02�j�M�^���k.,5���Z-Q�'��x�!�����gN�*���C913�L%y ��b�Z�t��ޛ�z�����������k�%��#s��t��%�	~�ow�d�>�崮j�г�;���B�Y���q]E@�Ll�4�/ܫk��U4�^��c�����M�R%^��
�}�T��a<o���\;��Xa�(8v`��F�������6���Mǝ�7�����Q��~\�X/�<�\w�ϐ<:�ٸCT��]�J'ͬ�M�b�㝞�}`�U�cR,�2de<$_L�E^ ڈֻ)����?a�S.=ȇ��d�D 
�94��!�▪��>D�2����V�����7��.�.���xI�MƂ������~���Yv�̅%oá��{X�,%�h`��b��uk�J��`��LT�q�v9b�ܷЏ\JR���G�0�&o%mD��o<��O�E0?�4�rӻ�}�)X�0M�<���� F�X�{qJ���pU����[g�C��s\�/�� Rh�Z�0i�-qk���l��W������ A�]��G�[�H�al�+�F��	Հ�A�ao��Pν��o,sMT�11���9 �}3_MX��/�6[��]UT��s�3φ_Cg6Τ��S/�Ϥ�F�J�1ѦI�vʁ��(������}�Gޚﶁ�Q�;b�һ�!H�xa�9ɛk�VqgV-�V9�g�G�* v��EX����M�a�7s�ϖI1 k���y�fĊi�%V�o�d3��ﱕ��6���I��R��_���{��n���X@��D��g2
H\5-	a�����0��[L4�٬���َ�(.�9z���P���EJ
�jB�?
PաԪ���hM��S��}�	�?�	:�Ҟ���)�H���4]T]��y��v l��.��8K)����(#�\�0�	�خ7R4w�͔�A?r��8X���g!�b�5�4#7��Y7�O�X�?��P��)Ϛ��C;NK�ѥ��_�.'	�u;ޘ�E?�[�p>����]h�5m[쒾Y���9�<�ͦLlh�^%rE
o�0UY��5Ѡ��P�<;e���m�Iʣ���m�͔z箻/��X�˜�\d���_;�C�OscYZz�]�f?��Vj
�:Is<ع�F/�]�5pj4�"�.鸤���=�*�]2�͡'�F�Tv^��x�� �پ!t-iW_b^�:��7��1���6�H�_WËW�	l������3�d�#�q�)Xا|�����n2�F<�/l�voS��6A�r����%��-���}�"�7�J�T��#�$���n�HD�6�����%�H���Jv���{�7��uT���2Y���*U�lL�)P}����G�#Y��D�����8�y�������E[��q����)��ĳZ0H6���R�I��K��Z���n�2⌷]ܻ�D�K�"��̶5�(S�xm���N�Q�i���a�W�k�H�s��#ܐ�p��ѵ�J;d���o���[f�OZK��JP��A΢i/�w�Co�2lD��߿{���!�v�
x��9K�
��C@`�����k���!��T8�4P)$�p	q� ��x��&���_f�G>�?wⓕ'�r ����Ko,@�۳��9�d���&�.�������Eي��(/V	��v����6�-�;�R�v5t��&+�H�b��
��P�bofI*��39�@�KK�r�$O'�eD&��+���[�%���At�]��JC��L�M�T���Z5.��AxDw�or5y,0?Y�=�A�.���o���-��7-�-7����v�[�"k�)�a4c�ˉf�f�� �L�)Z�j�BD	���6�������bi�MX��U8���5�H�DT�Fbc(�N,��~�g׉��v	ず~�p��v��$j���B����c|�sep�h7�0B;�d}5���`w�z�^���-���A���v7 ��˫���2��}�<2��Kĭ�N��3�z_�tJ�E�JيU#��R��.��I��md}��`��	�U;��4З���]�Q��$��y�TC�ɐF�Ǧ��ZŤ�)W�b㬲b@La�Ͷ,�'��N���"A5h�
�es�m%���^O6�Ȫ\��)&�{��411�/L��I��Zdϊ��F���t66��,�S�u�<_���܆�n����k��^���@�ݨ���U;BE�xH��������%>{�8Mj�m`;1�u����d�r ���r/�1i�5��H�_��[x;�z��u�y��8`BWn�cv`ԧ'(�v,D��1?���&�	�##���	�H��n><4��rF�D�o0����&c ���S���h��?�<k��<*	���u����|�k���$�Zqe��lba�� ȫ�k�[䯚1zOlÖ '��]ƶ�w�txQ��Pkr$ya�>�Z3�h�� �
��p�i�M�N"���6 +W�SC��~�[#���<�M�����gˎY�b�G୰yf�=7�q�mܕ�����m�c놏@�m��ij<qh�uDo�-	F
�����w�	c�35�:�l���1�-���=Q]��R���m�Z�������Ne����>3�t�8���p�n�d�<+��� x~ L�*ˉ�M, ��yU�@^ֈ��E5��7�.���*�6bu���L�}7f�*Ƈ�)��'C�ә+�.�*yR���}�D����j%8@�'��_:�(`<�C{�*?��?k�ˁ�A4[Ռ�۾��T�*k�NQ�=U���ؿbo�<srD�!�HY���8��Ib��Ȼ+ƨ��� ��q4tt��{ZK~
�64#c�$YH���
x-3��%2ңBx[˽����e�����b�c�y��* a���d����3�r�s���P#�ȼy������\�:��w��m�ᡋ��wa��յ?�Y[i�s�����.iMj��Ռ�\�[�S��8ش);Ќ��J�|�SP�\l����H����������u	�8m�\���jIۋ����@�샟S}���n}@ ��Յ�
�DM��M�:���yw�}���J���Q<�F�F�T��VX�ؓ�/����>����N���:Xt��@�o_;���s?#�ШαPYW�R�,9�d� &R#�	��6�i���Aŀo���"�B���v��R"����f�8=�Jz/������mV���Z�H
��)E�'`J.�Z��h,��t���i� 7� [n���o:,Xq��W}�P��MU'�i�I�鄀{8+|�1M��Qa=�����R���	,�7�L��U?���G,�\�>S,m�j?4�2Cm�V��x�&G/0��y�N7�#A����Q�΢�fv�)F�9�39t�M�����M� ��T[}���0ʵď�<Ca��koq�u�4�s����;�d��*�_��:C�b�.+��h�
&%@_�(~}K���^¯o�g��bM0�+�}��L��M�W��,��"� ��ev����Ԓ����_��]MCi]��딘G/�	�8/'m>�o)C7�.~+{��iRߨ����#:^�C���	~]����N�o��9��[��p�g�O���c	�g}u6�v�+����)_Q�So����ī/��(�N;o�J�6}���!G�? D�V
�|��;eE�0���>C�E�^���pcFI�a-��=���gJ]�����Q�����Ze
;��k��m�J����D-d<�G@<I�z&�fX������4���]��ݦ���w��hD����!�g�um}>&��"p����v���qd��P{��cԴW~�<{���D�\	sxz���s���l�j��0٤L(i&C);"�aO2��6�rg���$�Ϩ慂d^k$�o.Q?"I�%��MgR����p�N�����Y�V�X�F��]􂮏�����D7��=�@�+���v�@|�p����]�e��	)1A8`Q�7�^�jQk�����8����~@�F*��Č���0�n����@�m���o��Y�?��(j9Y����u+sA)�A����PdЁ"�8�tI��� ��፫�/,SF�N�Tc��AϺ��OF��C �i����R�PbB����.Q.�����,�U돺/��R�=�X�7�[�qM}[�����2n&�ϡX�	�fw���}��K�Rp����r��=�:�8F������,r
�O��b5�T�@3��S��\ d��h,���up,;8%��_�����PJӈK>Q�Z-2���iu�tb�ج96/��ිO��������%{<�2{�J�bmeT-�ppwJM͢�c�{÷s��c��D���2M��,/��)�_�e����Y�@�b<,5�e��@�#>����)ا����<�)6?L@AX�zv~�X�C��u;�w�\H��4z�گ���L2��~�P��J7��#C��\AK����N������E�@���k@�f#X��F2�8ǻ�k{�3"d|
�R�M��b!�����ȒP�ݿ��:⒬<�&��盏N,`# ����6ɀq�|n%iP� ��a��bv���>�L�NH��?r�c�ay"���,,���� ӷ|����P1��ò��=m!�R��/x[RB/�#�~�`y���a��w\g5�g]�m�R��[�˫B�U�5�J�I��d:��i�[�V�9B��$��:Th_'AW�e�E�𬭔<���,:B��`C�Qug'V�U6]A�G�P1�QOc݀�<��u�8�B�c��3�g�'��_��Q�:��Ε��W[�,�ֲ)_[�Vy�����p˕���ƛ��Tz�#-'\x�L��Ӣ���ĭj,��H�n/������ �'y@����e����Q�5#Z
��51��6���bm9��7ו�����i#��=��M��c�s ����_zD��3/��49^�g�\K���O�U4`o�G�|�1�/�8�b���cA��Z�o�+�%(m�C=(r�/�+%U�(:� �w��	{�[��~f|�D������v�j�����.��	X�OW<�E㓲Ƿ���b��-�	��1�!����m�,R?�򄄿҂��� r��f���T�	��K���3�ǥ��Qi5t��*w�����z�����ĵr Y%k�|%��\|���T��?B��������n�o,���UP؀5���lN�9!���� Ev��D%���~��֒���|�1 ��S>`s5��\a�w�d� �u�|���GC�V�m$L\��_9"�w�4��*��Xb��w0�����=�Z4�:�t�9w+�yO�J�X�:c���_;�*�c��
R�dW�K>X�3'�re��s�5�|�-���;E3�x����	�D���菸��φzh+�'�L[#�;*�X06���EMf N^�����9'Xh�D�l #���i!w���ǚ7��bn ��Sу��dX�3����5G>��2�t��A9��jm��y`��A�RB���׿"��G�`0d�R��$�B��|�n}�5�g�vt�JttK�ӝ�z?$�װ`�����tn]�x����9�J1�\��&�;9�lR��O
S`��<e&2�d?ߩ��Zk��� G"�kv��h�NnRS1"��kt��P�AC^>4��d�FX��x����@XXޛ�)����gH�R��yrj-07N��1�#b��+m�tԭ�>��L��5�P�l�� �K�8�]̍��7�ޛIG��_'�R�����&��f�+k
��a���o��6�ક~�1�ע�C�l��}@uz�0�'����~q��i}=Z��j��|�oz�Ӹ	\�7Ѭ]�'�~��$����x��+� T�Lo��9�l�_�%��{$NwV�KG�m��y��db��5�w��yH}/e����&i���S<1^Fp�����C& ]֣j�f�k�U0b��� ���4��;"�>;�Iޢ2Z��Ӣ��x�.57�� ����N�ߥ��{rɇ�$�SA�g�={P�#Q���^�jy�c �A��z/��YC,`[dOɐ�{�>��0e|��(q��="��
�����J���tm[6L7�6T6���ʺ�c��n̈C7�%TzA�I&�Cٸ�-!�n��e������G����r)�x��7����i��l:���`^>�,����}|���#C�w��JvC�����R���#�D7\�j|QQ	5�S�(�g��:d�?d߱�Q�'r�f�6�-h��L�-����3�y�X��[O���߲�=�I��'5TBz�dm@_��FA	�zBo�v�}�u���}��-�^�{�e���Ⱥ�+�������5Xm�Kk�q����n�#OJ�<s��͹�8)4�i���6&|�jG���)�0c1�_h���#�W��uI��k`�ւ�݃��h��&�v�;F��Ox�ņ�0�H��FD�6���d���qEeK��d˯J�i?���
1��w�QC�$n���_�P�m}�p�)�u�Qģ���Q�Ѧv �]Ā�����2������;� �����g�1f��p�F@3���u`�������9V�Y�v��PAU*P_���a�`pC�V%w�����j[�����؜t� naw��5sj4�]ƀ���[)=�Ba�|C�d�O܂���H͡]t��d1�X8WV�TF�5$�P0���~�gt픅A]Bh,P�p�6�+y�,�;�iz�P�Xӄ� v&WRvGݤ#r� �7�ۧ:틂-qPʋ5�|�;>��i�݈3NB�L-���}��q�ur��_Z&�WV6!�y�%=�[>mH��u�]����\�m�z��ȓ����+M�/(�&���f�1��=���1������B9n��$���be���v��r_���[	}�ۄ�1 d�޷������]5Y ��7�������C���uuu����LC��x���愆��p_g�Γ�P��z�Z$�Q�s�"2�T������[�wl��Y�-��iGKƠ��d��4�D�!���P/�s%���
`�&�<a�@�Q����tR�a���fAz4.��v��w�I�Ϋ�*�e�����Cx�~I=��Zx��t��&���q�51� i�:����	=�R��;��G��S4Q <��{�ݷ���	�Ϭ����#�/��X���Y���v��y��b�'���W��!��R!��z���x$���X-�D_WnK�{�З����j�W����Mq���:���8.�~g
붘��<d�N�h�ILsB��U��dbO�v�nh�Lӧ�cf?"n�iy�,y��ͭk{(�=M�a�Ĕ_[nG 󫄨��-��^69�~���|,X�=������z���,V �����B�]O�#T�g{4�Õ���+xg�a=6;�@<���T���As>�8���mB��i��y��3�����C��[��<](?��?�� ,>AL��p��Wp*����z��q9�ll���\���Q��j�DD��fT`���+�z�H,p�q��Fk�}�`�Dd��>x�T�Z^�2�Nv`d���t;����g|D�g�����w(����1끓/�ޝ}Rd�� Jq�r/g"����f�U����h��QH�ג��D���Wx���'�fS����xeCr�C�&��L�AzX&`Q�=e]���
�9>!R��bX�<�[�}��`���K������R̽�K"��� k��}�UM����|�����܊��zx2����N3\� ��̃O�B��@Ig]�=��Fa�o��R�TFM�r�ևv��I�/�	����/I����CJ��w�ϏN&�<'}B/w�&�&�O^��"�*B/�^<�5�s���y���>����a��%��ɒ��u��Vә�Yh-��� ������YY�ݻ��uvjn��;�!� �8�XȔ�2{O�4yV�H7P�W���
	�αC��g��I��[�'1��d�K+�͉k[�P�Q�
����L��=���U@z���#~L��Ψ����t��}�+��O)��z��_���^	��.�fNd"~䊅 ���[����R	e�.p~��X>J��L�F'�%��A8��(��� vRUq��	3qV=2!{����#D	5�a-�|�ټK�N�ts��A쳣�s�_��I6s2a�j!�s�g�ϱ��D��*]�UkF`���l��������+���Y��4�/%�E�X��i�jjv�U���͒�&%��x<�+LO��c�=VH19���z��&n��E݃�ƥ��:�cˍ���(��E�__���Gl�j-Q��v_ՙ�)	x1�F�i����EG��l�W]S��������9�rQ�Y�ӽ��_o��*2��@!���B���`��XM���Sz�1"Y��x긜~�h�������o�����+Ȏn��� �9����I΄���/>���/ǅ�fw�����v�}gj�j�ʙm� ��Fd�T3�K� ,�w��
�Y�.�x�:>���C�7��b{��^|Y)'��C'��9�.�!�.��~,�*+��T�h���)����6^">e�H)tl������U���f����WN�0buA�A��}�X�`��k�v]�'�4�j8��5SKo�<��x�<�t��_z���N��)��i�E�C2,��b��1UC���%�~�(R�2�Ķ�}�''����7,{��X�b:�*G�*tHr�q���Iy�	���|���L��cR Y�[�!8���Bڭ��� 4�񬌸y�Yy��3��4ʖ�5�N}b1�;9�F�0��4�(��Oh���l#��仰�՟B�|7�g��+��3jpӆ��Q�{�RRr �r�9�r�v\���
;+s�tYIMp�@��1o96y��ڏ��x��A >�J�M��lU&�tN�U��2�*���c<��So�i�����Y��z�m;�c�KC�V7[Yr��(������Ǿ})��"��BX1(��a�r#M��@��ń�7$u*1{�ȧ�
ck��h��S!�#��T`ʐ4��rʫ��hj<{�� J����}��b����z�Q^HEKw�����y>+<�m}�y�S�P�~@k7���X�.�Ӎ���#�����: 43%m'O��h-�\�ץ$���ե�GM�,���uO�(���0,�-�f#�3O��n<�Š���(���o.~w9�E�����o��t/��4�J2{���<4����AL�� ��Egwϗ�Մ�湛�g�����I���D�������4U�O�=�h>i�X./w�l\�U�dbܛy��"t�Bz��I��]p��� ��� ���H����vr��g4iY���z��~C���kr��<��*R4�o�7�<����&7�qg,��V(�,�w�+��sZf��Ƙ�2����!�z)� ��r��dd���c�JCu��h��Z,?�u�@�ܷsڋ=�ǔ��Gg��vc�R���X�U'x~M���Nw3J��B�����a*nH��y���T�X�G���/��wf���`�)z`�d?s��\��Ϣ>�X�'�ƒG#t���fc~��={t�@|R"*�9��s��:��O��!K�1�rE�K{,qw؜mC�o'R.�x��h��U�Y �����	��h��ن�3 2�Nm���g9v�bs�;��A�!�W-y˲U����[���|�O�U��Hn~�T���cU0���W�t_0M�|֎�d�t���!�H=��в�V��eX!\	��``=D�¦�s���zcʜg�I#h��
��G�����V +i�"?=���bE�3b${uU^?�9{w��~m�`�ۭ�(��J�=��r�ou�o�E!�Ƭl��^�'�:*�;m�SKc�nh�n�ǽ#VK�RI��pi�@�d)��nlP�g���o��ߎ���xku�%�p���F��Vhh���;9��B�q��7��.*�ٔ���b'E����8�,g�)�d�3�5���Q�j)t�����]�I�_'�aI�6z�:$ժ��p⥉<}f�0�I���U!�n>8@�����;����r֓����̍O|x����Q��Y������ii3���x�oyJ�L:�)Jp؅�T�㗕B����v-�Dm� �7V�R����=���B�(c��r��+����˔B�75�Lf��>J{�Z��U��3t���������BN�M?F��	�⦰��������$r�/7��놿;�K�Wy>�yh	)��cw^n�i^�q�1vYh�J���P\�@��.�49� ��)�j�N�X⎂N���.\�16���F����&������E:�C�2�b���y�o�����G7�ՙ��6�5E.�2�A�T#�LT�����ؑ�[�~|�/;WկI��S6�s"�l��'C)�qp������Ŋ�,dyF$�zxx(�W�k�v���:6�FT��/�ޞ�*'^�\�/�ޚ�)��'̃���#�s��D�E<;ə{��
3��m~������qI�k�L�H���Q��,ΐC��
�ۅs���|1":������O=�r�����T$If*�	m�4�qUMR���� �O`�'���	��~c�wͩ`��9;ԍ�XP�X��ur3BȊ���@8�Y��D�BQy��hL4*�����B�v[����n���/�!��m��L$E��-�;��FV.��� V�����褗��X��.Ʈ!��$l��w� loo.��Ag���$�~fi<������&��f~j�.��9u���x(GS!�nu��%M+]�jZ%�ť繀��7��p8Q^��9�� wخ<]��>Úq��94�7lTX�&�H~� 33Qh����:Y4_���ym%��v��}��R*Q����� jY�V������ _��Ja^�f���zcy�=��8�	�Ow�Vo�[S��F+�����i=�<x�0ř� ���t4�YD��/"L-�e�1Y�P&+Ze�ٯ-�`4��u֝a��_��T��6�"Ք�]�"��LR�~#R7�G����3�w.j�j_*>������J90���������(Ӳ��!Dތ��M	���{�@��:Dƽ�}Ѳ�����0w_+?��g���kˍ��(̴h�z��[����(�ۻ����;�p��n�����;vѿ'5�,N�T����gN�kȡbu��zb��ރ�Ɨ�B�v�#+?�U�>���W�#5T�i��Jmq��Hh,��Y��e㍛�~�vT���ʉy�^g|Ǉn�T��� ]9�ªɤ���A�8�s���Mca�&UN��2����G��tvj��R��x���&���.u��~j�hu(}k�����è.�Kɀ"������	N�p{�<ю9˧û��g�s�_�8�,<����O�ZWL/����i�k�	�"ܶV(O��
�Ȓ�C ��4�A���-�"c��Xj%.鐈�[��|��b���&|�Ykd�-���9C���Ki�s����~1?TU5ewP�0L����r,�<�I�t���G�9�$���ńBn��u,n��P0v8�婖�'�aZ�鸘�d�Ë%� ��sx�d�j���3�76�?P�u	�r��F�6HJg��FB���ԯ� ��YX������`	��'���X���C�s�)L��_��fG�� �FT^���d�X$�`��vb̈́W��W=]tj���7ŦD��pr0��oht�nl��'��:���7�y�!=׸Ϋ�K��y���	f���x�C�l��w���?��j����^u[���.�`ۜ����Af.��Xȧ��:?�D��8����v����*������q3�@&��m����<pi�lYO�t"��&�J}E>��kj��EI۞�Իu�O���I\�B�̔�&d��I����Y��6��.IIr����^y�~ԉA)ӛ�v���-�����gb��E��\���2^�/6�)��+�Zτ�|":N:БC��.X�4�����A|�jbx���`Y�AB��y��^'�R'⸬�Fɭ7�~�߱��1Hg�SE;I>��al֫
G���(�=��=��m6�x�#�{�����]w�|c\��q��0q.��~��Z�~� 
$T}_����hy�j|��)»Yu���FZ�t�g��Eaְ�+���͂�4~	����:�} j������il�@[$�,Gݘ�p3p��^n
r����x������o�$*��y���`RD�S��4��J�������KI���W�͕x(���Q�%�KJ�c��"|�ճ��R�cr����
0���z��1�[����
/>���jU�B�������'�Wh^� �Χa�#����5�@����^��'�,T}Ь��rj�"���1ȗf���~���ȟ����po�F �ُ`���L�ʇ��>�b|�JH�[��P`����'L�\�"�}>պ�~��3Y��B.Ajox�ol����ݹ�BJ�����7%stD���]c���\	��M��`�I*{�T���Ha`8C�;�,E�&�[�v�h�1��=#t��,��cTD7�`���Ix���f�8|����_������~#�Ng��b��Bh�Ǘ?�T�z�
�~[ïP�Vv竿�0�ٲJ�%�N���o��!z�⡆��-R��.E �w��M9�d�l��} s`�������ы��(��ǽ����*��� �����Q!
�rg�ȇI�Q�]`�@#������1���Y��6��֙�K��^l�\���:�������tv��J
�w�$� �ߋ�������+�rY2K�v�����fz�Ȋ�`���<���QA^�g�ʇ�r�?���i���>�2'�C�
	�M�v����q`����z�]H씐c��ot���]#�vV���ɘ.P����4�$���O�`J�5W��6����Sbn�]���'y��]�I��%��aP��AgE�d��{K<<��6����z~�u�a,����^�5~q��I;�#[�z˘^<UM��!�Y� ��-���o���`�Qb�M�rW��qג�$���� !�l���v�Lm�F���v=Z�p0��3/�������vĢHBi(�p����q�{�S� ��>�i���
/h
��)�1��'@��Z�T��>�x��ȗX��Tf���J� ���A0��j�V���e�M�G�	[H�k�Om����'���Zvy��2[��HXB�0�/^B��wjh!8��s�
}f��W�a3��](T� ��r����Q���)���M��d���Ia��dȆ'̼�7���5	�;-�����;ߍ'mc��6�wi�6ԉ4n6��F�`��"ܮmr�D�{��,�7>������=�f��w��O��O�d1.��00YYb �5�������Y�ͱn>(Fv� ����[�à`�#�P������՛d+�&��>�� ����~�c��"qod���2f�t���#�C6����x ��,j����Z�y�a#sZT+m��`���Q
�v�������x���Yt+ZXH�9O���cN �RDla��!��tgQ�ϟ�^G�@+�׸y�����>�bHF��X0�x~������ۓi�`��bvhE� ]R��6�E>�)'.�o����p��;nz��á�u>]#�S�r�j���wR;��[�w���_������[yY��h1M3.�c(������ /�d��F�*U�KֲY<G�_̻�)��1l�#֐9�>f�m�	"f�x�[���a�h���s�;�+פ.�EO8o|�7s����צ��F��
�k3�����1�m�XUP,���&�
����Qf�b�4��e��Q#�Aͯy�+����0`�:�a�dmNA(	���Y�D��ڲ�1���e�)��@xg �򒖜�߽xV�>���̯+�B+�""�w�ns��3l��I+W�iC�d*��p^�j0��G��bC���'<�_B��3��x3�A�܍�"��p��,ѹ����M��yv�	$u������d�-�{R�$D��`\��q���Ӏ�`n�����/^Ju�c^�%gG��d�7�`� q�勏�s(�ek=�������~e��&q�=u�E�X�d��r�����}�w�Z����*��*R��<�i�
�yL	v̯h��7<�E�U�W��C&�X��a	����;L�����x�+H�{o��Ў��� |�� �n�co	s���]v���1&Yo����l�X6b��qۘ(�v�$턾�"�3��j�c%����!礿�.���N�W�v%� ���&�_z�� J X���`Q� m^O���Hb�˘1v��~\�v"+�5f7�S�no��ؔ4��)�
`��IED䬒-�J}b�<�#ݖ�\o�m7YO�$X�&�fȽI�A��j�N;���{��|w�W�"ت�K�+�쟕�G��71��{�0���|�8�~����Q˯A%PJ��da�[���.�ϥa8@z�~�+�R�~R���;R;�U��ٵ�Z�G�l�Y�0Z�pvdka�	/<߹���	s� KJ�l�V���O�m(B$O�zS
C���y�;����M���)>�`0I�SK�#��e���I��f�z����07h��"����X�M�&���8����0AZ�Xq�u@�+H��Tc�Gd{�O�����o��_����~��|�b�B���|��c��"n&�)��4n��#�6���?=���Rq/�Ù4��|���'�-���ʛ�n0���C�dU�2W�y޴��diq�O�f�I�kfZ��� �ݝ��m��aW��H�'f���3�`���5�	R��.j\T������cU�d�"�<l�����l~�`���
���q��S��(ʸ"��s�D)�?՘y��R�׈������O�x��k-�!1����Bu�J����w���ak(��7�g�L�=�pc+?{o��{���g�)t~�\�M]dTy�@Zex� �[��3('`P�=]0	�LM�M���~�Ϡرi��&V�s�Yҫ�Ѥ�Κ��B+,Fv��P��������%�� �q?�Yy�����d{�H3�9Θ��}�*t�rD��;`t��U�<�ӿ���9�g ��pB�a�*RRƏx��e��TF;�
����W���*˓�LV�<���;�O���1�?&�Ώ�ѐ���YM�C�w��A��B�JW�f��K��<���3�w��}D�E)ȒϤLyT8�*59i8�g��AT,���a��W���n6����FN���O(�A�O����o	��h/�=�o�FBk����k�`s��֤3��y��ʿ�8/�m�f+�.��_��X��S8A�zz�;�bdx�_X��_��y��8��H_�����<М"J^`�Rf���:�Y��x�O��u&;>�t��!��Ag��#�ށ6gq�@��+!�����.�1�K�ӳ����>��� �V8�����|Lr%BvY��$$י�;|<��5�?�����o�Cdm���<�30P�5l��؂��Y�'ը<G���,ކN_���~Jٸ��͐X�)���!�%#� �� ��̟AU-�M�� �B�,-�� �R3	�p�^"�W����Ϻ��#�N+�9��� �؄��.lC$iT�V��H���q�@�~j�s�_>�@�!�Q��8;77}�Q� ׉L��k&�����@mN�77���Băr��I��^e#�Q�|�
f����_��Zmpa����Sp���Z.x�������0S,ZP�.�]Lz�[��kGʐ�����{����t[�d��Ar$݉���u���j���ȗ��45�p�,����
+���;�,F&�	��|S�3�G��ҹ1�g���Cl�z�v��Q�8�8� �z�^�����w���a`$ p=_�C�^��.�r����2�3���]#'�2�&�v��a�2�������>S'��7[(�<�ಓ��F�2�fz@��+��~6\ဗ?���@Z@���E�>�� �}
}����h�!�T)�G#�g_����K74��/3�z2���3(l�B/o�m�o�w��"�%��f�&\�أtI��'��AF�'[U��Y5)(TR~�}�*����G8�B@^��f7�����ǬE����:N�6G��v��T���6�i��>)�N�Yg�D���.��x���W�s�Ծb}W��m�/���x`޷��X�O�g�hﹼ���ze�y�ڞ���O!�ڵ�-��W��BTQ��!s��u�!g�Ig���x�R�r�%����ǁc6���ߕ�x�M����8�̥`�A r��oV_��x�B��1EϺJSSA9o^�V5�w�ūd���ظEU}|uѴ�%�Zufu�n�8@�w�cN���g�ҕ�7w��sv��U�����o�A!>�;v��f�wM��7�;Q��
��K�(�ĵ;�DR��Qݴ�6�)�1���~�嶭��jp�6n�������`��T/�#t�q�0�iLE��K;)�6Jl�-�@���tPA�V͹&��A���g��������L�-?�_S�[�4pEN/�$�����~hZ�z&�QG� <$�x�0d���8�n1�_e\�!��Jn���</���sC�Z�1 KL� ��T�G�5�bL$�Z�e���8�߳�kc�ƋZ��>��o[�S~�|��O��ziX��&����}7h�Aw���[G��T/��8P>(,`l�RF�IC���4�٭wC��l9!�d�~�y<+�O��3&�O0VU:\>[MO޷J�o���Լ�|U��}��p�dbyCIT��U�A)��7��a� }*nL��.g/Q"�~(*��N�>H3{����Ṵ-߾�����@|�]�R.j���j��K���A�f������~�5_�4x���hR�8̺Lx�"4 �[�E����H�翓VS|�.4,lȻ��-�ʦ=���7��h�=���Co���?y�4�_Z��vɏ?]�Z5WϒE�T��xd.޶�7HR&4j;�4n+�Ǟ3�?-�n����~��0S�;�<��[�Z&@о�0���4r�ѹ*9ʖR�L���P����˴���/�(\��(�@=�����p��1�9�~|q�.�8���w,,Q�\�Y��?�rv�-
|��j��Ȏ��f�����#�\�=F\�ߛ�'�9���ȃ�c�Ғ@q�ڎh��"C��u��j�-�"����Xs��(��l�v^��x^%n��Y'���Og��U��mw�ޜi�v$��C!闇Ĭ*��3 ,����%l��vR6tH' U�'��Aj-�`X���vQnE�E�b��F�/>��5V�G�%������(�%�~�j�A#1]T�(	
��B�u��X��xk"��=�{�-#NŲ���ckY0d=\��O�O�[b[��ml�$WjA�4X;��mi4���!Z`l9��Đ���-ߩ�ɣ��*��� y{��X���ׯS�Z3Ҝ���P�`	&z-ݼ�ڟ=䩏 9��Vu��v[�?d��ז y�ӏ:����L����������(x��)�`�6q�Ix� ǧ�Ĕ-q�ߌv��@3�Gn�.���~�`E1�Z�Ljmx�G��5�9�n����K]��u��q�vH��m�q����.�r?�����c��0�}]v�pW�6�N�j���	gT���(��tO��{>,;�HC$g��3	_�����	���f�����+S�'Xp��/��S��2&0�>Q�s$EP��'�ʄ�H�����~E�G�_��ِo�Xb�����hV��F�eMqD����S�~|EC���5��������n�t<�҉t6uZ�9��;z�x�iI�*{���
`q�<	$Tޛ=��d?#���IZ|��k�i�i盵�.�<�Rܬ+�>Ϸ]��gĞא��M6:|�φq�L�~ǯ"���
OUb+5/��23���uoP�˕f]#0Ǿ���4��ȬL��u�1
t�SY���X����B�Qi�z�A��E|�N��
78�x��\���ޟ�t��2L�5�sW}�?�+�J��=����������B,�H����$�7H -�ͦW���!�=���xL�x�0��ۯ]O�c������-����:���q�a\�e��&����S���࡟U�4�/n�/�ZM��- �Hv�k0�_��7���)q��|3�ıF�[���y�]Lg�CV�WٝH�0ɡٙts����_g���O�(�)G\j��������U��{���~�ǀ��hV*/�z�#�]��\�޾a���X1&�y�@@����`K��3�Dҕ3��1�����	K%��
�i<>/Q�%�s���H'�(LV�+�p��5Kr��(ܑ0��l���� �e��jC�iA-*�0@|,^y4W]%GU�r��dȟ6��a�{����D�.MSHu�A��o_��>���Ȁrxu/�/��pͧ�5A�F�J�OF/��ہc1�uN��W"gH;C�@Ka}#�Vz����.�G_搆A(YM�B��X�77����PěXt6�@����)�`�-��U�Vmˉs�� �L9o�SO�'E�l�g�P7�B�6;�pymG3��R��KP��R�_��������焆:���rk��H�;أd��N3�;AJ�h0����Uц#P���*(�|�4�ԫ(N��z�C��l(���b�u�t	��d7��2�i!'�YE<��-���$�4�n��ç���!�0�3U�������lH�pJ/&d�@����5XX�'ԕ�~w��B�x(~��Cj��x�%Mz���.���R'��@9�G�1ULX���y-±�&�=%Ӥ�!Z��d�A�0�64I��!ċŅ��%YPs�@��9����Oa��'���>hظ�]�k�������M�ߍdp�ۧo�2o��$�"��~t�����.����U/��0�3����1�2�}�L�ʪK�R]�غ��1��N1������Vq�Sr{�}a^��x�`�<��4$F�tً��52�p�*�Qg�G{;�9w��ٗ�]��!V�yBP��������ʮ*Rg�b���,xj�-\�F����iG�3r�6�-��e�j`�v�u��pTAerClI.�B�k�0 �]c�b��.U�Oج��V��[��c�[V�"ע��Y�+(���
�[
���v�Q�^�t�%���_�̊N�B�,_�5���78�� ���0���K�٤�薙5��ͺ��P]_H:�,�X?��9J ���[ze��!��������X�{8�����	��΀O# �̶�G$faU��Dg�@��	+���3�ɟ�o���<�k:+М4bҴ�
��G/G�5E���?ƨ2�Ǖվl�F�Ѽ��)�'��C��[�ǋܠʂ�)�1<O�Y5~�(�e�$HÍ��!�h���_�����udʭBm_t�xWg��ϟDv�J��c]�zО�"�| F��:���d���~�D�2O�E��0���P�?��+�t(6�G���ߴ�ޢ'ߕ���+k|B7��\z�� 9��K�-���ҲM��ׁ`�`�~�q��m��y��9Z�؅�
�,�hU�3�nj�9���������W�+��%��0%x�*�ݍ�F�_��@�0�gأx:�E���P#P��l�����s�ge�����D����c��,��;K���'�' F#=�$�S��{	 �A�Uxr�����ݧ����W�6Q��AS��N�_|��/u����[}a6p�r��o����9<Ѽ���,�w�a�\6!>\X�,��Z��R�=~ܹC�*��`@h ����+�>��t�>R����T7���7��#Eh������~��k!�	��J��ă�ew01���K/����3��a��f�m�{�
)N���x�6���ݻ�0D��
����jT��Rz ��z^ʡ�,1����HӂE�ʹWe�bh�A�T�Nü�0f�BX�8��ÿ&(��R��I��щ�7�/��A=� 4�"1ǐ0�U�I w�n���lP��:����4y�}*.���6�ՆCӀ:�7ڗZ�T�������$ؗ ����㬰�|����>�'��"���F%�x����g�;W��H�=�P&%Q������*�
��s�ah����p�Fo�5���6�'c�5�st�	x���t��D�U5ȺЇ���<Tl��
��l��m� ��R���&5��-��'�3��j�(��}Rw�Ab!m����P�6R��"f����#��������������LQC�h�l��&P5R�U����P@/�[��F�Z��/��������~�d�KpʋW�{rr$1`B�x���ىKs�����p1�Kg3����I�~�r�� ���r>=���.fea�h������b�]��`��I�B<u$�#��˽"}m�!��ť0�1����E�I��U#��b�-v��E�# K4�ً�P���%bJ������W� $Z"�1�����\f��v�z��h[����H��V��E����P�Y��I!��<^��+)d÷�C}��Wo�A�~܄���g+�<j�h�o,Y������d�@0;�}�����{&����/����N�����q��Yo����]KG[�3
q;NOY�k�Dq���Z����ۏ%6V�xz3Y�=q� `�cmK�O3���~B�v�Q�ƕ���k�n���2�Nc "2����<���y���5c�m�6�H�9X`R	�QB�����Ka���mZ%%�<:�q��J,�W�%� 2>�F�tГb�\N�k-�9�@@Ţ�!�j5���m�O�������,l�}e��n�u��UQ�k�ď��A*�t��>�A�"��t�$���*] E���ά0]�%!k��ů#�Ж^��4��r���}Y�/�T�LC�dے-����C����x}�2{���q�ux+�f�{Ìm>��B��)�J�9�;\�p�q̕"O�H�b��t@$}�o����9���I�}�[���T1�\ˊ��
6 �w�������y%f$��_08��Z�(�W�}�q]�3�b���K�:��]�.g�O�OB��i����n'�Z]��S�!��+)W��� �0�V��%�`Pz`X���o%�a����X�z�2�e.b��a$�<[�o]鄫8�uh�.���M�6��q������F�Q@����ҙ�]>���A��m���D�?���,Ϛ�܃S��{-�{BS]�((co�#�sxÀ��:Փj�1T$c�fc�];J�Z�%�/��C�	�/R��vX��ֿ�U�T��}-�'�,9}�ye?*�V�f���c<h@ą�O��@�d��x4���aD�����?��`�|������`��JPnH���1��q�zFׇ�d���oux����4!4W0D>�5�"Z=)�ñPXt�b�,��8c}ߴ�6��z�����V�'��4��"���L��r�ɟ��FM�b�>e�U%����a����G����(�^�j
�3z�� ��6�d?�0��tO�� �/��Э�Y�3H{�"�»���3c�!�9�9��u���*�Z�'L�A5��͠27"p��I�FG*Y�y��I>�R{�و�cKC'���F&#�����SE�3|5��R�F���|%V1	V�+y�����SL��r�o	u>����50����N�7>�Y'u ���Z���d���;��X:nM�\�}��G�r��UkP�@��ueL):?|�J+�L�W�]k�jN��xf�|����G֥|q�B�j����kú�g��T�@��y;F�g;Ph�״q֗�eV �Ռ�iJ�kj@{H�K��'pw�ɡN{��w1�b�$�]=G���<9���n�e�|��L��Z�G��e��ܶU�Ɂ�����P�!^_xR�RD=3P�r���F�/70�Y�T�5`��1:D* `a���ю�� �p����~K�g��P�р	{�=t0^���!��A��^�Jt-߹�iF�9���|}�M|y�f����=�Թ5�Ԏ��rB�%'��Γ+y�����-�,�E%\��//���ح�r���r��#Z79_�r���#�ov�����_��\5is[��$���Um�I&#��l@/?�W��K_��E�������b���;���M�"Y�:s�vT6��z����^S���f'Mњے��E�������y�+q
;�L���y�|0��٧�3�܄H���@�ȡ�1���l��V�"I�pO� �������E�fX��IFFc`�::�Z��Q����I�}ۊ�:k��t0d�~ъ�݃r��,��i�Aާ�������!���3 ��[)���izZ�d�*�76�V˚����~u�I&gY��.(pѲ fOY��
��,�-s���Ӡ2;�NT��)��=&{�<
�Z�4͎��d���f�����`��{�˕z�j�U���d-��#��-�ڗ)-��"���Ƚb>[�|��l�'��1e�jԖ����xA׫�b�~�����}=�:�����\���W���e�{ �>r�y}����y�g�cj�o�@��;�L���/���{'�N �q{c��C˛�f������@o�r���B�s;�����i��j�z�5���U�u�Nu�½v'����g�H-f����(c������iT��b��Y�[E��v"��[���^斏h!RI*�a�q+GN��*E��/i����0^�����!�@)���!�x���ϳT��0�ZvOLW�I�þ�t��{�-�Q1N ����к]�7���u�}[�o�פG�B���4�:�jDL<��$�䣛��|�R4A<؝��}�$�ز@�umf�Զ�H�u{����=�'�{�>�+zz_ⓘ�@�À��L���D���:��'�v�ȋ!���}ҋ���u�K�A���1Dȯ�����}�벸	4���g]3W�R�g��
t�@��m;�jܹݥw�I��q��B�5K����f3���s4n����iUѣ��p� A��@��ZHܵ9��@��#���Sj����=c�KwM�-V�}����D(f0�{�%�1��42MrK���a\����H��\O}ZQ[��i��,�����C$�W=6Qs�I�ĺ �F�qX�4�L���ha"k��/Pm��o�D~2�~�2n��C�t�b�u�.xP�Ŕ����Y+�]�}�f<U�f�)bM�%ݾ��Ip��}ia����b�4��D�A�������Y��t��|uT�M���+�pR��9Z'�/|��"8YH���^~��U�&MS��kxF''����v��b6o��䟮�8XQ��y�$ŎHmϬO�bH<<��ր�i˟��op��+�	�+�A��z]H��3Rz-��/����*׊��/��8C�Կ��}�*@�#����	K=r�3�+t����������t�9R��f���=�qA��1�9́��0�6~}�����{�����j[ى��ɥ�]��:J9+ӈ����A%��ۮ�'�EF��!$�����q<�eu����)j<�!x���Ñ������[?`[��̷�c`}�9J�P_����}�g��0�+<��o�-Ԡ��U�uzUBP����vy�:��%�a/�� �L4�DK��,��|����0=����^��r���>0�A�gjx�.e8
�9�{�b�8\j����Yo�B|�E)@��u��U�TV����P��ж��5�
0R�[�w�)��au��ەu�倆ҙ3� n��OC��m//��u�-*���jxs3���(����ч��d}E�6E�l�����KH$�rq���A9�Q!ᙷ���v�N�2{ۮ���˸��n���5q�D⾉G������`�&&��@�OcO��J�S�ǂ?Q�˙�+iP8��j�4��4��/�.�5	�������Q��n����&��cs��Z�a Sh��"z�))K��}:�z|���=Wx�7��M-'�[�x�5��k��K\���{!{���7�v�ʦd�2h�K�t�5"#�����>��IqB{�� j�����W`��!�2\��1�w��#����:=7H���B%�itx]�����uRSRٿo�|If��Wg��^�ޡ�0,�'�����|ʨf�EDn@(���k*D{WB4,�-L{2�~��Sڿ�S��!Lv,��j$)�Da�D!i�����J����D@�+M��2��U��[��h��9�]FL�߿���>�j�#- 5�~<rH}-{p(Y-s��5�؁6�ә�,`�5�m�kS�u���$�c<؏���� 46gm��+�X��K�޵�A7����B�C�����؅����b��*�#9�g��at4H}!JDJ���ʾ���mjh�ʓ��
��:�{����kF���j������G7=Ռh$ҕ������N�T='���1� ��Ç��D�3�%�54	��
��N���'G ��"0���Q�a7�ܡ*����`�r~�ܤ�$�Oϥh�
��4��eb�q��c_�ȓ�1�*U�؞�+AE+������� �j|�3i��>�����V}|V��J�]P5��"����z	�8(f�_4ԉPj�k�����m�,���p�g�>&	��}�Y����w&gU~�읂B\U�*�+�|��5o��6�^���R[lxPC��N���G#Ve ��͉Iov��ӿ4%74i����˅���f ���p yd_��J�P]"��Ft6�'�1A��jaܑ,R��v+��>:?wY ��N:@�W�̍!��f�8�.����6NeH�bP5�*[r@�dO\Q<�#��SI;��-���5�ͮN>/�D�H��\���Ʀ����r�J��L ��}7\�?������[�mC�{,��� ֗c��&�<̄H9�E�&��gC��T��H�[��m*/�ʖ��ޏ(J&��������Bٓ�VG5�
8\{�\j8{�t6���t���n��&8%����D�B�t����͍l��IY(��*�M�ME׏hu��|�S�a�w�C��z��#s��.��ݑ��1S�Lav+��
�㷀��o;c��Ϟc��ڄ�l� �����i=tm��c
q�W�I��$�����H~���EIl9�q��x�hG̖:�bl�ֿt��>����^8@�!�b�/%��2j�?3�s���k)�~�h�6��]S<�j�_^�g_T����KE��J�n��}���`s�]+Vy1ʘ��~G���n���jc�u�3�R���<�Ĭ?��V]�NYOJ�Dn}�N��3Yv*]��̮��+`2&�F R�����r#�`�^mp�hӺ������p��.>�~�bf�J<�3�TYO!����OlϜW���){��&��re/�m�z��1�x���YˀgG]e�@=A���ܯ������u�b�����KZ�:5_�D��x;��,�����r=�4�A6!��T���-��9�s�[R ���6�}��ub1��B��|D�Nܟ ��X:<��6����c�d�(R�K�K*�P�B �a��W�C��R����[Y:��CB�e�EԚ���bc�r��`�Ī�n���"�i�zcՅ�����#5YQJ��_Mh���t,$X!�L����o"�8@<|�]C�T�'B�>4�u�~��`��kN�H��L �Q������QU��mtU�m׌O]�^�+3��N���S�=A���p�v�?s��V@���`-F�%�.Sѻ�m���
<�ʒCh���<��n+�d�!�2ڄ=xHk6��x8V��kg��hv5���M��3H�uNĲVrl��6H*U��L
�5uEqWN6>��Sa��7Қ�������{k^[��D��d�ʈ��qA�����<��֘��\yw,��&|��q�Q	��W����]h��tЫ�)h��V7�j���ܚ*���������?�^��S��zG����W�
�$��-���S�#�����\����T�0f�ͣB�N��§�����s0~z��{qK���D�N�@𙈔������s�[X��g��Y���j;�dl�,��7]�l�QH5�y�|dxO�S��/�
C���>E�����@Vf*&1 %����Aő�.��m�l�J��NR��T�K}ޡ�������]�������8¨ї�~�{0���=0.�a�;S��_�.!��!����y��ít5!�c�(�� #����7��o�J�kR��,dn� n^�T]��OvEIܠn�����ɵ;��H�g���+F.P���������k+��<l|�4�4l�r��q����Qs'���`=��9��rD��@����� .\,Bm8���r�1ߓ�9�V�`D1���9ה�����S����Ζ��@b����ݫ�����K�*��*�{j��y��8D.�NS�bȼ��yB�o���)���k�InP �-:��(�(-��Yd�m4���%p!bs��J��:ᬛ��ag��Y���׍r���@Q�@7�� ��iP�cr�%Vϑ�t�b��D2U�u�Ou�X;Hܷ_X��W��Qk�1�u���1���QjD2��3/x𜴨! Xz��O�@˴�C6����Ƈ��'�t̉�O?ce�jg�1 J�hFⰝt/:IwF����n[}3u��� :H���}
���	��۪�vſ�Q�N���(w'�����N�ef�r��d�bZO,��C�;[r@���������Ro������?bԋ�������}��u}}��8άCF���d�R�4��~��������Dr���̆�p��i������6n�5�z� \J+�#��Yj�	c�+����CJ�����W�rPY�\��ܑ����b�k�)iљ��j&1@��u�9�&#��H� =K�t����4�Awz~#T������q%af�AQ�\��%���Ů�(�fzY5���@��y�:{/_ <u�,�� ;��ZTBg�OD�����|�Vv�F�����hߵK�j��R+�^T]T@T��i6Sp� l��j��ꜭ�U{ =A��	,b��f)��&���,ɐ£��AύZ��ya���ٹ���x�V4�e �<�e�D�v�qt,\�]4��Y��S�s�^���&���Qb<���-5��,ZX�C��.�i0�J�9[��0�*�[3\�9�%/�h�MA���9�3jC�����@&�p.LtPl�hx�sdp}��Fx��_�\n�C5\5�~=N�L����i
\<�>��a��!��0�맟�-z�qa1��7�rġ�N�1�g�E�d��W�rb��_�6�X�أ��C��9v7�)��"�u��~�go4��BJL`���Μ�mW8��+�.@7�F��O 5�P�26F�A����\i��8nD����k��~-�N�êM��T@�QG�m��J&�@ã+n�;+�8m��B*��"�K�9�^hc�}8ЈF��i������vF���p��0�4i�S�(��8*�ǎ��\]SI��|�J��C�}qp��{�W�*�R�����5j"�^��o��Y���h���4ipMHot��t]m�H�p�Hk�N��m[��ܗ���I�����v١`���6,W(�*I�C��Y��
V�1ϼ�l�QB����C�"
�EݔW�E>��+#gi�&��[gJ������1,+b`D����z�p�l��� ='������{�о��	6+�X[�/��b`�-�`m�H	���xFζ �#m�$DW�<��bF5O��~?�w�J-���KYa-w�<�١��Pԡ�e{t_��+��/>U���4��>��W�MFxYlC�����D�+#K�pV0�1�Zg1��-��RI~�kL��٥���Lc���|1.�a>�>��v�_�n쥼�r�r��*B@nƴ�RX}�Ѯm��.#��Eo������p��I�R5��_�K���JЇx�	���m~ЬS�ƀ4���!�:��]���6;w�݇�(~ZYR����{���=�*SԵ,����2rV�^�㢌��!!�q�+���5d#���iPk�q�us�]���j�`+Ht��hp��XPe��1��3���W�n�C?��zm���[Q+��p܂��`��'�ֻu�� ���ͤy����"@���h{�<�	�]�+#��흗�fZ�cAڡ-WG�_+�ڤyاl� WI	�=��,CmXb{'���XT�du���D�U���6]U'E�Ӆ�����-�3��j%3k��F]��J�����Iu��X�m�}KL�;2%�q
,� |yz�Ӌ#4�8{�O��E4�v��M9ŜK\�O��(?,�*(x7޸���q5�����l�a�S�=���/��o�oE.+g�����0��7:ٯ��s�r�<��t#��Ը|郄��Z�+�L̻iA�o ���Y��2P��Cτ�w ɴ��j��.K�ˆ`�\!�V�<��wX�E+��AHc�����&��!t����y�>Bn\3T�Sm,0P�
Ihr�C�d�L$�
�Oh�Dh�(n�Y9|n����B�-[�9���6Tg)HCP���,W˧���0�
�i����#��w�/dw#x��>ʞ[���c���Y�~ FnU�}��\s��2������ E��؝����Mt]�Q�M��cI��-"���gD�����z��~y�#��Đ�:�k�o鷤^����E��5r�*h�'ҟ�p�����ec���0v�}@�Y��s�u���������9����q�����[�G��I4�'&,�<
��Q��,㳘�J/��=�V"��R���X��|tt�#����e؛�֒\�vh��pW��9�o?����1��NӴ��|��Խ't���q�h:�R�<�΋$�$U��	��$�����d�����r��(+�$N�|��vre�2�[62g�1�_?従��ɘ^E��:�2 �*���̟��2�l�?��hP<)�����o,�§PM�E���X��m�S�{}&�,v5	�1ہ|.i�%rѰ%I3�!���.��_�Q4�������Ѣ� �j�j�	7[=@�7s���};g�'i��ƭ���`�����36�k���÷f)���Ӈ���}aI��-��]��Q�YZ���`�ᢢ�kR�Ҿ1ֽ�)���_�g8c�ǘ�|2�������{H�l«.7�@C,���%y^�(� ]Ctќd�
e�9��K�G��F��bYz���	����g���3�dg�k�+IdU�H��5%��
����| KN!S�9���MJ�j=����F�Cp~�"0�6<���OA���ɴ^�����k�r�J�S���f#�{��P�����<��H�7>[<��(d�1��h�Ȫ���U������,zd)0Ģ+ ������ �ݧѹ�W>ML���p�m��K�D�)w��6�K)Tk��;h_8]u��U��
���?  �[���9�&�C�2O;p֮x��r��*�h1Ĺ�F�h�civ�F
�����ާT�S���-�9�>7,C|H]����Cs��Ǜ�G��&6�7,�� �e!e�����f\��-B�BA��Y��X`j��O>]��1�Jny���� FQ?�x�����1�V�(���ٻ��AHr�v�ܩ�d�1<�W�MJT!Vn�_���j�Q�i�v�Q�ok�}���8KPJY��rE��@�w��>�C��ivߎ�;�!q��z�T�	7:BKOS��U�INJ�&�ծ8��5\��^�WxG=R�P�fr:/ �Ȯ*��q�砍8�H�+���6��W�>�!|s�qk�L�&;H�}�*�mf�a�����Ci�a��]�ދ�VF�3�5i1ō�>�4�_A>l��+�G�.aVk��{��؟g�S�z�~���#su�>���x�����=�P��e����� ?j�I�*"�U�2�-���Ꜹ2z�W�Tg�U�k16�w��T�Q�CtVӭҥ:�&��D�ՙ���V���=�))��8g}���zI���~ڿ��5`����'�0�t��� �L��{��b��@��gLl��)�9�{$�������1OD���x���_���.��<~4ڷB�q[�WV�q�R9�$�<�C�K��_�϶�r4�a"¾A�d_���2N÷�����V���CM���ïS�d��x]��'ڥ@տ ��mL�Y�b7n�ڊ�Δ��3ϥ���f�a����A��
�Y�0���@�SW��V��G�%$������3�s!L9�%a�u�t0D>��h��X�_�5�#^�D�����d'9�]��J9��(��v5t�@hv���7:�1'}j�O�&�7���}�Lϸ=��:@ż�%�F�R�)�AJV>󦝧2¯bg ����v )��q)�lU����5ԝ�,��=[����_h'o��q��6��3W'�w}�#��}_Q���������"�X ���%��?�r켊�0���̼z�X�7oòM�u�����R0�ݣ2��,����Ǥ�X�A� ����-���BﲃZYRD��6�V\��u�pJ�y�L=X�	�&�w�]%-T h����41tc��n����|����������kJ����a��S$��DQ>��m�c�����1ٷޕ��a�x��bׂ(�D2sB�ы:&���0f�Q�Y񵞠�P�U�^f�:#J
3�犆����A
��r$�������5���T�
8Z�ψ���ܖ�e1���|0]X�����T��|�u�1b��@s����ě����R��[��&̑c��E����Pʶ��=mq�K���ֹ��[�Kvfկ5s7���B`f3'��*�|��]�.a����^�a��!�K�S*�rw�rgm�_��RTf�g5Y�t_7Q��'3Ci;��O�<�$� � )�P�gY�Ư�� j% %����>
��n��<�� X졤�W���;q�5b�W����ｊ�4�&$�Ҫڌ�=oТ����qx4��YBN>��}')~�F�[7�paO�A���*q�(��k��Λm �0\|��"�:Z});��x�kMzoa����o���R���H*i3..��+��㷶&���K%o�q�{�`�	O� =2���Fx͕�/���H�]P�⌆�߈�`PD:n�����߷&���8��Zufڻ
F�J2آ5<�8��X #I��;��<�t�t���F�R��kB�p��n�+Yi�Z��;e�I��"K@�|Va�8��1�A��ʙG��
�5����W%�ͅ��:JPˋ|���]V>���õ�4> ��Q[H���!dP�.��LE�yF�kp6�H�!L�tP��]8f�m�����~��"=�n7�wa�b�N���y7J.�� 3j��-�m��Ü��4���Q���A4�<�s�G�sj��z����3'�k\!Tn#����V	gܧ[��W�)���E�%?Q�c�c)����ʨdC4VC��m�G���G� � �E͞���z�ש�I|ec��-��/L�x�G��xh�8i�SU�=a�?m/���m�������@�sӑ���Qj\�,S�����S�7m^d��4.�,+E��e$�C��*�!_5?��;�Zod���2Lm���u@�$���3�!��Ó%�(�I�?�.~�<-�[@�|�����}��f�U9�޲k���O-
��6�.��-ۑ�`��*g
!�c�ߦ(���BK+�����]J�ի@g�k>eaK�u��CWGu��q���� ���̔�c�񐘍�,Ԛ}o*)~�+ă�W(b�؃X�y��
_��aR�a���킣ۻ�h���L�i�����O�D�mWU�j����_蓤9%&�(i�=kc�L��2ȧ(��y1�	nZ�wg0�]`�fť��bh#�cބ!_ܸ�
�&A��Z�h�J�� '�^����m������Ԟ�*�p��e�#P��v1��[	VIڥ��s5�
��ct
�j8ҲP���V`��.G�/e��B1�" �`lRS��" ����+�4�+���0�<����m8�N��m`Ĉ���u�kh�ę~>%4rgzò�^�{C<=�m���K�/`XQ�4�\��@vme��	V\�V�3`o��څ��z�t�	��*!��U�m�g��5龸	\���od-��x�:���^�h��i�Ld;1}Ke@t����l�'��G}Tc�t	,���Nz�O�d�2W�Lj�X*�	��̚]�uAVmNg3�ID�Y���ͻ�� @�˔G_��E� �ҩ���ݷ��f������N!7<kUW���99����� �:�;�i���u����`0���[{n͆*dd�f����=��D#Vw0S91�Q *��<\c���<K�+r`�6����A�%&;V2T~&Mhb�L)���/����o4��y�|!4�
����2(�cHʦ����v���=)��kɀ-5��G!!��o��y�_�Fqrz����3DYg 0��O�@{��R��	o��?��~�#'�%�y��#�տH�'?��<�9��&=% l��@7f�;�g%����7������_]S�����C�G5��5��a�q��c���DE�"�G@2��O�����mLX�/�ߌ��w��2�c�LK�=K�{�0l-�j�~�;"WQ��_�&кisg��_�bX&Ud�(
�tt��sֶTE7����������b
0-P��5�{G��1��ǂd��!�n � ���ϓd��M����P
�k��D�}|���d+��読�V�v��Zfaۋ�C�.�[�DA=�����(��Y��2<(�����¸I�R�}P')��H�Ѝ�}��`Cm]�v����^�6�B�¤�m�Q`<G��"��7���.MXR7�8*@��O3�ZǓQ{	e66o��H���Muھb��S�n�Ⱦ�m���+�#�E
��1+;z�wNͤ���I^�@�пs��?8Q��T�4���}�@�?����QS��4�����s��#Q�T4G{RgXnH�~�=j���sM��s��� hFڠh 0\��:#q�<7(�L3��H���<��<Q��kmt��P�6@=st0�j�|	�|c�60k���|I��%��0�L$�� �m�6z�$�VTw�ۃG��z���W��n�)��<4�@:'�r�μ0cX�U�"�Kn&��;�����t�7Ь#RBcy���L)���F������[�=�\��2�?�Ȥ����BM��WCx�U�6� 3z�L���1�����]�6ο��w���v�Q����i��Z�,������~Rx�T7��jv�h)�����[X<X�`sO�G_b��v�~p.�_���Nk��g�< Gth��Po�o����!WXqĳ_�uʔg�2��Q".6�BD���s���I�?�L����'7x���{L�2�r�ڶrh:n	�i,B:W��r>��Zp|zJ)��l�(^����6ς	�f|�H�ٱ[\����e��VCY��Z�X��9dw�M���>��Л-�0������VR?ܧ�6޶���CX=B�<B������M�+^	oE�o������4ֵǀo���s��认.
��"*R���h�JY��A���\P��QZ��(&Rac�:�l�&��&,+�uW	֐ARW�#5�lU�+I�N)А8�*�|6��Dk8�d����g|@���7���M�
ۙ8�K�
���5b�>zc��a�	��6 Q��{��+x������Q�"35>��\��h#G��ӟYB��7w�e�������w�Ƥ��6���!⼕֠��(3V��n#�*���9�$bЙh�@O��Fw� �� 퐭�5�1?]G��}�\�mr���:ǵ���Q�2>�͙���&��7��H2�4 S������p���s���F���^RZ�4����g��ݰ��B>ڸ��H������)����aU�N�_���V�1�lm���O� ��8�����"��3I�XO��|ɷ�DW��9.���;�_�/�`#^e+K,�w�c�~�)#���փ$�K�T ��tk��aV��ⴍw �Pc��K�HM2�ԁ~v^���2�G����»�l=���Q8B9m�Qt>MN/kL=̙RS� �>m�4}��c�"���ɉ�_����F����6}~'��[�!��k=�|+F4
Q�����)e����	N�(��R�:�-�H�]	j��
 ��`4�e߹�YfHU}��`�-�q��5�?Y���%�̜,������e�5��k8D��"��i�m��� z�=�;�ho��yX�_�`����S�����CKB�ݥً:@)�k/��0����� ̵ɐ���Ff2�(p��x�d�Xj�":J�
������Pt��4Z
H43�m����U��A�*fN��F�]צs�#�0 �#%�A��K���3co_�f9��Ikf�n�d@ޡLdI�c-�����k�O3��s�D��H��e��N�DC��䓏"�u���U�k�������9�Tt�п��PL4�r�jr$咍%"5�������$Np%��FSy�����-�7�BO_�����u.�):�VI}&��r�L1�A��&��јd	�/�e!��T�h�`�)��f�����a+T���\��t~[��m2��5�ա�Ӌ*�;��*�X�Y\p33s���bu`5���́t���Ռ�L&{(ȍ�q-?(�p9SX��VM�n�臟�����
�^;��yֻ_�f*���f�{.�5�����R��k-f�A4�"�"5������Ы�)SWl���Cw��j:d7K�m쩹�ܐ�Bu;��Ӯ��%(������4�MO��fI���%���Q�J�h
�x\L;�2]���1K�;	�ayˢc����+��1�Ё�wB���V�׎b��d�^�9��ֱT� Z����ϙ�p�����ֽM�,��=��i���V���w��M��6��B6JN�h#��#sł��i>�Y3^�[��J�
sz�@�*��k2��_mڶ���S5~�.m�^W��K~�ԃ`��2�J�j��ª�P��NV˂n���i����ə,�?��ms�Ԟ��)n�i���і�P��^��j�����N�[$/�Sr�STЙm.�MWr[8=� Tn����0�)Ă�����j+$�h�p�2����h��u	۱Dc��}���I�VطV{��܃��Qj@�'�"F�uyW��vd-����u�ьQ!�P�ߘƫe�i��G���t�?�
Fw`����P+� �n�͌�O'ɀkSF���B!"1@�sˊ���Z�{��i�A<�fӃL,YN����cScn��ͩ��Vg�9 /�sv�����$�����sh�잘������1}�C� ���,�	�0�U�&����)9
���u<�E�s�Y��R1��lz���׆yr;6/�L4����	�}��2���s�y38��>�G�2L�w|	a�ng�*��H�#jn�4�uL�@�@\��f�bv�s-�Yp԰�¾��D��|%��(s�ֻ6h_p+������X��9�x�:�ŋJ�i�g|؉C�3���4���X1�W*�,3��q����u��L	őB�A�u��c������Y�{0[�p����QP�m�Ј�����\��> �H�l
�Z��g��0s�!��Q�V��m>�kVQ��!�qx��L ��A���U��C�D�p�>X��w|��1þ5I�=I��A�T��+�p�3�>!՜R����	=q��q 
t+�A(�g._�0�?1HR��܄x��X�����ݤύbBl�y6���kwM�(�מΆ�rp��nȓ- s�rA��6fA(���(�q�V�v���D�}C�zC�]G���/�S���x#�f:!��W:���uc�"nmW��?���ͼ��Y璽d@�OVs�n~�V`��NE?��t�B`�����W�$�>n�����ɯ�y�r�-��1 mv��A�=⸑���x���� /���^�?d��yei��y��/��6s\="a/T[���&rP�9����6��/x�D���ݘ=��x���sݿ[�>����^� �R,\.%Q�O�o�*H��h������Ọ'X��ʾ=q��"�w��R&�h�%-Uh#Ա
��%����a؀x��s4U:Ca싰�ak㏎�х����0 �0�4DD�q{1a�,l_��΁>�}�E���4�h���w !q֩�"�f6S�Q����z��K��A�m�v�YÃ+�B�K�|6����^�Z���=+���X�#�&�ڤ�qFD.��2O=m�x_�7<��nI*�?.�� lE��[<����%�}'�n�I"���S˳ɚ���Ni�S��o�5d��{Z�	O��.����ɞ4�mCB+��
�6p���&�ڏV#G�I�VR��])�����\��:�u���rNr3��� ���Q�(ۄl��Ds;C����ں���炅����
��!<
���EZ�I�]�������#�Q�K�7.�Qz<F�`|�fZ�4�����O0�Ǎs��K�(�@'9��pIJ+���\�>�?�v@��b ��b�Pe����F��o���[�_\����y�P75�7��
�����.]\�?S�- d�4��.Kx6�+)�b��V",M��8�B��D�.F"�dJ�-���_�����̏�x����~�r\�0I��K��?`t^C��w�e���S��.��cT2�9l�M�壤i�.�C��2�;��'�9Q�R����Z����x�"(-ī)������NC�q�Uq�U��eo������嬌&����,��=�V�7j}���4�
|I%�cj�;��1Th�/��U@|�sNb��ؿ��獭6��4w�(��\N?�:�������h�p*K.r��'������q���r-��G���Zf�ټ�+ndKzk��h@��f�@z(���C�X�pa���G�	B���<`F�:a�[Agw�`k�u�����Us��N�;T3qP�v�f���L�>�|f�������6�T�Y��?�%�"'h�q���⎻����������.!H��7���^a	�3Q��2?˅$���e=��,��1��s-xD�%w\9B+����rv����ɻ;�k�� 4ɀ<���C��l0&ƀ��)�Ma���np�|*�R+�k��t��$C��TS!El��N,�9�)Q~��j=�%���$xI "Q��\��;8_��G�2�+�o�(v�Τ��~~z�/XL�aʇ�~*��:nqӲ3�����l�q��|���4��:_�X*��m�8�K {гG2��CV)��?.��X��P	��Mb\DNL7Ox�f)M��.a����U[SC�w�gL&������r���� w�������Ѓ���P�4�h3F9����<�"�m���DRu�Ϟ1C��~,��L�
�-�n����G>Z->�����wE'1	�l�y	�F�L����~�F�.���yɒӅ;	jBz��e����[�[���u"ķ`�"�e��r���%�Dn{����K(si�r�(�2������NSZF���r�j�DǞ�Mv�U��%Y�ΐZO������;d���Ą	��O�L��坞"��QpI��G��3�lr�� �f��|���\_�1��,��N���Ċ�~I�4's����� bD|,�Ϳ�w��A�.<��z�bFs�$�j��x�|�zR�,oabve����+�?���۸	�)��
��J��v?����5��	��B�1ҷF	��g�"�驹�&�#���1\�يU�Z�u/f�8�d�"�_��/� �z<]���R������G�
-x�vG�`J�6>����[����s2��>3�d��	 f��2�''�Ʃ�rH��@��ˏ{T��F���=J���-g�8?�q�L��/~�^r�T����� �`������s&�d�y�Gv�	��Oۘ�.�<@�ZT�ïNxH\F��3�kD9/�?dAg��.x)�P�v-��������wG��y>��r���i��Z��+���$gH���KY������-9\�]4v!�<�KZq���C�ȹMWGζ��Cׇ�6읾���	���1�P�b��\��͗*0B܇& ���n�Q3���@v����jnn0P(��f����G�Χ4������0����*D�~�Soeǲ!�:��3�Ѡs�䋄�,7" ��u�o#9�� �#��
�}�Jy!�_�/�ɞ���h�r�j҂ðN��`��E<{���.j��;[K �0`��㜕6H���ƛ�E�g�3�>0fqZ���0ӜATB�X��rDJ4$�b�V=��a��J���3���ƪP�s�/� ����7��Hۃ���ϼI�B[ g����W)���e���L��w��v�#�[,�։]$ ��x`���ô�l����C����n�no)���tu�}'J%̼���\�P?J ^�ϙ?٬J�X��$V$.�P�G���:�Q�ͫ�=���wYp�e���$����(
���q�X6O��b\V���ٌ2~���ݐ ;mh:����>�z~6�43�b���N�t�2�josjb@z��xi���}�ҕ��f��s��ӯe��\�c����~X����b��F�a�^�@��-��g���J06a��� E30�2�)�x�}���v�c�+�VP)d=Q���JfOjm1X�<� ʸ��tҿ��J��u�*[�+�V�7 ���~sbWo&��:��4���F��~#���-�R`J2�q��ҹ�r\A�BF����������9���]�7'�R�J���z��Q+���n�'.^��q+�]k7���ݜ<6��|��`�8�P3T%H�G|�<i���e��rL�6o8Ð���S�gY��t�3O8�S����xm݇�[����@��+�>�֣Ux0��#wƧT18�1�p X��+}� u|1��X�_���v�O����U��7-��z�\�n|[��G��_���'��)�v�AT���Q[�~�P��ă�����bS���5��Aa(����g����%ޞ����rڽ<���2�F>X �僡1����ԃ<p��[���;���0��`�ǧ	-�\�>:E���{���W�4O{�� Ւ�s��`I��H�x���s17m%�����&fn����U� �Hᇓ���3�)����ɯg�2$	�w�>��k����ο3���3�]Ɍ����ڬ����������vY���j>�a]�[7������Z�e�a5`śt,?�� ?�aG�:T:&����m��}��I�`���t�m���H9�G��Fw������J��}�+�z}H�j�v*���8��2V�Lߍ~(�$�G��sTf
V�Jb[����� ��Čk��}�!�z�Fg���-�髴��¶��Q�L9���E� �j_{so�X��Y���M�=a��ّ��}�@qbb@�k�8�<�ci�Z:�8/���A&vH��)Y��Z[|Н��%K�P�����Q���,_4�cI�;�		A&��}�6��n�c��J��Q�j�"P�#��4"��HS�R�׌�O���Vs.=,$���z�dr�v:%�9�?J�H�S�bqb��� {<�!ɠ� A��3����T���x�l��ݨ����MsMEA��,�I�,�*L���7&M����nҫ��4�%aL�dn|åLVky(lĺ�x�ڊ9��o�V��q�r��h��U��Ғ�����g�^�u9�o���]�u��QJk���ک��� GpQo�#;��h8GEQ'����F��G�	G��2z��/�+��L��g���%�ޗ�c_Ay���&���S9�R�h�|?��x��A*�� ��"J������$�2K���H����^���-��K�$"F�7��m�௴W,��p3�v���pqa���-.��M��/�7�����E2Oq|3���$JD����sE :,� *���ľ���ܙ���o���i��$���L��<�y�I,���c�I�\aƵ�AT� ��
��A�G���rNM��a��𦰖��_m�Ȯgn��A#fO�'�v�����n��ڕP�ܠ�[($���ࠡ6{c�nw`rL�5"{ �"x�@V!,s�����%^WDU&���rJ�s�#�v�>Z~:�Ĭ#4�)���k�:Υ��>
Xӱ�æ�\&�{�`�H(f����{l+t���iB�[�)��k���z��['[S%�ʢ�m@:�����8d�c%i���M�Ţ7�p���]�=�} ��������QB6���_g/a��ʽ+���ɦ��<����[ܵ2��T�I�bZ��T@��>#qf�|��t�k��#xd�*�9'U�C�U��@n�r���!��7����|mF�T(\)�˽�=J�����qQ1
�d�%f�����})*X�u���/��;�2;�!��3�)��2vS�hC�����}:���}ѹ�D�2z��18�/���Y'�',�I֒Qk�9R����&�X��@���+���C�ihN�DcFw熴VC�6�{����]1�n��7m	��#�;���w���෨�����K���JLU=�r��%�}�f�_4��W	0ʶ���A��vJWB;�= pa����,�� �`8��3�IF�������C8hBw�]��ω� d[z�84|������>;~�2JC:�'K�W�F��j����Fڏ�\W ;C�=���m�����	�v�s<��izܟkPG��S��;�[vO�!�֤=n�cpBvS��(��r~w\�Oc�p8�[�v�S�,��Vb���Y���S�5���S�Sޥ��^�e�,�Z��~_�K��4�Ĭa��Iz�M�Ԋ���E|�eBPɨ\W�lp�a����	�#xW������;��!�����qJ�'gr*�X2Y߃m��䑶�z��h��!5'HC.��PqZ�`��v����7T�D��S�����2ŧ�������!$�4&��X!�]o�8�}�Bk�|�B�}�	�f_
�*�9��EP�r�h9�60ғ��
b�֔����Y���G`���o��8�կx�M����D��2�fz/��R��������%˛.��Wx����؅�*�m6���ą��!�jz�5n:`D?�`��&\���M ��!�"�,��{i�PXM{<�>
D�D�<=f�7X�*_Qs���܅��O"��MU��Y=)
���r�5�1�%�<�+<�47EE �q���4eMh��P�g=�Ʀ�>��`S���U��;=J*�<���]R��/n%v9�w����?�%i��;�d:2H��:K�JDй�!��ȂS�$jt���J�E�Y���z�ջ4,?�\�u�-m2U-�`λ�J���e��pWbX�8(�������D\�lO��t��O�Z�A��F{�1YD��-��ct
���c���������=�^ g����@��03��O�@m���Ύ&>	�k�TԘAĲH��,0V��7�8A��܆t�a�1�C8N��6��?R�Ե�R(�sx������EgW�a�k8%�,#	>EM̔1l���̷�wr�s��n��M{]yXk{���byq�zC�l�/�r���b:dmM̃[im��jЅ�1�ǥ����U��*bk�<�܄)�hy쭫���s�������l��qb�����qa��% :��|�̪3���;�_���T��_�]v��5w15�>�a�:���
`n��lFNZ
�Ac�H���̚T���������!��5�7�߶��MR�ݮ�=��:?*&�����v�(�� ��?��K��(R� U�(���Q���Y�T��c8��G���%x�����<-8��BϺ�Ѷ������t�0�|�M�$�KO�j�ܧ�NK�ĉ��n0�Xl�|���L�7�ضB["ۍ$<'�FlC#3���x���U�����
���p�)���]W2���HU�r��H�n�}��e����Y͍����2�|�@�
��AKl��PG��Z��A��j1(�\�qY%�/�� Mj8�.�#o�]ux�al���	�e�-f ��+֤��y^�|�>��[�)bԩ�%�5Z!#B.�V����w�=�oF���n�����Ih9���M۝[&�؅Ƞ\r�|
��׎�����v��ۭ��&����xa9+�}�x�Q�Q����P�:7�q���=t�h���Hj9W(�=�J*�U���w{ךQ=��d._����0>�˫�>��26k�2d���2?�����\�Q/TQ���BJ�>�?SQ�>�_:+s-�$8��$[����ʂ5g� C_�;p$���[_�u����ᾎ�T���hT:OدҸ����v<'�(�����p�Y~���LϞ��/ۓˀ�vx��3Q�D$�9��F�رU�R5�Ȋ�ԱU���>�w���G���E�1����U�o�y�[�
C�U��\��[;��R{��*w3�W�1M�ź�H���3_��=����*<dhHQ�a�6yO�öb�[gd��#̋���;7ˠh�Z�_v���
�L� �UX\
M*!xg|0�=���^b�l�v/�fGű�K��w�u�;�o�>��c
����3m�ʏ2���0$r6[?<3��)��y��Em�K�X 	���6	T��������2B�w����0Dڸ.�t�f�s���	�x���=*|`�1Zx�lU�\Q�p}�7G�D���ɹ��f�{f۪��&H+��?�4���@��O��ˮfMc0�u'��E��<�e씤��k�k3ƭ�*ѣ�'����k!��슁�D�O2�L�0	$6i��kB�e��h�;�O:k4vӻ�W��k�&�P�w�:��l��ћe"��G���!�K@��$O�s��|��!w�)�1.�����������_��44P�}�N�#\����$�ݭ��)1��U�V����/�(�;z�r��-v��!���#�?���1E���>�{DPQ�ט�R	�\�Q6V���[��<(�6(o\,�h^#Yf��vA.����؉*"�>A����DJ�d/"k{5���@�Uܐ��V���B7+��#���~���;� (+5�`�%}7lvf�Z��$��j"h�坩t���ځ�̦��qwB[-m���I�m�d�:�U�/c�kD�I�Pp����7!����)��b^%��
_�G �f�L��z+�`K8�^k�Vڄ�O����j��Ѕ��l])��T��uR��d�mAw���A�Ů���l����)�3r�Y�>j��I̛���ܝ��?�gh��)j�����`���D��w�Dη��a���l���H�h�����c�����TWH����u\/ ��/��#w�l�r2�$���:%��Y>J{LC�a-P��+a�����M�1�����o��w2�����^K�����gn��׫جN����dR~�ʞq���[����k�v��S-/ߍ��N�ӢHA=b�j�eH���ć N1�	��LuS�,�����z�JF��-������迒 ��t��:�r,s@�1壅'&��G�=*r`�W���~GY����^�Y�tl�L��_�4��#� ��{��OV���I�����;�R08Y�~ tΓ0�ѯ���S��o#��,����b/�j��w�`���f�}0����y�������,1.���}3�ML���fr��k����4LՐ������B;�]����E�6����+ ������C�>Sd�3�Ǳ\,[�F�Sj�a��x� 	�23z��!%��ց���^"J��
)eGw#�����K����rL��'�ʲ�������-�OJ�R<Oꀀ�5��?���g&$0��
p��s��oSf�#ok75�2�D�d+��i[��~�Hʳ���4��"���f��0V�h��z���ub*�68�J/���b��1B�A��}rŹ�@_�����;���/Wt��D�q����X�3��Ο��X���@�yf�#s�Hm �5��k&u��@?wG ��=\ˊYe���lұ`뚢l6�7����U�5{O����F�^���-�.�<�(b�$��N��s|�A'l8~����w�TX�/m����|���4 A��`�'�>�_4`�#�b]��G��w&�AHIx	uj�q�!�V^Ԓ5�"d���,)����Z0�����
=������0��'�u!� �!������	 �ө�a0fJj����b��	E>�O[踋�6K���̑&Xv '�ՙ:]Z���ڷj*���a�| [�!���f��L��Ej.���{�n�R�?�8��|� 9>���r� �/K�-�R~�C��W�o� f;�Bv6��\`6�t�.CϮ}���56[�Xd��q$�����C��e0.��B�_x S��c�;�Ч�$O|��A����2%|܇N�7o���ɲ*��������N����꿴Lu?Ǽ�+;�B�J��Q���Ր���L/"��#}���Fs�t\)���s!E �Ot��~���<޹���$?IM�z~�4��#1w%�,B�+��y5(�-��i3�h�����=*{X�B行(7�P�������MY�$摆+<C��T�FF�X�6 ��qpwF(�(}�l���Ci��ވ^��ձ��PϜ=w�C��71��Ӂ�N���<��@���Q4'D*���W7��*59A��"	$ȱ'sݜ;���#�h����ɍ����Z��Z�8�'"�vPd#��yUf�&5���9�Y�M	�F9!�>�-[W��8�B_����.���Lv+8/��K�z�w��9� ��m,P}��:�*mk>- �i�jP��r�ɤz��_&�������\�Y3�a��ͫ��t���4��U��ap���^�@��=�Ɋ�ι4]	��ߨ
�D���f�E��j Xh,=s�g�ֶ�gn�T�V��ـ�{F��|nE�Wp���`�ï�J1�A�4x����w��~�SeӋ�)Ne��8-�z�3�AM¬�l�G%��=�F�'t<��BQe��B���s�Z�0͐�T�o�(�)X��|q8Q��(����sO����_q���P������엉��Ď����LC� � ]�V�ӧR������~��Ն�����-�~_�b�mk�n�7��cuY��S7(��.���"fX�'�u���s�؎�K�|�d�Ē���s7�h-.���⎡y^��kܖo �U�H���r�m�h��V[�@cs���a�����0����6΅צ9�5�/��Z�c:!X�I�٭���j45z�y�(7��OR���:�,�	oa� ��2ʁf��J"xXL#��?�2q���A�:�	�)��~-��_/?)W�|R�T[��̍Y�L瘫�Bk���!�͐�[y��N%�l(�����F2���+c��뻾Eej��yG4�=���\��D^�/6Y�~1�����:��������E��ex����^��s;���͎��?�d�G ��,�.��ѰO�"�P��P��-l,C��0":���c\5���Y<
GUm����v��(��li�����6�����H��u*��;�\���=\��o*�C5M�6E���z�-��#�ǫ���O�q"��K�i��k�}���+3�%$'402�J/�+����/��B��IGIot�Qܑ*v!u��>A9Jrbh�����η���Ѕeq�c��߶d՛�����L!�U�IG�P/�A|$�8`Q�QI�Z-�K(M��z.�`�/q<�}�F ���*��)PN����XB�SB�p�$7
|~�|('��ڊ]]�����Y���!ȏ,��LI������D���ō&^ >e��UZ&=҆��-,1� *!��й�c�Vi�@�#�Ysf�x��y�� l����d�5��1|a���FZ�0$�!@x�;Te���R��7 �l�s4〔��P� ������h$q�N�~��F�#'��{��1�!d����[��%{���+eEdm��������I��d�ʎ��C�d��7�1.�/�4�,m5��jK�U�ГR�^C��XA:{����9�<o��?1,*�k�K�����)Ⱦ�q�0-ȍꊨ*�b��`�aW���z�ޢf��E���O�4�	�8c�L��h�?X��Pn��
s^A�j�Y�S��ή�§�,B�K��/��%Z��}��s����7q�P����7��� cc"�����W�3�"'��27��:��ӈ�cXr��/���@C��.	�05u�V3��@�%`Gs�C���;6�KPD�Io���9���z��_�b�$�Œ��{xL��퀛��s��J��8y��J*�A�h�#��^����R{��/��{Q@�\0��n�.�TM6�6��Npj0:���e�J�����Vn�(�%�C�����֦i�֖?^l�P5��I-29�&��"�AonL���0���C� �l���+�t��5�L|�'@�{1�����w-�C��L������>f8&W��QV�m=��|Id���+�SҬ��oULֵ��6%e���W��dѤ2T����7�v�6���o����L��T�R�#8�L�KC'\��ȩ��.�8_ݎ���nV|xTMmF���GO�(d�ϗ�"�eλ��#��%Y��ܧ��x�3�P�����w�Xk9n�+����͟���3�}	�:aQ���MI���X��ih��8�o4�`_�'|<,���.pp�/�r0Y%o
�Q,�Ě
间�Z� ���ydGoz�9���^���+.">��b!�RP����f�W!y��SN$K�_2�gͰ���� �#F��l[>��֦�r� o*_�>J��7���k҆����+zo���*Y���}6�F�kB����N�:ą �2^2`"ݛ@�5�#A����5���Q%֕�������׬�l�٩ݑ�=X�\���4R�b"���'e���>�0�qD�j7���쎲o@Y%��%-�k�r��@���B�X��%ބ�?+Oy3��X1(��P�T�Ȑ_Oo����M�7"VG��K~a޼k��z�2ri��97P�c�*�hC����Sx8� TB>��o�A�`�3B��i�b^.~.mτ�F��0�$$"_�,��$oSb@Ӯ�Z�=���N�P;��Ɯ0�$�*��7i
YD�5\f���1Z"�L �I����+]�����`�Be�cq/&����"�x��C��t�I�������E�\y�K"''�����H�'�ݸD[3�o�{(�Ɇ��/�C�tT�	��:Z��/��<�1U	���Zǥ܈��[�)Np����ϑ�^�	^�ok�-*���\�I��e�֓;-]Mނ���YM�!��#�*�8}U�GDǕ���[�,G|)�K��3��z�c�;9t|��!�'�<|/�> ��	���Z�~�p��Ɖ2yGdr��8ױm�Y��*�A����/"&�T�zwxQ��ck<LPݍ|�V�/�^<��)�����P�lXIK�.��=!G����<ɻ�'�ob�=������o�,m���K��T�����>��O�˵�����i1�ٲ�V��=��9�qL��S`����-�������X�n�;�^\Oa���V	;��;Ǐ�ΐ	�A��F���x�rL�8�^�Z�&�S��/��9��.�ȩ4_��I�&%M2��u^C>��[N�2�"&A@PP^s3�Bc��uT��jR�gGw�|��C�*����'��|ūN� �h�D֊G�
�LQ��9�y�.�T
��:pV}�y6��K+LN�������%�t{\���v��)�(+gwF;�F��هQY�U��F��-��,��	DzX+�)��Rn�LO�(M�O��G���)-@q�&���01�]�ռۺ�m�^)/�m�D�l*Dw�2r��<��ǆ���oS���Y6N�k�a�^�-*~���jSI����]������f�>l|�G��H�P�>r�lF��t$H�.�v�+��9R�"�0b���>�)���wi���p_�/T��.ؙ2�g�����ڏNO�<��	����6��T�!�dfc����J�#��Jc�*��9���\|_�fZ
Z�����;����_Nf]����$��זH��e��6��&�!�m��b��^�췺&%�}r���
��K���;��p�np��k]k4�ua�,��o!ğik.gRCQ�<�����X��JQY��&���1�Q�6	!x̾L&�d<˶n���?�LP%�,��:s$K�!6�۾�"�`yU��³�8��!�U�YH�� Ibx���\�w��A�Һ�}`�î0�-��Yd���/�[� Ұ��:'�g��م�^��*dXްI�/U���䔃:,���㎝L��ڪ�-/�FF��*a���� s@%D�I
�����X-�7>�����}o��ؐ�{A��z��M;��b�Zb'M�kȒ:q��p3��a�R$�xt:*G�)<ʩ�J�&_ ^;��F�S�oGX���d�Aj_�o�
O�l��'N9���G�hv�8��b�Y��S#^><�<��ê�g��c�I�~�BC��r5�p7�����jU�a��s��0�����rRQ��#Jκ�/^߂�^'Ӈ�Li�kf��=T��y�TWe��lL%�۸gN�̩pG/�����
v&�adRoV����?��w[�k2C �c�P�$
�Hء~����^�hb ���^�
 �#O��Ư��')�N��
�Cw�]�AS��څ����G������������trCw����F#�栓��M��*etI(^G�MF����xl5��Fɡ���J��堛�3�86�}#Q��KU�B/ن�l0��?��,Fr�;�D/o	P������W1��xfvn0Z�dO�&����P�{�6�'��Z�����3�w�u����ַ�W�uLX�k7w����ӟ����M��?���V���-SS���Ԩ��z(����K����Ft�S���`�iϢCk�7_�:Q�#����������iS^9�j���

��w���'k�{����ǲ�e  &����F��͜��T�<�:�7��O��!K�?T?�>1A��\�� ��0fzC�m:�o^��"��}���1�7�;|��b�:b͸���B[�8'���!4������~�Sÿ�!W�E�1Ǯ����k�\�=�'��'Z���zŵ)#���쓯�9CO����(Ű�Rf��t�+U��ۚ� zҳ�6�j�FJPK���*9�ZF��&�XGb*���� �rt4TĀ8#�[�v�= �Z���y�5^�4��Cd=	v��)������Â�$�@B\�iDP9�U��"x�.�^�Xs8R,����ת�jj��s��F����"=�z�Fo������?�=���@|������#���i����x+��	]�b��}9f`d��Z��7��p�-9�Vi�Y�ўt�V�k59]Iw���H�.jݳCrjׂ��ݙ�ͳs���&y�o��#�	$�κZ+>�T��:�-4˼��!��5Fh�]����,��}���8��p��#I�ʄ��f,.t��8ҾޭI�� ��Wz������V�ƺ����ty�,Ì˞;���R�u�i<���Q���L��Q��t���XՆ]>�=�]G?#t-����<�����<�f%焧t~�5�7���#���t��ؘ0��5*ѹ��X$��u��N]��z�Rr>�1�"m��
Gx�N#(���Ԏ({� ��� ��"4��.4^���f+�V�����k���(�����:O��
�9XY�`R56�#��ԙ��R.����]�K��|JE
�4f�H�nP��&\��b]^"}�r6q�ZyV}j�&�-wr���������~GX*�"�����RH=��`�.��|��/�8�>E^��a�D�!�����3��$�����+K���,��y�1[h��b[�ڳ�%2A[zՎY@������_"��h��(c�v����P$��XQ�-ZV��ۍXZJ���U��'҂޺�e4��{`8@�5��{?� �:�zp�Dc0�^s&}aN WD:ޅ���̑� [W�R_���Q<޽���b>��8���[��(�#	v� q6�)Gcd	��헙��,T��p�L]�.����Ut�L��,��q���+m���G�E���X����5`�<�w�x��%;�f�я���7�B�@���C��4�F�I�O�{#�~Ml�G�a���(��Iɸt?��:~,����C�S*��3!�)u<3��Zm��Ǚ�o���X���d�،Sgb�S[0�e�c�>߳�Q)<�WU}��U��u� g�N,�&�0��ʆ�`��<���eb	7���+` ��F���K�qu$�?ǎ��H�2�_R�=��Z��������R%�;��s�ƈ8:����жI�/��@85@6[����8��܄��PW�x�]�ƍ�1d�@\�IW��H,nl���qP7�P
�⇏����k����1����ߨ�ݲ���.�Ѕ����߻����b�{1eś�j� \�q��n�0QX6P��ɘQ�uFw��D'�<�Ҿa��³.ۥ�3��ԭT��m
�յ�x��S���s���vB��N�!L��C�D��3ٲU����s��:�Jq|;��+�g�۵]z H����?��Ҕ�͞� �Ofs�'=ZK��}�64V���_��tw4�T���U�M�HĬ�[��]n9~{]�:��[e��:\��w�#��O�ګ��u����bg�>�� c��U*�-��V��/�k�xz(U��o:���b�N�\�&�}:��M�/�x6�X��p�����~�h1Tz����m�uز@yuXQz���<�����G������5;�ݗ��/a5+S?`/�/v�z�0�q����N��W(۝^gsL����b�s��9��+�sد���":�P�>��ap9qJ-x�s�#a�v%Eep���UH�Q�_?��F�之�<A�H�[ω�?\!�yq���pz	rn�A�����o}KU���b�go�IpFtMEnz2��{"10��_Ë!:9�P=b�z��7�\�vt�!�u��F�J��"49�|�����Ic��xg?�dbr���v�,٩5Y�#=���kF�BWQ�~��9�����D�-\�������ث/��k��f��-�a�1����n�����}5�ok@bsf�'�@̜e��jՋ���7ӱ%<��Q���if �k:���5�ע'��� ��eF���d�Z��A�V�U��߀�h�xu{/s2)��)�SZ������]�������$G �u����6<���Eg|PN���	�������	���oMz{_	FpR0�C8d��B�gk��{�5�����-��!�E�`��_��'؜�e{���ZN�:��G��D�+c#}����ӵ{��L��Ǵ��AS�Y���ͺ���/����m��==֡��M���ɪjoW,t�8"D�3�l
�C��NT��.����^�^��=%`y����?E���U��Լ����&��n�27?fL7�l7K���K<<]�qw��	ђ���92'�6<��+M�q��NT2�^kL�V�ex���G
�mX搣Í,�ɚ���0i�b��W�5%L/�v��(�
j��U���n�ߴ�+�fd��{7��y\|�}�&6[ ���l�j��խY�7(}��/5��J:®����_��Ԃ1��(!�1,��u+�~���tbC�gd��x�JI~����ՈEAC�6���oϕ'�;�41�`_u�8N�Q [�3G%H��v͖���&[���x�bǡ�%�ߒ|��iOX�����g|��e.2�� �W:h��Q�Μ�`5���r/�6j����6]��76,6	ܪM��]a�?�ule͒���u�k�|AYSlk�}�9��g��E���r��x��8��~A� ���p��݈&��f�Nc����	J����d��8���猪\	 t�ߑ�"9��S����b0*G�n��CZ�+n0���O�| ��2�Rf����Nq�R��'�ߒ�>��,��m�
���{Z�k>��IZ�o0��/$R����q:d��s�+�K���,4��LD����Q5c��5+��y���\o~Has�˿sPj�Q|���P���
��坺���f�	�w�e'5O�]�>��dLt5�K��)�p�
;��X�s���X�)�1�ԁ��\ `D	�n"zZ��<�9Xc�h�Y�}��zq�FB����=7��.K�N���5���hB�&o6$
ɧ�pԊ�d1s�nr���i��4�[L�잓6���V_�J�gZ7ZY qX�\n8�vޥ�W����#�ʜ{ZY�p��]�oh�c�Fڬ	y��j�T��cDU�VϽ]|�M�
��3SШ��lft��8���DU�|e�:�gՅP
�ŷ��eqS�6���c=��/-�į=�=�o���0���\]ҾN���ߣCܱ��]��=-�w�Y��7�"{�"���9Q=�z^�'���S���K�dT�ҝ�X`����hz��&n��|����x�Y��P1�c>t��]�W�;���#���Sg��P)�<�h�����y���`�dR��6�U#JA9ɬ��\�u<f��=��m�'@SU�}1zQ�T��	����b�vZ��:2V�0�p|W�{پ��%C0���>�b8�R����s�a�M��
�(�RS�3k��\h���<f�1#�&m��E X��UEm�d
���V�Wo�0u��FyEr1!
$ꇒʜ�q`�uB2w�6�\�@�L~������P�	��+ֻ�r-Joo)���(���;Pյ9V����2�[��bD�H�J�E����}�Va��V_�P����H�z�x��jo	�Es��!�2��ں�׉��"�ޖ����ã��֌����Gt�N(.y:xe\���/���y-R�d=�-�b !u����z�i�ӽ����P?�N�誺$S�ؖv�5�a*+���)m=6фP�6-�/[ksC�o��'Q�<=����C���f����mU�v"��acD� }%�ޛ&�v]V��HK8��H�N�엫�����6W��~��P� u�ŐE2�)\�W���STg3&���Ԃ3ˡ���%���t+Ir$Qb�v���=����`��4�e�`�#�9+�;���?�E�r[�i�X�����ȿ_._=g+���ʻ	/K�Y[�,�����
N]�v�P��H���p�,lAR��VY�V[�7��=�zn��=�j]/�ƌ#�9{q�I:�uq�W:7�m��j�'y]ե*z�qŰ�1�]
�#��J��W����%.������g��3q����ּho���df#������;�f�z�T�� �{��D�(�5#k�~���1A�)�B��o���.�)�|���1�!�����>T�w�����Д�J��ǩ�Cx�� g"}�Qb�H1���ۘ� ��HZ(\:�*�#g��W�����S�\iIB�\f�>X�3�I�СD7��t��W�7�e��I�ҨM�.�j�H�Vg�Mn�O��coB�� �\�s�>0�G�:�~ft4RI�`�����6刪��C-UQ&�J���ˊ�;̎r+a#�c�K�5�AO�̕�-_��˕LV�v�Tt�����ǋ���[�J��U.��!��1#d4��ռ#��1/�Y��Q��
od,�Ҟ��<mB@D掦Ƅ�C�W���#;� \�[5Օ?{�@�{�7K\M�5[m��0�޳�B0��	JG���=)ik�q�_�hQ���^�@�K�֧�c%��e��	�=�C����Ș���nrΘP����7��Q��[_�RrNꘀ�����z[4�֞��)(��"�� 	0�;�m��Z]l�e���>,w�m�f3�><�9�7�+�T5��ɪ͡���N1���\@��������tl=��V7�g�ň���~��%G�|�y�q��م�\��!+��q�/�]�m��Gp�͞�R�5!�+������CL0�V��~(���=%ݗ���p琦��
uq$�y����;Y���	��:������J������Y:ȗ�&���s�,M��e@��� ����
���B�3M�xS����4�T�oBW��SP�C��73�Үp���m�?eQ��oK����UԂo�T'��V��lN�!��E��幎�PSZ��!bT��rv��sS�ӗ�ʇ-�r!�d�_-)(1��=�C&��f��u#^�yK�UF�D�������h֏%���W#C9-�E�r�A�?����l*�y�~���yE��tl�t)K7	>����6}���4��f�xDӢW�W`?
��pO�S���ˣs�ӆ�S8/�@9�5_�ܔ�[�7Ɉv���+��m��ѥJ_��;H=4���仯ɓ�́�)�n��p:����jKiRd�P��o���w{m����_��1�ޒY�5Bϸ���VT��\2Ϩ�̑%��c�a���	�������~�۲�e�Ud�2#�Ǜ�I?�9�e�m��c*��'�G���8�+M��Y:���mW���?�>��(j	V�S������-�� ��wZ25�P��3.�����:�H9�?��*��39�U8;�g��&l�������ed։xx�3����BgׂCĀP4ܘN5V\�y��`{���#�p��fz��+X%�EK[�\���e���TK�1d��V6B�����T��MG��-e��(��kZ�f�hp�ɯ�
A.}4�B	{�:�d����uKg@�i��{�=�lr3�&.�������oCb1xw�V��&�a7N���<�\%�Z,O�G;��������x8sUo�e��d���c��n8X}8���{�Z�z�0��5�\�:ա���-��!��$}�1�\;k^_RD%+h�f�����҂R^�����Ѱ��������x
/�t�^28>��l<0�Їe���$y��۝�:=�d}<O�i�q�CSע�yƚ�΢�1��%��;�%�_��i�He����s%��<��=��6�?c;�����f�]�ł��|�F۠�\y3^ȹv:_�$�L�#(�&>;�a��"x]}�&X� �~�AͲ!h�r+w�1�8�$b�����\%�%`R}A0�@C\���h���Ϙ��x�φ�>pBC&jP*�׾�wa��8!�ϟ��?�+��ò��t���}�2�XLk�4�ؖ��c���O��=w]��X�|Ի���%o��!>3ɱ��\��|-����S�E5�#��82��qH}OIӑ� ����������0��[?a����k��O�3����܀�� =v>���#,��N���m�)���)o��η��� &�8�:�ըQy.'�|�����Q�1�������jxB��y��� ��%+����T�-7�-
��R�1�0i�os���Hv[�{t߽Q׬����e?J�YzT!�|�pv�},&[�S@�by����C�yI�>`R����t]�lS�0F�Kw��u�6�/�,��zn�q_��׹Т\���l��Pכ��rL�ږ>��[�(��nz5���ᗌ��s�T�l�8s��l�I��,�^��&Z�ݏ@�l~�z�C�ػ�N ��3�}U፶x��x'+�D�Q+�x�u��G��Jy��x~��5�����	��&�`��:F.�(wT�abD��D-B�Ҟ�14X��t�'�ho]Y%g��d�\�fCl��i���ԛ���ߨ06�H�}y(蹜��Å�\�;Dk�#?�&E�g;c�����:�I������XWSġ����
�	����F��e:�����V�J����	��:�a���aR�G���8�w�H��i�NY*�1k}���LW�F��)��HB��gp�Lޱ~���!/ͯ�sMFWL����u�o2�S�A��q����2���8,Y���jpVX��'ݏ��$�D:�SC��b��g�O�h������t��P���4���/?w��o��B���\r��^�wҕ����d�7�r�h��}!��#=��y6omB��xD!��͕���},~�L�B�F��G$F�^%� �+zr�;���[�6�ֽONK�#5m��&^�9�i�onc��qO�+Y�	=g,^�o��&Q��qE�L`�OY�E-~�h}+ٺ���t-I�#{���s��w����/st���2�NM����ձ��O׆&.+���I\��hF1m���`���� �
B�M!�3�)���i��ϼ��J��釸|�G��w#�*�N=b�����5�E^�"2���)lm������OU�8�1i�:��mU����]\��;�jn��T��-ђhv�&�\��#k�����]A@�![ɠ&������q�x_����5-l�wݿR�y�J�z�� ��;�5��&b]ho�Ό:0� �#��UUSw�/Aq>,y2V(�f�K|���@��2 ��`�K�eq�;��V��Ĵ��,1?��#D�>�8�m��yH�-9�*6�|x/��E���S��{s�U���M���]Si�Ǫ�2^w�~��V\�Ap�JF�����ʫ�B�B~�"\v����VTJ��F{���R7�����<�Y���~�:U�td��f�=�7������>��^>���Ӛ�?��p�>�烩3��u�����f���7��
�o�<���PC[���h~G�RٴM�¢��h�E�t�[W���T����vך�bu&��}��g�$�՛�z�S�}
JhS; �wK���/_S>h�b{yi1Y�j��$�ew��#K������w')�&��;���X��j"�U�����F9�S9�H�����Ķ�+�[�Ӊ(���I""�ӐtaN,.����S�Ӂ�_�'&ŋس�+��Mc�u��-E�KW4�?�%���hԑ")�y�J�1��W�����-A{o��%�nU�UNDGLg%P�#��Q�^;V�J#��!��h@f*�A���ŧRjO�MvJ�����DF0R�F~���M�
���ov���80��N�}�ݟ�)�vGHP�j���Qp�PŲ���5#�$gbmܔt����o9%~���pZ���`i��} ]�,�tF'��a�_l��{��y׋d+�����7� >v�q�J�0SBT���s֬���*��e�vy�8E��ְ���l� �|<�p��{�ٞ!I�#[y-���،G�C1�yf젧]�Ͷ�ƣp�?�&l���J�(�)ز�X���A��U{g������f	GЙ_�u�kL�3Ñ�"tjr���� �ſc����K����nQ����S��l�rM7����iȂ�O#�s=xF*t�աj
*�N���N�=��4Urmօi�ؖg$�'z��= d��LԴ������(�>*y�t�ua���ɇ�Zy;_a�)���~�*7���T�sRa���k(������
9X�i�+Ǟ2�Kl _e|��)��p�ѣir���ͮ֧��ЭSbch8�<���PI���ո��n�Z曧��(P'��"�"IO_7��V������|�O��Z��Oaw���
]��5��61���w2K�Ms+F<Q�U��y�uQ�o0&-�bۛ���
��+w^���f>,ME�����^ Q+��$��{ �I�~��� �)T�y��(�����o&�j"�,|���Y�q�2gD.^���MA���=����ٳ��CMl+a�U[7b��r��7� -w�����C�^��6:����;� �UK]�gb�>'���߇|~�@%��ɊG0_��3����x\�j�[*t��;�?nB���|��J�.R��~��ӥ�E۸Vl��7f��j���Kp�o�}�y�يe:�QI�����.�Pq�4�_T��u�/lt����d��7)`��#P�z��*8�e���!
��~���`ҫ��E���ə䳡l�H�~��Ȫқ�f�Dl�˔��7�*2p �h����!�D���ͣ�C�@{dt�j�k�����&�#�h���� D�d�s��
w�t�̆���=�!ʬ�<�al��>Ѵsɟ��O���!�$��XJ�f��f`�K����.�����.��I_��Q��Ч���a�j���Z�,[).��	L���U�L �׻ȋ��E7����𺢮��/��+`���߱�k�op�g�[q�t+	�6��	B�J� �x3�װ�&���Ek�9�__�	�_9vw<!g��	ĥiH�Lv�!~s�[���ՙ�# ���Gɰz�2l�JH"Ή	s-�J���p�EP������TG04U�]R"�ߣr��Gg���2b��"..�����by�t��V>q!��TPr�K����ft2w��#���rM�Z
�O���v��٤X�ĵ��XJ��'-Y��0������Nٽ0x�Ao�)hn���>R�+w�FT��:x���|��a�~�Q�h(IGh�&m�TR"OeO�`�3ihs�rEc�T W��U�̭AjT$`|W:E����j�=a��3�	�Xcd�%���VE:A0^я�hܒTfj��r������1��%��j5�4.|!�L���|�����Ȅ��L�;�����n���f<�]��9翏^�U����T���Bܹ�Do��پ-�H�k�u�8�E�5�������m�q:�����3x۾Ź�z�1����C[w��fQN��� ���xgӬ/��B|���l��Ϛd�T����EĔ�O��N/Qb�zn{����t�8hF5N�D��L�L��9&{��5�������I��L�W2'p�J�
Fg*���l�q#pkH� JNL���>6��L����~{�� �E���������ǿ����A��Qcҷ�Q�z,Ƴ�N�;c���t:����p����I'Ʊ���;�0�����Rtp�������܀m�货�jQ�/���L6��=�.v�LN�~��<��n�H�;���mK5���Q_��y Q/�"cm4Ɠ�`>(��`��8A��k1߆��c �A���F�u���B��0τg���R������hY{�!��vHq����Ў9S5Cf��*T$��N/����Q�Є)j�a���ǌQ$��*�7���f cf�ko�V�M��bx�@^8�����^s��7RI_5�Z�a0)!�W�F�6�Ie��PP�:����Y������S��W���R������l��R��hѺ�i�g��Bw�,Fk��g��T(G��7�V���^]�3[^���ho&�;��k�w%��o�Mq�K+����'�hC4	
u��b���N� h����N'H�#ᮦ����=�:_�5�@Fy'.�-1�V�JVI�Ÿz�n�+��56.��#^7&� �h\<� ǭ>�;��]����Xx�.ۨ4����Jsfj�Z��|�f�����h��L;c�K�[F��|���kWe����	��V�k��C��k��1V�۩�16�%fZ-�������b�2��J�"�k�t�I��~h�pA1(����,�Y��b�H�%*n#�g�O&�Ϯa�dK*���1c8*'}R��_ߘ���6��dp��C���ob���c��c�K�q8n>)]���.���wZ�v�xn�������Y�Q{�F�_N/�#ﻝ���h�g�6��ΣN�2�L�Ȕh�5�.|:��I:[ҠAlf�<��Ͽs	.�%d62� ��1Gܑ��feqp���/	;,ƪ`۱Y���}��.v&GgB�����@��Iex��_C��˗J%��gTW��1��W��0혲;�� V�H���=ZQ�R��L�qQ\�sc(ްdY�Al��UO%,�����]!jw
��α�ܾIjpu����>�XĂ+��i3���	|cEo��qȖe8�;b8M�/ʫѸ:��atW��BWԷk����5$�x�c�L����sZ��*� ����,l��D�i`�tv����  ��9��ʉ�P�ó;��'�ё��C���h���9R�t�[���įvbCr��V�J�xN�xD�����Șx�GH���*�4ϧ�ݓ�]1_�3���/rg|NoT�h8�QW�i�Z��#��F` R
qڐ0^��c��	��= r<n��l6lg{3o����jFYH��g�E���G�6�:
5�oq[� ��L�ICGL3�!�dN�q���<��B�z�+��)I�-�L^e���qy-�F��]�< "c怳E��1#��%�Tv�}V5÷g?~���lF�n�cGr
]�w9/�MN�8 �=C=�]�F���O牿:�����V5A���1������!�-!M�G��|.����O_�pU��4�۵0���VR�ԥ�N�����Rmu>�Y
UA��y�>cı�H���c�ޥ�:�����?��!�B���7d�6�(�ldM):�j�C5�Q5��譔�HJp�L�6$����[�Jb�:���ep$Ԃ~'u�c�L�D��vn��}����fc���=	Gf�Ӻ�g$��>��awd�S����F���W�ן�cLj���*A`9/�2P�F�	��~pb�5� �ߩ	\���+<�e�m`W�}�ڀ�W�[6�����8V�����;F�4�Q�m��z�Zr���P��R�h�,X�� ����8�[�>�Q���IR$h���*�Ť )�M�]�AV��%w�����/#�`�yə	�3>V�F����Q��H=�kz���}�����J*Y���J��
�$���)��z
����%�+�Y�H[`@��S���#O�}}�܊ڦA���-n�K-l�H�<��3ug2D��u��W�0��J"��~��*�Ο�ޱ>Tp�T5",�2����`�Ċ�h�9���Z�ٍ����RЪ�� �?�W��ɇ5�Ѳ�&�%
m��^���vO[��4�Ɣ�[P��H�*�.��' ���#��zm�Ɯ�>S����Z������*���C��)pp��{��Y3X�JULE���HN�I0ĵ�n�c ��G�Д8*������L�S`9�m{&��V�#Γ��<llvw_ˣ���ټ mc0�x�'��<���7N��c�3�D~\����ڒa7�����3,\����T˄�<U�l�׻D�c@y��ƌ=w&U~�q��MM�0Z��}q�;����Fto ���4U��8v�@�.Q���/!a����AL�N�� �3ľQ�����"�8s0�xѕ��a��Z9���,��N��9�����P竚I{XRx͢���\&�^|vt�֜���Hr���2>�'��x=�d��foT�X1m���7gg[�x�G�����?��0����
�2�9}[$-4)Y� gW���:ߘiZr{����iT�^�m�%��~o�9+ۚ!��N촡��UI-+�$Ɇ��8�10��m̍ۗHQ�e� Nk,g�F�����v��h%�3��E�-���35�C@�2
w��6P!ӂ�Ge�*�V��Q��k�/Y^�?9b]�d9�;L���b3ý��N'��
��AJ<����f�k7�����v�Q�k���Km��41����5��U��K� ��j��ѫ�O}d���ؑ� ������Ł��cDi �s�Ө�,	���r�W���D��¦Y�Ӫ1�r̎���ԃ���|�LՁ�����r�*��A���ԟ~t��E���^��V:t�&=S�"W��+���4W�Ů]t	lIFBZ�k��������`�	�&���&O-�����k� ���|�~����y1�G\�u���$�Ŧ�c����7%��~
"'7� T�/��0�o$��:ߜC�[3bp����q`���4`���!�6�XC[誟�u�p���ϼ_��d�}�����?������Ni 	�FDy�������#�a8�c�,CҎƨ���,��p&�?������bV��0��H!���~�a�̂@����'I�[2�0�,���j£��,��a�|�^[vF�A�e�6����C��[�/��"Q�8��d��$a����N08B-{+�,)x�3����Li���'���pkg���E���c�6.���=WF��U���/ݛ�?����WJ+����u�J��B�V�9�n���C�����kSS ĩ�����I��] 4�2f�xs+���Kv<a�o���TB[e���~PN�0�ժg�z�Ar/i�Z;?x�q(�`iS�^�ۼ�2T'�haPL��lh���J��$��qA��8B�A�����px���?�B6:�}h�/��'����f�U�g�V��E�Krş���v���zXW�u� 	��Gt�?F�#��6�u}獣�I��o_���X=I�P�������|�U�ϥ�D��]SS���$шG�z#����Ή��w7Ԕ��x� �V����}�U���T�c,�2��,)��ݞt�����_��:�+�h�[n !���A��yȔi�,'ᆢ �x���OsE U���u��N�dl?�o*d��
;������i��c�����YD'���6o�I���kh�;�s[p�Z�3��h~R��Wǡ���ki� �'�\�r�y��%�q�bƷ���5�aP�W���o��������C��{�!P�T�V{t���5Ƣ�,;8��T���C��ǰ2�7Mj'���l_�����T@�_4ֻ굵G�d�gY:� �5������l�v!		�c��*���ͧ�wvꊙ�ЉVݞ�|�n6�FCb��6�8�i��=�/�]�G�g[M��o�û^���|9Prd�Xx(�h��z����f���[�s�2�x�8��ƃ����~%��X�8C���2W3��#N�~��e�-/�h�&�?M@+M0�}�{?�����/�N8�wC�b�|�%����/]��������җ�S�U6�!��X4p�K�I[=��ї�{���0�k{���X�,c���q�~���'��Fvi~M� |*ZzQЇ�V��#�P��M��<�U��ԃ�[%�e(����.<`��h2�O܈[q����\��3ᙜ�͇#*���Af����KGq�Q�6�8��6��a�6�D9e[�0&��͠�A���C��8����;ؒ[���HD6�����#UKƮ�-a�{�[�#���i���}���獏�L��(na�,��ș2����ƀ����4��r���j.,\��3���O�G������z�j`��
@GzF	mha?����v0��T�X7�E�d���hR����0r�.���ۘQ���L Y!�;C@�����Ln�6D��x:_���h�9�A��t����	P��6h�ܜ�$�)��u��^)p,G͉{�x���!n'���fT_�H{�����QRm�f�N�
���� ��Hs�� �dn5���L��4M9^v�� ��p@�L�ujy?*Rv3_2����H�����Cސ��3��E����<H���#'_�]��'[��R��(�'��vwYz�H/#�<�����}�A��k�*e5�,ͪ��1�'IZzQ�5r�LuU��=�ߔLk&lr�g\��q�׫r����𑤣���(L3"ɠ��7d��Ւ-�IdZ����"$h��!�,�5���J&�te���O�|1�x�g�P�T�G��	/?���G��1�)�Hh��"�ݦ�."��U����h:�C=�9ݰ���m5�1%0�IisX�=�w�˰o�p�9J�!S��`���lէ���g�d���1�����ȟ���_@�Ph��os��w!�jW?�������E�O��쌒��៏/��R����te<go��y����M/�X]V�C}߼�0Z��[�u�5����В����{M%;t��q4R��eW��tƵ�N����[���ŵd���h3���<"�q���^p��`T-Q�;�U�yj��m��!��q^��i�@7m��qػ�.d�E�l�����ā,r"�W�Ԭ�7�a
Vp#u�]�5���u�S2
�3�
�+U��W�-7*ryZ���b;�zd�<�<��i�ط�u��W$��.	d�n��,�h^��*S2�-�������L��L|5�6O��6]"� 9RI⋵tf�X���,��W$�s#���J�:�Hm��)�~p[��5Z��N����ڍW.;\�2��Ơ�E:�d��2H���¶�
��*�<��J}�I��oY�g9ݥ��L䆹�,�հ8f�����0`B)��ZKb���䯌_�L��HA��Ϭ9����,���7Ua	�S�CC�X����]�`��k&��ô�25r!�P��p��m"�T��"�~�tX���$3��6�.Z\Њ/�m�uW@CF|-��ȝ�u��jŨ 8O�d3)�:�m�"|ƌ�^��D񌝰CQm�񮃝�x��^j]ׄ��SA������[����B(,͔�M��mU��	e�����L�����T8�����A~�+w��ߥH~L5��^�RM���3�a�"���[1��Z�M|~,�T��G������}=1�S��\,�Y���9��O_�N}��4o-�ϟj�"���TOV+�6U�GƆ������?�ׅ��y�н/�� #=�F��� ��6p��}�O�W��"���)L���h�J��]���B�!��n��kT�s���^�Z8q>@�Dr	��ѹdk�|�����"e�T���\%��i�JKg��|����U��q����y�&$y��D���~p��M�ny�K%,K��4��y	����Bu���eP>��鲢�2B�r?:�����r4�Pal'�����G}\��-�UqT
��29Ies�EGM������r,��I7`)Q��/��|M'����کU��Q�9�Fg��[S���K�0�����#���;0��6'	���S�?YגZ^��`'�)�)�ĖGɽ]���d��p��1�4�����?����m�7%���d�d/���A!K'@(~6^�[�!���1؃���c�]ۥ�S�t64ƙ?�6��@��>��r�0�IC�N�(x�J9m'�4W��'��z8
N�E"f�	�q}Z��"?T���YG�E��h����K��{�����8�OяC^#/��J��Izfݭǭ�h��������L�@9��t��H̎>�4�-344��rS���H|��<��s�c4�+2��f�8�Цپx4\������^+��ڪ��0���:�ˇ��Z��v����PX�q�qx�����uo������A��H�nH�K�Ԭ߀ݩҘ�&���~���vc�AV&�ގB��FE@���^k�V-��XE���(�{KEh���t'���3�bo���>a��у��F�T�r�kp������1��N5\#�I����������.��O�겳��MHP�g�y�,� ������,���ﳉ�S~�9�L�����7�m��Z�ha��i�iCԐf!�h���J6+���=*8�'����[qxJ���p��yi����n���YQ�k� W�Ʋ����R�	d��|5iR=�d��g?R��8:��G8��$>:�.3X�����U>vC%IVPM�Ԃ	��4س��\���3ʗ�ȥ�^�����^��|[����;�qy����̄�"�)[D�����[��$�V�1��e����R��k�c�5��d(�$F6m�m^���<�Ⱦr�?���٫���q�+��"�V+��2ک�+��I��f���:�?�(bk�K+/�CM�nv/5�2!��Loid��V�r%�E��P$P���2��z9I96pd��Z��Z�G��=c/R�&c�-\��GSt����>�"��$�����Θ��$z=(цUm"�A�@)�էs	��6����e�ޭ�� �U��ZO�3��щ�5�T���Ֆ#ֆ�����x�/�^�C�5'I&𫱑�ԑ9n3��o[�9�/n�c�����Dy�R�J�=�Q�.�)�RO�@��y��^��Ҭ�[���~Pe};��� �xr��PX|$VH��r0ڕ}m*���&���ߟ!��P ?Y���A�1�C�m��P�������K]��9,�&i_���'�p
�
�9��)�+�.y)�Y��YHAp
�w�k2LN���0��^��1��u�����E�n�0x��M#8��&�?ݑl�����`ћ_k�D�8���1��n<�['.��$-�z�5��;��=Y챈�F�TÕX�s��p�~]u���9r��e���=[H�$�]�6K>�CǼEEO��u�\�n`���bT2�D�v]����������*:V�����t��!`&��������w���7k�*	�0�UkP�m���0����
�
��Z�f�I�J<tl�Y�ń㷼�H�9�Vl�4�����]�R���g��¬ Ⱦ�~�����oK\N���ﹶ�1�n��|�q��zI�R�3��H��t)� �^�8<�:�J��lw��c��a���6�<O)�4����"*\�҅�z�&��Ai7^2��W�_��l�j+!��,�U`���=<H2�j��O�i��i�ɋo�֖��Q��\�YF��Շ@	آh �26��w�Y��U���KxkrP���ˑKbO�*,����,,.�8��v/���GyY�?W�>c��c���T8��[���1�KӢ��aL�S	ne����iXIŬҼ�\�ј�y����@,w*�G�������d�7���Y�g{���;��O�����jy	�rj��&��}:��>蔬���Q$FmV.&7�(�<��	�Hpy+��Dz�P���x99b� i�R�����3�����e�7lI�d�oچŵd�ʑ�GQ]�����*�`�|룲E-�������5��$y�����;���qo7��:�?�s[�1��\�EՒ��P}:�R����C��]�	Έ�h��>\���A/��f��G���+ z��`PD�g21�)[����7��+�\��3��?
��e<9�L�:��T~���Ȥhm��ʏ/ga�*ְ���Y@s艖R,������Q���%��F	/#I=��uk��տ�⅕�G_�-�d���7fܱ]�ێ��Dgm@e�t0*L�D�~^�q$��x�dT�����t��StY��ۢ�t1�D�D	�A~c��3��,;@#��k@'���ܜ�$����Ri3�Az���U;����v�m݃�o�z�\s�Ԍ���ô|�06��[`��Ge=�v���8J,Fq0��p(�5��b ��"{�Р,4��k��{����-���,��j���«rmXI��	͍�TjO�ǩ�\n��
�|
\��^@�UJJ�W>��;ˠR|[z����J�Aί���y��;��SZUg�܏/vxi��UtXm��Q��J ���˘�J�=�����LI�%0����s!j�rY�Ȝ����٢&v�*�3������-jR�j~�C�"�D�&a���3vgS*:O��l�-exTP4w�-�<DlJ�̖�5��
S�9+Y8���d�*錻Ke�"�>|�V_��5��]$�| d����1���C����k�S�y]����#�vk�8�g���*�U�F	���(c4d��$��*�d�_�!㇘�~�	���?q�PŮc>�9�8H��"|��+��	!��Qz8D0�`�ϴ=G7�B�ҡ�H������3�:1�������Iu�i���e�*�BQ�{47�r<���k�,�����L�H���������Al��NK�6���\1�!�N�a:D�D��.(��Z�n���vG�:��xԚ3t�}�s��zu�-��	8���$��i��V��\���O��c ���j�v@��؂q�S`M����Ƅ�iU���F��&ڼ���O�Ѣ�}�P/|~D��(�43{�A��3�F�ܖ����!��EYk���ۻB*�tt�X�:��̼F.�IP{�+��ƾD��X�Gٛm� �z_�8����\��9��@!��A�p��o<I] T��H��	Kr�����|-�5�p���yH�z�0�De���1l�Yﵮx�*z�Ƽ�98Y����LO��x��;/���x�*�]���Ա����Ռ-�����V@=C��>�b'��p@x?g��H�(?	�|�1��\#ı`�eB2w�D�p�.�"1�	�8�؍{��Ez���۔B)gt�aVF�����)���d6<@�P�T���YVoi�`Fm%�H��Z��;:�^;����nuj*� 4�i�R�y�uG��<�t�ĸ#i�]�O�n2y�£����3ة��C�F���#*|�.�ό\P`�G�~��B�?1���A�$ �9}��QT�����~2�専EQ��w��\*M���l�_�f;0c4����=Y\��4Ph7q!�4�@$������`��agi�u���%��(v�U�.%F�K��ҟ�I���c9��x�2�M�<�=����ϕ�//��Ǳ��b�J�w�e�2z�v]�>g�=6�|)�6	.<�_v���B$��u?
.1��ׯX|^ɖ+��0����F��=�FH�a뽕�C�����%��$���9a�d`���H�(`Fx'�ײ��f�3�i��-{��e����2?���p{"'.�Z�S>�lX��A�B����)�폞��W�Vw�d���W����f��}Fs���y����f��0d�[	���VT�cTor� ٩-�
�kF"9D���ו�@��s^TF�����l�r9ٺ�M^�{ .���eX�����6P>=������8��*�v�k[&�h���*��2Z��r�7��r_�q(�C�;	+=o{�r��%|Y�	rB���|�}��_7�RފX�D�h�u7떣��>9ūcٴB�%s�\��h2cu*�Ϻ�	>�Gul���71�^���5
�Z��9׼8��T��(��xPB�#��K�îg��R+���?Q���eCs���F���D�x4%%�4Q�c' s��T'ԯN�:B-W�P��^ 0�7e�JW��,����vS�F'K��[��s�/B���fِQM��=�YqA��_�_��Up�T�-��WYV���NɎ%~���Z�P���*GT[�Z?.�Gd�n��q򕝢�|1�y2{NY��y���%�'6��e6B9�мL`]K/�;l�;ǽ]����C���|a��!���*P����+BE��].>�ʤ�����{�64fQ�t��?t\���|����CR1B},'�4
k9� �]�bo�y?���	���*�Ty;�Xd��{id�3���b����@o	)� �D�%�cY�_7��i���}��SC�� 
�쾤#�0Ȥq-_ �X�U��+���D���*G��(�Q�6�����#�<������»��W��ם�G�XZ�D,1���%�X?�(?Lq�*�a����~��++YX��W��h�2���}erIo���O5
}Q�͕�H�:d��n
"O��"e�4|CX�W�9�e�!����!�PJNj�L�j5{�Gq��bsnEr���.VG*�v=x�U��,7>��Gx��b�0j��S��e�Gtw=g����8��4�$����q�	Z�h�K�,��2[t��!���Ļ�6)[60��G�͕@s����<��ςKM���7N����e��1�(�G��<�#~���--��ڨ_�\t�2�A�y��e�l��V)C�������3�}d�Yǎ��5��0+
�A����t��!l%L�,�
\
�{j%�IHϽ2� ⿒�s"��7�T2�8�J�e��O��!���X��z2�θ �G��
c��S��G�8�����ɱ������Z��ն��O2�� ��e��[�@�@!.X ��k����y�a��El+_)�>��HV�!j37gR�T�D4S�����y������U.f�f`�
x�|[;�Ѽ��ග�f' x�R]/�$�d�z�^|�� o }�B��:�h\� Au�}h�a��6�Q�-G�D^����?�<]vd��"�wb=� Ǌ8��$]cZ��N�������Xui2���8T�<�t���F�j:zT��e��֍����0�^��i&�~{���u���Y�0HYC��n���M������X�U��h�dڄ�d� W�|�)y��BՋ�%a��W)􀪅���L_C��)�nK��z��D�{����;�#9FzHg �������יr�m?X�k������A�!�%�&�K��0M���t+�2�������_�����!ǅ�y=��k�93@��׉�S _�#���_��8b��v��7�L�����MmO�Q/��	���5�N�#lކ�1��xu##�z�*a�rJ�2��Ϯ��N���|�UV3���ݣң�++�H�@���
��֤���1���@b&�QA�E4HX_���l䀠��<���4S�P�&}()���[_J��~����7A�)���'Z���r<��]�����O4ܱ傚v��y��{���^g��/*�%�K$���ۍ�#>}78=3���' �{��f恈1m�Xhm���Q���P�,��s?�bCr�Wf�a@�cL��#�
2��5��űah����ß�݁��8�2�j ���ZT�F��'�b�O7l���u�{�h����`�/ ���5
��MR3A9�!A�A6�N��!y���=y�����64���v9z���"bcV�������I��<_#��Q�p焤�׀�y�;���/}���Z� �x���aCk�q�O��9�K^DV�۴�698���5Qfz��|0��/�k��4\�6xv��c��Y˹I�T[�~C)T��]p����,f�b:��ƃ�K ��t����gha�SX��o_�<A>����ظTE��7��<D��O�z����񏠖آ'`�?A�(
���R�����+Kֆ�˗jC�x ��j�fѳk����<����w[���eq�6�w��X�%��N'�.��qg��zV�[��X���K���ßqk%�+u�fPp�S��_>�<܍�M<͕��MC"#U�y-�h�4#"��^��EV���GbcOE+`<t�<xk�e=L��L�"�-���8���h��ʴJ�kf���w�o!��h����.�w��DaE��=��/���>WV�q*˰��.��x��
1��CV�>���C�^Ő���Q��E/����ann
�d�Y\�`�Pҟ������&�P'��W=>_�K�o*��H�y���?��Z���up:^dB;:+�X�����/t^ ��V�s.F��Z�� ���	�$wk�+�pz�3j�`<Pe�mWXo>=�[If ��>l�JJ�;�&}������/�$�q7Όc�+�ʈL�iS��5��C3���[��ϧ���G��h_Z�ڡ�*��/;���	��`�w:M6Y�.$���l&e��C3-�C�Ti��;J�G�^j+��&�	�m�u��
�(�S{��c��:���X@��"8�9T�t��u���\���,�֣1�R�1�zq��$�%oSH�еB6q�t��8��5������q�벐��^ID�n}��ȧ�e]}�V�Q�>��d�e���0KDә/�k�!0TLY4�ů�-�F��i�����P��u.�u��V?���J��r��L)p�jz��rqN�m=�Wc3F	��A��ЃD���)خG�g<N��^��Z�uPu�O�����Aw��5b?�!�����tΞ#��C��T+�A�Y2,ej@z�+𶭂_����eJ��6���<�������lDx�3�$��:T#d;��*�-��[��IMܘs���J�~��P�gc�w� k�?f�(<r����͈9���9�Oh��s:���1ѿ�s4q��scY���$w���
2�Kv�%\��,� �kVҞaaI���7�8�bl�socp�S���;� F�m�9'�A�P�-0W@v�m�I�`R[�`\倻�m�n��_j����#���	�'t�����n�px���$[�b��	j�v�i�u�}O��G.4�몠���>~��b	w��[���FU*�:W�o�sRZ!�\ڸʒ�Ǐ7��G�4e�2��j�/���������\�m�kF]���d�0��y�\g�K�թ��O�{�B6�h=P���Nkiy#r�N�S�A��~��9��,X�Q	)źx��ޗ��\/ÅJ�FlƊ�ÅP��B]?�
P`ٽ�����%ǝ�w�p��M�d����V.���I �˶�ft�I�,h�I��<����5|;𑀕��1����f��cT���3�?�	�σN��k�#a��%�P}�­Df��[�'�,���:A�2�*%.��~���j�n����؜)~�~H�B�'�d�Mњ��G�Ajt_t!!}�e����2q&����Ȼ�k�2<��V���o�U{ޖA9�}�P��(�$���� �Gr+2�5Q	�E"����շY�tKr|�>��F�0q��3��95m*j�Ǭ�R��Q���2t���MJ���p�����W�����U�K,��̩��*�۫Q�	n"�V��RnK�=���7�#4E�,-<��t/P����q�_��:��/5Fzz,�e%'�IzSR��h�Fڋ��ҵ��iKLS��N���Ğkt.0}��o�Ǆ�� �7�{�I�����%]��^<i���`�9�^�Q�x8��n��y��1����ߐ|���:qd�}�aaR�p$��(���ȱ���*���g��k����s?�d�=��#��T~��47$9���!�yY��nB�0���W�ڙ�������h�������h��݆x@��WD6x�(56YX7�\���T����;J�jO9�773�"�k�B�'R1���A:�;0ݟ����.�\I�+۲�<$��c�����+���0\&�Ŀ�+��Km �JF�Q��u�3�#1���݇% o#R�X^U�p�~�5�W��.�Pg�����������2}����[2K��b�E9�#�V�ڽ���z@A.���灏x�y�(�K<��{�ט���$S�/�����wgEn��K�v�L�.���M���l[�����j�1����KG莆q6����k�S�{�[���D1=�t��l�s�!��0!�Tj{{�z��?jqA���X"t��	Ë�ݑUR�L��
6���/f��b'�d�+�'�nta0�K��T�;�K:�^]�����B���<�/��i��ѽ�T�Y�V�aJ��#�'^NC�bM;l�b)+v�>�PA ����eK\q��H��b�0-8�yTQR�u�{g�2�ߒ��\��KP`#�b�2���"��ǲt~P8cb�=L��̳��	7��Dw�S(��v�Y�ɽe��j�|sr���QN$׾��d�8";R��b�(�Z<#95J�]L}a>�njvn�I�-��K�[䔪ZV�- 5(m	�,%��R���u�6�A�y��I�x��KS2.�b�-\�O�;m_�&,��Q&�xC�>>Z�v�v�O�>-Y��7�\o^l��q�e4k�5�4'���I���I�
"�@��m�a;�`Jq�����*�i�;Q�~��
�W�� ��2�2���T��r�E�NfS�ǫe|�hC�?ķz!�J�[��\��)�\�a`����[u�Sz�ê�h��`*@���Åbj��|q �����1�?�"W�G��|����A�c�G�wo�[���:�h��J�}�Ds�Fn4��չ n���?���jVu�a��P�_s�'�Pĉ I�}c��&�O� ���δ�F:[S��3�Q�d���I��Q�!�h�Y���W���2�����%"^)	ؠa_�,X�Aj��˭�+�5�����	=B7V"��p,�<���~la���
�!\�|��b!��#�b�X�K��Gdm�lS2\��g��尦y�c1��xg�����Q�Mxv��q�<��ͤ�J}S���Ε�\B��HF*5�Std��V�|��F��#��:el��i(
^T�s��FUG�ad�*<;��B~��y>�~����^�x�㦥�H�3��Y��b�0ǹ?�:�G![Gn�J�ݑ�[��2�����ZeH��hq�V歧�gw3^��Q�����g�T��;z�|Mɞ��>h_�.��g�\�n���>r� Ou�]��KQ���ѵ���R�<�GR���K������p4n��Y�����v�.�j�`8�?o	�\E�������Z"���*�:Q�u^_�Ҙ����c�X�2KJ������p��,Fi1z�~7�J����9Q
�����8e��)�qfS�����~��ǰ2������,-|t=��"p�ڞإ���1��L���_��k���h�!�>�������O���j>WRΆT��$I��X�zp���Ƞ�\��=Z{�����~5����s�i/0πQ�'�H��Ov/��I�󶨾�r&)�'0& ���<W�����A5�F���kkdx�	YPC�� ��Y=UF^�h���^ r��M.�9,+�\�F2�l�*�nꉐ� ��{��QB��l�E) �L,��͘�N�{R�J"Y���#�ؗ�|;�����l��߲:7���	aȈ25w���v6�fB �iƖx�����BrR~nCO��c|���ErԜ���R &�v�}vETm.�p47d�G1���_FI��Qe8�v,�D:ƶ�GvUӛ�=�qp-��a=�����d�:O���>$]:5?�1^���Ls�6��뾨 ��TΦ[G0_�v�����cN�j�e�M)�D���ď�#;sS��'�ːe!g�Bm$c2��p�A�����wa5rI43T�rdT���Q)g�8�G�?}����mU����E�c%�k ՟��?/�6����!]i���#���-M��H���g�������zf����1`�訮� ��d�*Z��찔�H��b�aP�(VZa3Z�k��	ؔ�7�� �s:bg%�nD?s���{j�$�k��H����ձd)5S:Ţ�V6��`�,E<s+-�����#D������8��(g�����|�(�8�j��{[��?��E�ha2�Z�t��{bb�9��SL˶��c��e\�z�}���'�H r����U��էDkщa.FO721��բ��fL�]��c�b�=4��_��&��/<4��@�VQ�斣ٻk�u��P�y��>�zvR2��k�� ����z}�秭_{���Z���PN�6��6]HX�eX��-���]�H���#��@��<n����l/\B�;��@Ton$�@���8��"��1$�Ȇ�x@KR�z�6x@���FV-T܈�.��+B�\���Ȯ{8���Jر�'js�haw@�e��MF�|[�ǽj2�:�.`���ryZB�<���r�"���m=�Z����ّ�=d�3����}�~~�4�rZ�����N坜h���-��
:^�d2����e�}���QJ���u��  xT��(#1n�{��a��ĥ!4�O}D'��#I�\z�U/��h���:�§��%���N���l[~?�T�����`6�4y;�iw�k!� �)I�.�;լ�����W�h�8�)���m��7T2�'!:�Ӧ���Τ�Vo$��������z�f���&�_�;ه��E�L�k�k�yʎ6DđNGV�)�"��e�R�լv��B"�!���r�95X��x	�Sdf:�������]Lñ~X�}���E���D4�O�{WJ�����W~��炌A.�����5��m/���T�OD`�s�"�?Po(�����L+���D�KV�B�_���tW��#HwE1#g��8,!��CK1���y}�簼�P`�<�!���0��_�x�FÀفT0�C�8;�A�{6�e˝��N�˂6��!?v{l����4+�T5
T��D)ڜd! ހw����Y��P`?�'��v��P�r<wZ<�w�|[�be��kZ��ߛo�cqbu����șqF��f�ef��q|�,�f�X�l�[?��9�d2��\ƶ�AK�O�R̜u�e��n��������S�dg�.J�=o�(U��tF��m��&L�a�2�:����gX߾�A�j\%S�*	tZ ��-L�#6�� Ʉ3��J'�s+LG�*aчa4�2���:�W���h;���K���*��o�D0�1�DY���F�r$�)q�g�i9�U��Q4��{ErfP�&�N���]�C(�쇺��l��E�$D�.�#m����l��S����j8��EO/܇��͸�Ǹ�t�Q;�C��xT������ػ}�ǝ҆���N!��B�*�'��K��2�� �#��A͌$5M}GnYQ��E<��=9�v$����^�	���[ξ����
r���m���x�n3
���joe�9&��g	׫\P�$+���xH>��Dam�f�z!���C%������5 U
��7�M+��@K�<A�_�b)����:�d�l��[&������?}��HCy�͝{KCY���yE�>U_k��REЭyn���՘��d�"r������v��^�Y\8�Y�N�N��ke�����ģ�$���g�}��K���ٓ�o��Q�v��g*��{�*�
"��>�+����u��>0k���|��N5��!P�?)��Lg�s�{JM�&��d�i���#�\u�'��a�! ��N���Ø����#5T
�]a�~X�h����Y�]�,���A��^q�{�:�^�qD๣�V<�U1�����jP�$����u#G,t��Q�gwc{���X6�
<��R�wt<gs��m�m��8����.A� ���^��F���׸��.@�n��-bD���(�暁�mYP\?3�u�F�E�J�;{�?�]�Djv�֠��jpF����~<tc1W��1$�����.���`P��`2��*�jV_�Iu:�}h<����9[<u�e��f�F�)�zgHb�X;�XoaI[Ɖ�t[��p�˓���p�<��K�3U��X�� ���!�F����ǈ&�{�\�q��4�����8b"���V�tԅpx��֠"9E#ꑰg����� P��B�Vn֍�����I-��S��/���~��� �C���m�?�Ϣ���6�9�4�w�:%M���;}s����/��������3�Q��������B�}�XTW��0ۈ�T[���� �||o�@��J���h�g\��m������3if���|���.Xě�UY,E�]ҏ��D1]�=zp
����I���^Z'�:1�K��T2w?�Yo����9b���2��G�ڼ <�ݾ��XL�
�LZ�Mu�&T�$�)�q�?kU=��1I���Lݘk�8Z��o�	��N�������Yg��ֲ�&NI5�-�
%ps?9ŀ�|o�Zxθ�+�������y#UW��EI��D� �w�x��0�b�j=a0Gym�ͦ��?mT4M'�!F*��X�t��E��;�i�%�Y��;h�[Ē�]؏��t�vk�:��s��ʩ����p��ӡ��C�3r����"/�x,�}c(
m��xT�7]����]�ĭQ �/bXJ�`�S�$�@����40e�^�8�g�h���
FRP�� !歓ܗ2��&���d�S��(2pcKr,�{����@��`�lYt�����V�[����v.8�
�E�t���-��N &P
�|�
3�jj����!<E<���dJ!UZh*@��l�u[ ��)�M��T1��x���_�q	̩�Bn��+t��/����5�W��gM�X���qIG�Q(�<C"���h0t#�����0����n�u����"���ZD����iBmH����-��t}�/�-oI�d8^�j1ȓ���^��p�â7�e�S�K%'�a��'�`L`�L����&��]X�q	��zE��E�:��Y��� ���{�f���˪d�����H���ͭ����ƞ�1<8��)��>�(,;����Wɍ�K�ߟwl�����޿��<H�{~^KN+M�.�Z�rK� S�j���5A��L�F�ˋ�V��� �!$�E�����Q�$ ���(W
��8A����5w�ê���=�caM�����J(����'׳���X�D_vfG�Y	�~S</�� �3f��P�S����g�{w����?1o��ϋ{D�C�*���5�A@N��}���g/�dg�7�Ԯ��i�G
	O�s�/�O:�!�o��:�&����@�qI53��id�J)�S�����7B2�[�<�Zc�f�]��Bf:u^� �~�Q��������:���~衚E�?��Y���0�D��WO�h���A�7L���?��Y�~OԵ$�閱	��u����ښmB?��Di�=�V]1ZSok�R��w��P��Z@9�򍢥���]�}![z)�!-�ۧ��$y�h��<"�����p]�;��h��1�,aL�s	o1����x�J����ԗ����~��5*L*㹎���|7��!5�ȣ�}5�����m'���ouXl��,����Z�A��y�ф�i8�>�V�+�/�[�fX��w�t&;
�/ɕ���'m��Rr�cA�0:T2���P���	A$#Ya��I8��q��os��͝a�M��(� g)�H��V�b{769ɐ�9�N]7@����G���ë�g��!��0^H�wF��/-�j��a��[���̊��4P�4�ز�Jf��)�a��z���X@���^Ug��`�v���jMf�֠d�-��\{~�d0ܔ�>Ӭ�R�Ki>����ٓ��1>�!�IwC�u�݊��AgP��'�tM�"�!g�_G�H/�,D��7}�[4<�����@�7b>c���$o���3D8d�:���e�c
�z�=��F����'��Q;h�0,&�\�a��%}g�(��E�1n?�^}��O�1#N1��-h��OU-��R����I��/<����u>Փ����?Ԧ�B�3w��I#�O��ح
����
���l3Yג��Yx3��آ�<�תd}
3"����$1LDD����0|GF���(N�����A��2�����~u6����A�B��	������s��8�;a��ݬ�^�؃�@�繜|
p�p��Ӧ;2�ڴ�R^`�_�=2mS!
����������\m�9(�3�����Wډ[딚Kj��.��;t~��ڞq&�xFM� ���5�$|
ag�~Ǥ�ދ�<@-��-�����T�ߋk���"m�Ju�U�7:IZr/7��}��k?2CV�(��7�;�%�1���Q���m��(�������M��t1s����e��Y����~����9�9|=^'���RWjٔ����S0����*�L�zk��� r�}F'=���}.ʋ_M���8P;�B��-�Y�?�rf�B쑥� �!�����"����R��!����V�������w| i{�y���2J�n	>�;
r�;9���/�qk��gK��F�Q�=(Ɖ�pL5q���h?�5���O���oR��M���c� $���`O^����5CW���Y�s
Ac-�)���
�*��F���f�����S0�'yK��,�����fa���G�<��1���a�����J�_c3+��Un���Dv__tO���I"#�]���б2��u��\%;�ŉ�\ň��q~09��:�2�Gi�&� �U$mT��(��)��k\J�� �aX�խǜ�k��a1��$�ԑ�̴� !�Ɍ�`V��`��J����<,��n5��f�s,�:�sT���{�ڡ�Y:q�! 8���&N�	�r'�?��R���(��q���K��?o����^,�Xi��p���/N*��	���ڞ�C͑J�&�U��V8T��G8��v�c_�������'����}{��Z^�H�ExblC���k���R	(�E�}�h��e["��Y��ֲ�����Q/�<.�s����}m�Nܜ�p�Kl�;
�F��#��x��E��/M!�I�����f<�B��t�5��zp���o�ns�arl'՜)K�>�����Y�{�g���?�ψ��|?�(�p!������ٵ���L�H��5=��%ntz�ySH'�����ًk��$3�^H�+.t��ڣ�[��ܗ"`�e���i�C�"�ӗ�<t��O��?�=���+X�Q}΂~�&,Q���|�̬܂-��b��/z�g��Wz�ޟ��� Ow�v�ש�ݜO��4�#�q"XI(A⵸�^[��Q�1Nb�T���t�p``�U��Q��o����*[?$���P����nҤ� ~K�J0��R�c�gypF��&'3�~s �˺���U�!���D�/�^̲T�6�{#%�wzbޒ�2_�b�܌�W�[,���OSxק9��J�Vs�����6(��$*^��ņ����ש�G#a�p�'A��2����5��� ��-n/LbZ?���&+�:�P���q.�f#q|5>�.D.WP�D3q��;����A��T�}���DJ:՘�`ޕÖ���z�i�V��=�-�0n�����A�t���H���`
��d���6����K�#�ђ�P�f1�M��,�3+��Cf<���������`n	g���I���'H�,=��X
������a�'@z�MTB�@C_�U��爊���Vr{��>Ҟ$U,��})rE�9�0��K'�ކi�QJu����I�42n�r	XrvNV{u8�ц=��Y�H�4�o�y��q�q�Zi*��F�f��Փ���'�ǳ�Sb�R�Ș���|��=��{�g��c��܌��d���"�<�sL��L�j��G��3�[�h�_@��L��no�űހ�?�����e��������ń�@_�p��J��i!�_���u�(@+�q��|F�-��:s�����fi��G�g��Į��ՀGӢ��q� ܾԦ�d��7��Y���:޾Y#���s����L��hҔm��^\ �vuR7}��i���:w{t�]��m�D#�/d(�h5�3���!������"4s�4�)��63��bY�ۊ�J_���;Z�tpP�t�2����a�2�/�
3���>�3ۿ� %ao
�r����\3zBV���Y%=��A�t�?2���4�mX�Պv��Qy_�����5���6S|��)��7�1�3�X'������� �p^w���r�o�����-X����w��D���6ǊJ�4H�zJ����f�c\_�6��꓁�1,�E���ҏ��n�̔t׾�_V�%v�,����[��q<��}������m�%2��c4}�߇)@kd�Z��fx��.����w6�	���s�4�őy�k��	���%۰`� �����et��
B{��Y��[>/��q��(p�m$��ډZ*��8,
X�~�|BSx���;���p��X�Y�;��a��<��YV_)13/��9ا�1�\����ԝ�L���7�t;�2❉k��K$f#���(xN����]�<�U�e)0����8y���*j�B"��i~�ֹ��KrS^�gȅC�[O������������*��#��'�xJ1�`��N	3e�Z��G2["���S�d�.�Z�5M#/�m*���n>�fAn�Ý��&8�@"�\^>�'A�����İ�h�@J�H���N�?F�����9f�e��-���xv�yd�V����dc�&�طU@ӆ��"q�R��ַ[Bd�X���~͞��Nn
�4Ю�7���s�%D��o�l�/u)\8�J�(<���#�M����Ƒ���'\�wj�]@�#�#�(�|�IT"�s������d�r�grͬk�x-kp�m$_܋�0�Ϸ�G��S���yH[�
`��!PqH����h�֧��H��8e��+��X�`��RR�����k�|���(��@ '��2sz��*�g��<��7&���Gê/.8�4�o�K����� �i#��2���a��krS���|M9��}���H�a!��:��w~�d��>���K�m���2Xp�p"�T:���WK��֗؉�����!�R��O�.�Qt(`S�Gb#�g��`L���H	A�r�S^N}!�-��E҂����f�wH���:&V��D�,�5� �n4p�4"����A�W˖��Q��
S�x���1����9��ec�x�'��F3ewxֳ����"���OG�z�q�nF��������*�n�ؠ���Qܦ�-���?�X�@���D@��1
	�˅��9�e4�)B�+�a��jX�����>��z�����7�d^	0�,�u�C�y[���J�>)�b���o$Ԓ2����ֽ
�Ao�ϳ��#��GC�Elac�Pm,���K�M�g] �39w�0�	������ݵ��-�`:3L�y��\``ӏ��|e�)31�v�m$��e�re}�k_DXx���Ǔc!�B���U�H������¯�u������/Q1ࣈ���t�e�a4[�����N��%��;H��g1+�[Ú��|"
U�x��^�w؊z�sJ�M�;���Mr�!�g�s����`��[�����4��G�aR^se�$�7�}����\B�+�̤���%'�Jvv��I��}Ip�*Y�H�@�<v��h@��6�����l�R��1�#!�A³m��ZwT!C��L5]�ޤ\��G&#
a%��Y�"�ok�Bk���������� �?��gdާ����B�d��}2@q����۵�Q�@ʾ(��ԫ�dS!]�8)�9xy��:�YxO̰kT_*'w�˥X�Ku�"�#�BKA�K�|ll8� M��v�#.��V:#/���NcV�pȡ)��m��������[�S��ѽ�(�&�W3T3���|̇8r�ڢ;�*!�r���y���_���a>��c*�I\~���q�5�yϳb���*���\�>Y`^�����s�5|�M2R�b4�F��\|�i~r]~�ȰtB�{�tb����x�2�|!\�"I��ۅj��C��[6���g2.8��i�I^���C���� ��}#hTleR
��U���o}TMT���e~#é���й���+}�;��� ��Ԫi���k1�����-6�a{dz@p��H!�}.� q��ґ���rM�c"�/��v���yG�C�����yt��>ҪL���#I+�å%��~s�-m����~y�˜A�cWb���<N�Uv����NN, ����21.��Tp�.e����P'��@;w�G�=5��:Q$�E5q�Au�:����l�Vh!�~ �#4�b�l����j��[X��}"ڲ�[6�@^|\j+�t����*�����LZ�ǳ[a���n$����G�`�+ �5��WV>��cpT�@�n�z4	3��q9�6�%�hY��N�g����� &�ҥ!��6	z.�-w�&�x�:���� �)+���d[��y��M��H��������1.���"��[��˫��{��w/=�:'�gN��� D;�F�IRvF�q�H�r� ���U�i[�a������P��,��.�[�SR�Xr�=��HٖkR�o�m���נ{���Z�w�lP�vH�$.��wz��D"����KD��N_�dN���$���J����}����-%9DV[���Z����Tמi,	^����2�?�%|�F���}��{AVH��~)�2�J��	����C#L��W����ng�q�n�A"��8$Q?��,rԹ1�Ǹ~�$^�M;wy8�pB����M���j����D�5"�'ߧ''&9ޞ�.� D(f�%4̕�`�O@�h�i�U��=Ԙ� c��2P�3�\�?*��S8�濳rD/Y�u�)<�	P�2����p��][���*31����s+��	�����P����l[Xd�K��Ա�R�oi$�뚸}NAӽ}���'W'��Fu�ެ�7ާ�m�\��ƴh����xX�C�pr�G§>(�����lS��	��C?K�'����ږG�摐��-��� ���&�ݾ��%�8[S�&�v�a�BdҿI��f��%HUw}��sm^�L������\.�����y�C ؏�̛��I>	�����w[�ǻ`��������>�#9�TB�A�.�N>y6	���M�+j��kˎ&��!/"�4�vf�H��{v��؅t��U^�?�Vl밪v_�%|?Д_����>�|10���4*"�1�PB��B;U�sS�/%0���lxҨ�t�F���^.����NM���_�$�xqU��/�,R
.����%��t�62�1�oV�|���F�ɗ����\���7��2ڶHK�������h�Ц9 C�%^�)	�Z�s�Û�����5Sx7���<��dY9mi[�>�U���]�z���r�ʘz�O4x�6���-?��ؓD�(����9�-�F����ݩb퐈TcN�]�&��xz_�{�Ħ����PNg۱\�����w�����?��1��'Gl*$�_�La|�Do�ю�\g�AKء��~���c^]8��sI��˻���Q2�J�1O!����A���c�̑��t�����"���(��]�E�wF?�����7^5�`FT6���M��KJƞtq�<�MdX*�F�'�8kX�zD�{2D�'�3��w\S����i`�R'"5�Ś9�����!��ރ���#z5�rr�%gdP:g[?}�p�� ��-�FF�ҿA��<&~^�f�4X�_����û�.�z/k���oZL>L����Y�����g����e�o�-�G.Zt�a""���o��
�[�/7�����6�d>d��=�ޒ78�9�_��H��s���u��g����Դ �x�K2>�(Gr�3r�X���:�Fw�{��e�I���A��L} �ͺ<^�H��7�8K�^��B����.G~6�1���!��pנ/��O2y�(�2 ^�H���= A)� �w���I@E�Yb�˻�D	w�,�]�1��S{r�����-����r�p����O�� N���o=	=��[�Qw�Q���r�{�ضR|���TA����E<��K��ٜI$�*L�ȃ���6��aU�3yB2�C61��m��̬�x
r��!��;��������t�"Cj�N�Gh%����wv�b[���9���`����+�I�A���-{0Ti���%���;�9R��-����]�1��P�SLi�W��@�C��F�p@�u	�jo��A
4޺`�s���Kw I�,J��!Ȟ��?��*��%P�b�8���$Zqe��jF�b���c{ɡ�K�^���C���a(އ1�ì`;H"&(�3��I��R�HH���9�d�P�ͤ>?/�*Gҙ8��f�����7�%�Y��X��$��o9Ke�ڎ!��L�+TF/���'z<؉A��W	�d٠Ik�.��m@�(�Z�Up���N��txi�b~V�]5��đ�t�G���br��9���h�2�5�(�%f^+ǽt�I.�g��CJ�V�+��T�UG68����J�;�c�W�;P�Bpq0�dxlC�P�^��-��]����/��~h�4�(u ����jv�:U�;f�mk���k=�=��-<䒝�sU�l�ƫW)��G2�63�(ǎ��<\�mUEF�g[���	��
��ř����d�kĥf��z!` CW���8	�A	J���AMKD����-��>aÂ�ް����4
���ߨ P����FR��4�OK�@h�G4�Ƨk[�[Π��5,}b�$��=)\YU����3�go��'��������/+��{	�{wt�F$d{5[�]���Y{.:,.���I�r�*r+?YT��e�7���0l��9�u+J��q�j#\�ҫXī*},�T&���R<M��:G��]Z�}%�B1��&� ����e�Y�����c��t<���撆���+g{�c�`ARƤ�&f�$����w}x����}�C� ���3����ԍ
��YeZ�rY����؀.-��͒éϝ6�s��`z�������!���I�eZ��ctV�f(�m9CF����T;�d����R9�5f��}���e)un��?�i$	��h��E��	��硄��8�"\(O#�	q��c��������)��&��2�hS�W�oX����H(�a�����Uh[��/5�=��hI���c��T���r9��1S'6��'�ox^%�C�Fn���H4#�8�$-�y\M��\��A!���$b	���[�~Q	��-�o��G�i�4\��H����N��2����Qg�=�I�
�x�'s���P�]�e>���,����UQ��$-~!;we��6��5���)E���	�-����u�@�߃��X���lWK�E˳0���lW�n��ַ��C��Q��0g/N�������=}�,*M��/�E�;�M)��^��N���������ӹ"��H薉��(�K~��BG� ���e�Pa{d-n�	T�L#�)?o(v�O��0�u�a(��-�r,��fQ�=��oo^E~���u1C�HJD;���lT�.�v�HV��������
����0�b�x�.�Ӷh��R�;�4����G�����0���_V�0
�O-bi<E_�_5���z�>r䀇�A���(~}�g�oBd3��-��&%{���U��jƞ�-s���J�Y�M�ó4o�2�9%�ָ鵄�䙒E�V)��r���aɀ4�A�A�j�RX̽�o:�����1Y>fq��*da��&���~�,cT��M���!a�|�S�~Ac��9�F��l
d��+���V�/�W�B��v{�X��,�ʂ�����.��[W�Ը�fx��C��4��E��Q�Z=��Z�RQ�M�'G�b��&Q�޻��,h2����Ԋ��ȷ�Y���-�CrnC1w� p�)���8���Y�)_��*���)q~�T����N|Გ��:�I�Y���O��խ�� �7B~�$�_ֈ�����u�n�CWP���q�4�wr�ڷ������K<�������k�A�v4�l�$����q���Fy��L��+�K1�N�(8
t5O����&os���CcL���Ig�cW���L��/�4���s(�H� ����V�r����nQ]�
 �M-���;��6�i�Y��ZM��4%5my��|R_������^����,LP�n,>�r����=]��~e;6�n��pڋ�*��C��q��h��$���.�l��8I++�)��$Q��W��%��lEFW����*�	��2��>�r�&��1ޥx�DWG�H���$r�݇׃+�Y��f�[��_�6)����D�<2rө��I�����-m�a���b�_���&?��k��^(��.ۺ}X8�.�	ܩ���l�KYD�9:�A��������푺�7�)f_8�I�����ir���uݶ�PR��_Sf������:��<�2iش��e}~���~����M���
sf���ܦ����<�GY�צnŻ$��0�6��ƏX3��]���r=6R+����$R"Տ�m�ݛNY�^�f�r�f�8D�����֖����r=���-]F�J���Q���ΐ�Z�r�V�~N�vrsE�,R��*�|�Ȭ�ߝ}C$97и�����`�����	�9��!�ps��y���;���}!�x �=W�-�Veq��F19�CZs��%�f�;N��><�A��2�سߎ:�M��,R���}#8ɢGF�&��L�-�;��ZRÃ� �G��$C��:����vW���)u��b������F,�`��ͽ���\Lb�H�=w���~,ejpz�UO�OL�uK�ẝw��mE5�L����E���cA�/pSN0L�j�R��w���UV7I�C�f8U�ѝz~�JZ��^{ �v����d�Q�H}�0�� �)2p.���{x�
Ey]�j��>g��^bRO~�폭x�~O]ͫ�#G�ل<R�����us�Pk�}���wOXĨU��WZ�w���L�\�8�L�Ng���=��X�������'�v������������WE<c"A�Tz�'����r�.����?����+��l�q����]�y�ڕ��(�ڴ�A��p�}�ΟOX�v��E:�[l7��vq�Q�O�v�������!� ��P5��g>`�]h~��9�����_����3���+��Y��0�c�Y[�3|�ё�uzh
@�AB5�8���ƞ�|��J�2&���j���\W�f����PY�>�gn�<��w��-��?Z�Y�!}}���#�޾�/��׼Y�n��l�ǁl� ��������~pt>��� ڮ�Z���=�:Zj��'U��|���;=M�SK|�6���L��=�{e(�zSn�9DleW����up�<�.w�����E{�'m��'�!?��v���xT����	3d�q_!y�f(��$�2k!�y7���;��|�̚Xh�C:6&����d���E����ד�>�_��x�P���Uv�
�DOV�2I[R��I|wN*�>3K�n��0A{��,L]Iy��0W�zR���ޘ��O�D���Čmn.ʎ{��?�94�ĩP�m^Ջؤ+I?��x�.�C�ڿ�3�z�55��e=
�#�H-�RBn����4޸ lJ�)���e_���(�QٓoyT�bj��b.Ӊ;�Ԍ�`�B|�u||"Ռ��|,�t[�0��R�\��v�jU~ʐW9t䛵b�A� :Fqr�Y�t��/-���܆{>�"����X��q�!����E_��,�<���n� �����x	>t�����o)�,��݉F�Ō.���#e��YD��C	L�c?ȩ�����7V�^N�^~��ݭ���@��g���4����7a��UhE\��¿�9�'�����kH�B�G^�ֱ��;������Y2}�SY?H(Ц@����Y6�Q0MŗV�9�k,kZ�嫊*��
-j,�kP�D���dTY0���=�%"'����s^'ҙ�
«�`$&�q��Oo��b\�K���Ut�r�8���e|P�t�djBNŘ�q�@��J"$�ȁDz�ou�p�>�����EZ�t'�CS��ɫ�6`7�u�D�/�h8.،ӈȶ�>�h�h�JmZ��Z�FD�oQ�E�oM�es8����5Y����#?K�؈(⟬l��+*�+K��O�Xz�I�L !4����I�PE6nfV�P�᧛í��i���҉)"a��$�H�@�.�M��`j�4�V�dG��*�a%�gl
��@�[ b����<%���4>T�����	L��s��J�8��D�,�������a4���߸�$�5O[�ί������'-�x��G�K$���Ϸ��]�]����l�)���D����[.�1���n�p"�H�������	�4'����c&�m�<���)��w�v��M���*�
!`2h.f$ ��*��	�V$��:��5�C\ʃ��W)`N@&вw��ۂ���a����U�B�h
}e���٤B�ԙ	t�]V�K�m<f%�H���T�'4�+�v�!��9��ߩ_ιO��*�+�R�D7(���f���B�>a�C�1/�;'6Ú��vm�v08�
�6����>�u�|����f��-�*��}�~���!H��>� ���Vܬ���Vսe͐�k@������z�8Z���#./����Ck���i<`�3�j�mO~�������;%ƨ�]}�I_x�K�
͎��~1���瀃���j��G:�d�b�Ƚp��V�,|��sǆ������TnDd�`]�N[@&A��w�J�� n���]���-駽_���hJȸĴʥu4(㦉>�@�V���ٳY}�:u�aCʣ�����𵬷���6V�'<�M(z��q9�'��W�T#�ņ��I����mm��FEjf6���nA�HZ��������Kֳ~{g;,�M*��M�-2����C�=����ݸ�?J����
���F��xF�)��ۧ�kW �h�H��N!��#X)������sFQ�2ѕ�\MY-Xp>��9B�P��	��-w"�X�x~�]@zhD���E�\Fa:���8%y�	��L�"Dy�����&	$d����=�F?����p����PsP�*���,s�?�l��C���F�R��46���`�T��~����p��x��i=��	R��N!R�CO�#�F���
�����W��?#<�����ڔh��N�<�����p�����s\lo�kk�J��%�	Z���VX9��_2ԻZU�]o��e��_�y�Z&���Y ���lИ���4@��V��aRY���2���2���BȌ��s���~�5��klk�ԀD��:�4�sê}��@�����9�qo�E��K`D�M �B.Ґ�h���<���uf��I�l;>l��u���Ǻ��_A	�=�/����?B���0B���)r)O�\RJfY��p�"�D��{h�3��R��Lt�O���������O��"���a��O��b��
\<�w��O,��s�\��'/�� faU�n�K-����ج-�n�{2[1,�7����*�<<RG�i���sWWÎ���'�<����ד��.N�>Y��.�IN8���aRo��$F��S��� ]k�e\��Z��,L��8%�q%��nX}���8\�M��PLiӪ��N���N��LN���t(Ӎ�ʑV{)c8��%)߰�#��g���%����ز�|\�AUTU�~T� \�=�^.��X�6��qֳc���_+0���k��uj,MZh�L�-��.huG���.2Ji7����ћ�p�h�����5��?f�f1�7�߳��@��t�{[Y����T�K^5_�&,4÷0�kX >�/�qo�pQ��E2���D�/v�f�+s`t��X� ��z�,a��.��
��-a�,̀�oZr6N�sӜ�w�}.���-Z8Y��"�HH���?�.\�Z�/v��;��H=3oP'"�H����0��G^y�����>������U%IÊ���e�F!���O���	�K�5���5������*�j��@&l�A���`���ꨞ����P@\�6�'��[�}ȣ�����P��V�/�W��|����g��jö4,H-�O�]��&=����a�:Pp,<@Y��&;��E�#�?$���&4�5N8l"f�K6wdT�We #,��.���w@p��k����MҾ [�*���2����?|��b5�:�,ц<�*lj����#�Y�9q�1����Ň���"�;G�۟�R�O�0���,{�~"�&;mc�ӖuN<!�� �>�@a������آ��6�6#'�]�a�R���[.ˈ��	Atvs^4�c ��g>��í4;s����7��Ni��8�jȒ%����BK�΍΅.Zh̚h�%j�Ee���'
�=yX�uR
9z&��rr��&dZEܔ$x�*�#L��񵘢K[a'��*�+���U*�8-���M��+m&=4�D���L����������t鰘�xt��M�8CP�SCG*S=ܗFX��*_ֽkNu�9��j}L�Y&.�׎,��KM��+����1���9�0��q�Q�~��V�4�lxkPNЄ&z��$G?�ߎ���'z�a�>�Tr�9��,��:]�Vl��F��\�����Q�z�bu���ԯ�.�$���B���V��V�n-�΅:خ��A�n�G�ݾ�]M�S����T��d��3!$s�����ֲd�s������uǬ����<�f�{�&����W��}�SR�U�>��,��Q{���o����0N��N۟�gU��Q'�#�=�o�k�_��u�e"�3 ˧[@��bzk�,�,>�1�a.��<(rx���ٗx?g\ �[3��+u���$ML�����;�1�DW�x�����k��lg��h��n�*W���J�R��̆�����=���_�b��PlO��U�"G�/�Cd�w�6_�j�pX6]@�ÿ�4��44��񗂺���e��������������ת*䤂���k�x\�#w6d0<;E�r�?����׷H�Ω��l�N�x�=D�"���UHt��V�F�-S�����hp���Czb4^��v�YdD%�S|�+["�h�]��N�u�C�bЦb"r������'_E��eo��:M�&g��WHŬ�]+k|
�HmO�bf6��L���K� kO��K(bg��{��l�7K.Us��T�d&}&%���p*���.a�x?�q��h��]C\V$&Z�xL�| ���j���V΄/�Ct��%a/��(d��:7E�Σ,�%l(���h��j���n�1�A�����$8���փw����p����c�?��H=X��qP+X=���K�� %��A�Ms{[�\��@(A������n�/�]S*������5���=ǡ���5y+�K�
����|���߉	�h����  �rk��Wð�֋�/S][���������"o�2�"<ԏϝD�v�ў7L��>դ�=���`v+H�L�.�n"���������9�E���J6iY=\֢���wW��i-�\���E ��3ed*�WG�@�nWj5r-�ױp*x�S�+& �p"���χ��=�Y�B����k\:s��}�8�2����Jf����E��.&�y@�	���1��s,��A#ed�+4yn�+����8�K:�YG'�'�н)�-���[�������K ��c����)��{4�HD6�VY�|����6�r�D���?�y)��A7�˙E<1�Ͱ#Y�l��`oݚF��W�5ex� qa�Kjl�\��X���'7=9W$���033�n;��&�]��COsG�����_O t X>�������MTЇ2Ɍ��G�����ԩY&G�A�j*�7:���lj���'�������|z�� Z�!Q���̡��Vp�`'3d7C�#�E�'vn%@s3tP#v0��#�t5 ��3�(��!�Vw�(�[�]`� ���"*��`�Q�f��Bmnn�sp��� v��*hT�r��1~�g��o����
7���]C
x���j�'���NN������)�wl���`�)���}l�W��g��5$	kBp@�����I��������S��n�}��
�琞4>�ٴ���N}&4��%o�z/�2��n(=S=1mH���6[���+�3�e�/���)�72�Ҏexk���f�X������).}oW�o-F�$?�h���]���ţ���W�3I]?N�7w���2�n����B�.X%v�Y8�#��pC��>R�#�����t���ۭU�B�>�PBF�M;��ậ�g���-k*8�U3  ������h���0�S�T:79ޞ�Ƥr��K�j�~��7�f��e���ԙ��} v�	M�E͇T��V�g�4�z\�ao7��d<�n8v$@*�N�p�v��ۘڞyU�����%�Y��$���vgK� s
�U��#�	���x��ͤN��/��l��W"鳈�*!�
`�{~T��5^to?�f���n�΁�,s�4�h[��*5�
���Bk�V<s�,��]���	��#=�����-N�NŞ�ǧ.t]�p^zoĳ���cNLC���n�^����p�W��9��T�$���!j�O��0��~!�˷D2޶�l�1Cw,��'E`U�v2i5'oM��;�����")f��a�6GYE�����|f�+�j!��撉Z� Չ@R{�RalJ�du��,���Ele7}4">�i��ޥ˗�`�-�-�X����Y�@CLq�c-��y��Qр6��	Y���Iq��YUna~�%�a�)�Ǟg::ң�"/�3�7�?FC�5�#j��J�{w�6�H�a��v�.2n��T�BG^'aԗ�)-�A{��M��EB��Ԧ��w�W�2��~�-�@�}�� �>.�:7�a�ߦ�o�5Vv�h�,H��w��t.���
�j���<�� �;�iC3�c3zlD4"��Һ6�W����%o�q)҅�	�7欯�찵n��I_-?��Y�8�#�z����[3:Y�A�t�H����*ɻe��ͫ]C?�g��CF/'h��������,�'���=ؐq��T���ŏ�N9��Ҩ�U֔lE�Cti;${&>��j���`җ4�R|�$,N�i>�?��(��_��D\�(Ù������3��>��+I ��[�� +,Cѽ�Ds|cYa?U���:N@
Ib"*�Ay��$1��E� ���y{X1̤u"[V�C����e�?@�z�Lg��X�"���iv����^/X��ANK�񼭜<iC� ּ}�{�{Ȭ���w�G��kei��9%kS���]m�~g��^%�'��T<R?��bG��fA������1�>"��>B�j��T��u"����Ӌ^u��my8��$7mj.I\=�����=Ȭ�mv�
���.f�#�6&] 4)kk�� �����s���NXUN��h~T%��	�u#1�[��CJ�� ����!��\�q"a���p&�5�J�hū��6K���4/�@z�K6O9��Y�	��B䢝$�~d���>8/�.{��wN�<9B���rioʺ�b<
L����.�f�t'�Ʃ���!�)�i����z������gkq^P �5�n�\��d0�m�G[$K�����'�x�dU�8	�J�������]6ڇPɳ��Z����b.c�g�#���8
�����a>�I�h�Xw���I,�B�#��qG��U�\�����;x�3,�5���xL,7�a[O��J$�V�!�2���@��GIOuìnL1�o����9��BLMe�b� ׉���;u *�CGw���1�ոnT%MW��5L1���� ���������An��m 7V��V�L��3y�[�`wr�0ݳ�A�z� �Ei�#��Q-?|��l�&�\�Rx����/r��.ý/�q�B�M�H�F�Ej;r����r��+��cҪ��?�ׄ-n��6k����Z�B ?r\J
�t� �x:˄�n��K[X��hE{��d�z]�) �V���56���υ�uۭ�Fl��!��ۏ*��;*H�8 ��u��׌j�^Ԙ��=�r���{y��alD�1��è���rK2t7"�T��;��-�R��m=���SB.�y���BO�~�JEg��@����h(��ߓ-"�a[�T�M�~İ|�U#a���M��d����j,��W�Ձ����g�G{�v|�0�2q����D����T��\����@Ff$�Ү�|�be��ۇ��R�>$���tZQ�1|��Pt�n.�\��x����s���PL��ݧ�=�r�ɡ�����EC'��}���!�3pĸ�"���!P\�B}lz�u;K�y������u��E]���˽²��Q���jbD�y�S.Q �7CMe�ʈ�N�����ns������0��?�$o��R��<[o��LG.�b���EX?��}�����m.��+����)Τ`�{�YF2<#�����ŏ(;$�2�	:|l���޴����W����^uC�b]:�B�ɵ�2�X�R��XzEJ�6�B ���!�n=̗������"��ǈh��fmgo��7� �-�]��v3�\:�g�	>͂��U�栃�d���i�*&��Ht�>�L�np�T�AD�x�����I�؟�Օ����k8ǵ�E$�p���gJB}�Q5gM$��ے��i���A�ƹP#�rMU#q0i��<!1*4J�αMG6��-_{y_��q�OxK������h8lok�F�}z�yp�W���ȉK
��G&�_����(�v1˔���(��	\;n�~[
ޛ���r��G�:�j�*[�V�+��K�4��\���MZ���-(:�/q"XO�f��nw��1�=Y�qQ$�?q+�^ ݘ31���T���Y�e�W��!�9=D+�Z� Ppt�v�Ş��O<�[�Й-Bl*[R��]Gg���&�����0�D8ܱ*��ُ�P=%�����N��_8?Y�hi����0�fʍ��?:�kQ$!�Q��9�l�lP�.�Z�����?iU)2�
� N�pښI��)^=�ĝ�:�*��K����ѥ95�v~4��� d�����џ%,��/%��j>�p��2?]� ��j��������3�:<q7��u}<=�g1G}��ʏ߳�4����e��&	.�Q������ ��kٴ2�4�	rA�P�p�3D����s�e1rY�A���m�\�V;���Na����x�CP[����ЈFz}�s�\��4���f�T�.�������<*�Bj�� �(���[�R���_oҲ���g4�@^��y9�x݋a������eU����m5Jq��k��C؅�U���T�fo+�I�[s8$$Ը}J�Oxx����}Ć��K��E��U�3]�Ӷ�B�ր��Ç����)��a�Ӹ/ˇXl�S-�v>^�Q^�R�$ZRC�r=�!��{��s�=M���dI�.]�����������z�#����Äl0Ul��F�;o��M<�:1V"\"7H8O$d������~c�afZ&N7F�F�F����[�� ����\�c˅�� ��gO�-�E����[��G�ҹ+�"˥6c ���6KR�`��ldr�)C�Xm�E�����>�?7�=�CZ�(�i;��X��زϺ܃=Q�	E�4R��H�it�ᴈ&.���-�˿��|�#���A�k1k�I$d�k,��CR�!ض�"h^�@d��-Ԕ%"n8.�xELEÕӬ��j�2���mu�|��SA��7\��� W���`�6}fS<�m�G�+�J�y�ߎ
����Ȅ�P6�r�(R2/�1�S>�3E@�E0��`�<6�;ħV�i7.T���)��u�P��qwK�f��l(��3#󨪫F4Rnzf���Ь�����GN�ߟ��?`�q��,��2?VD�V N�ш��Г�l���&��pz,��&ފ�������[nm�?��/�,��%L���-%X�C��kfj���:�S�}"	�V�D"�i��W_&3M��D$Ab��WP~p�FM��z�[D��>��'|5�n�{�yl���|�TGtn�z�+���Ƶ�As�rK�C8�"^�yM{���$*ċ[�ct�W`V�����x���)�=&\&`5�^�c<o�ca�lX�47*@143���I5pw����I�T�J�ϔ�I͛~��D*&�T2',B��ϫ
��i,��du��|�A��(��������c�c7��WC#��Ս�z�n-`�I3e�����&?T9���Ys���{;����bZ��,"65�x�c(�@�o�������=؄��.��uk
�7��It�������͍��8��M��>�##�9�?e�vsh�'�YmJPI��1����"Xen�����6�d<��_�k�+,��ݵ�B�]��{ٻ<��-+��A]�ٜ��*���S��T�]�֋a�4�Csa'��b���*��-����fF��c��d?g^�ʷq=b�2�ɀ��4*L�;U'�����n���5��y+�r��/��^Bk�ĳՇ�_V�
o�Gn�[Y��Ne���"����86dmZ`�1�.E,z�ޑ�ͪP��锸���MUکR��f��*� �m��'JF�5� ����&�԰�J���T�4o��`c��6�.�շ���3�
���$��yƗ�����Ҡ����t�h��C��V�t'I�B�ڡ��J^s�=��@��u\����NE�0>�Uo�Ǧ'8|�2\���g.^��]K���
���E3(�d]���ю^�A�A-�)7�Q/���:x-I�9�#�AL'gaU�XL
Cm	gZ��Iz-o��";��q������Z�ң�.�~|�T���4'�q�Uw
�D'�OX�7��}��y�-�e/!�Or��g"F���=I�H@"�xJҏ?6���9̭���_�v�)d,3'�1�'ڠ�R6�Э�Y���]�������OfV�_�q�H�|�b#��MGE�ZTlam�wf~��a�\Q&��`�
t�dj�I�9K3D ,�������A�����ȼW&܉��D�䨤z�o�Zbo�;{t�
4�mq{ޡ�h��$��}�U	���@ޘ"��ë�O�d=fo%#��3x�i����ȡo�[t�͑ځW�e�n�N$`yf�h@kZ�ſ���*z���������pB�x��N%&�� .p]�X���ʡ�����C��k�I�����ieLeH��S�,�w�ڤF�{��b�5dT!�7W��Y$��|��6��{L/������`q�z��^ +�xb�s���EtF����2���W�y������^���x���
�b�*��>��A�����ז",���O�nu,^�׎X�1�F=�����_��ߐCb�+=(��6��0��EWH`9��$�1"4�:��:��v%��
����@��G��*"�
��V i0��/B�Jr��ev�1�O���>])+W�[ o9N}�����8�a�F/���D^�*̱�kt3��h�ٕh,�Ua~j����]K�Z��J����O�4,���l��.a�3�L�SK�}�;�p��X�YP����8"�&̼�=:�6xD�l5G�էF! x�&E���.ԲULC��7D�k�b�����6���툘�wP��~U���=C6��IbX�a����j��~�� �}Fp�����E7���]BHz������i!�TL'���DB�':Ƈ���@y*{c0��vm�%���V���P��܀_�Nu�VJ�W�w͑A7Rc�_ؽ6S�c�XEl ��|H�ԛ��j��Ԅ(Yǽof!Τ�_um��tsY��#���� /�C��{��!A�v(�/(��V�S�C�2�钮`bv�{�L�B�{�i�3RV�t��z�7ͪbx޸��Y�	�$I�����r����H�������c0 n��7��Xm��ɮ�R�f~-��Vj0Д��_&�H���m�H�`�,��j�@���o;M
|L{[[2�-$uI͌�nO �}�����J���ِ�ئ��c�GQiU��@���A�-�� b�`��;����f���9�z�#�O�%���-܌��"��"x�����'E��A^��ru�T�����҈~���΀��7��`�"!��c�u���M��t��sa����s>� LF!d�;�� ����&�C���3� �#�������2��a�8�[X	�ݩKO�p�o�q>jŕ������=:A�,`mh��[�$*�HA�B�,0&r�~�~�*�7X}^�X��~5K�q<+Vz��Hd�ڈ^��Y�Dp2Ɗ��4w�ţ�(���s�Oi?H��(��2���f;jۮ��~vk:��7aW��A�;���rVim�煨�V9N�YaK!0���	�� ����$���$�B�������� ��ĝ�d6V����V�S"
M��Ev�&!G����æ�&�3&j=f�G]ϯ���ZA�u*��|�=�4�Ο>.�o�oA�0'��2k�kZpBW~�n7��$w�p��_�����<�ru���+9��Ri����+Ud�V&���p0�`2�TK����;���\��H\?p��
rɐ��O��w�|��
-Jkg}���������	��,�7p~�����)]q����_����>�,��ݺ�Wz�����!
�&���f��AKdf�Uy@���H+&���M�Fy٧���J�*6ۈ@�W� qD�w�m�s�\��H��>5�2��O�?t\����|�G�d�͔�$P. m:Xr��O̢#�W$�bxM��;6�{�e;+O6��Ƹ2e�2�-�U���v����_i>^7�h	�����l��3�y��kf����÷&f>��e��'�����o��A�|)ұ��j6������P���(2��\v��[ȋ�1�k:���j�R�������QHJ��m���u�hܯ�4�=C_����2G��ufB`��4��AKNw��f�!.Iu�ɟ��\��Ğ#񔏵������qF��F\}�i�Y��w�NK+G���N��Ī�'��0be{+/G^���	��>��� �!���hL��QZFu�<�S����&&]�Ѭ���z����Zi���V�%g���;��PI�9܈��2�9Lb�&�*i3]bo=!�h�y�0ޥ��;F�]�y�A����� �њ�ʬk�]���t�B�Zڼ� ��l��q��x ���h�55?�
�a��6��۱(>�L�pY�D�� ��ް�T�!zm��dԪ�az��ʂ�T+�/kf9��v��[-�*b��b���U6x��YΛ��v:�P%�T�ϵ�͚=��M�T/.�.s1��_T0��©X����K	��FN�(�V]��n�䄎)������	�^��#�����v��:R��ۺ�& ���hM��hR�;l��cYb�n?8�7@պP"l��"���de25�Ԙd���瀏9^ h�.�4�N�'0�K{z��6�Hi|4�u|��H�etc�ZG�2�M�Ѳ�5�@��X��N���ר�F��`��^�Z�&Ն���!��*bʁ����q2
߁����0�c<���[������c\�oH?g1�(c(�ԟ��"^�7���n�ݵ�ᱷ�H�y�p�mQ|e�p�`o&�jw� Q/�5����A��,��?�E��ٷ�H���
��|��oj�-�7��*�٭;�g����jƝ�S����L�ƩH�"L%������re�kSq�>��e��1z!�k�,*f����_�ɸpϨ\A�W��Úz��z�׍"�%O(d0�+6(k[<��o�{ۂ�U�m���� ;�P��0�{s���	5x��[�h�Dv� K�F�,"���t!ےoe�j~ZF�h�.Nɀ��8э�d����[@b�8��| D0"�wϕ���A��r+O�C߈�
�u�<{��7��-��im��~Oy�o���kl,N�+��
<Gؠ�j Qi�k�D�b$d0".��J�x�;#|��y|3���8vʹ^�0�u3�G�?��R|�.���5��0����l���]�z��Hx�"�o���P�=r�h���=�G��=�]s>C��&J�-��>�ي"A(�U�o��h�B�yXr�{�q��Ԙ�����]W��wbv��I�G�w�ց��]beŗ7�lW�KG�F���{FƓP*4}�t<��/�Ul? ɶΰ���������Q���3M��n)9�%���EoG��	��j®�A��1�"y>Pj՘��c�0/J��5Y��72x�#sX!��+RDY�N��ІU��Wc�S�'ܲ�?o��͍�=��c����Hf�m|�=��qpp�o��	���!����K
 ����+{��V���L�~
?����&��0NOC�ƪ�ßs�q�ﺮ��P���QhՁ�5�u�h�H�I��?}���a�K���5 �i�W�&DH'��`��a� �"r�)�k�*�l6o�#�Y>�c5��P/�PY�au�q�osa���Ȁٴ����+,|�Nt��p y���I?"
ck���P��жZ/L
u��Ή7R,�ۼ����"�Њh' ��]���!�Y���?d����!�W,"|9V}�H�v�M:��{�X��l>k�[9b8/Mʃ��@S��	8<u���x�	����Ǽ���.��=���x_�4��w���CW�������}��sPFjɸ�J����L��A��@n*����]�玲�:�X�j���DN"g�E��J�R�pɎ����k(��d\5pV����+��k�(��.���o8�����)h-6��:�m�&�Y�� ���o�vɥ�ܥ�M�:�3a�U�'(��_`��b:�^/q�4��x�R�t�>{�����"�/,Q
E�ً⧅DE꺲~Om+�;..�U���G6�������j �%�.E)�I�_���V+]��D<�n������U:�b>�v���zѼאf��3�p(�@V���fъ3��5���K���e���K�����1}R  �Ɏq�¦�Y��4���7ƈ�U���^4Zx_��p�鐕ç�J����Ċ� ��_�gH^�rz�q�?u�25�-�{<@gd�c��<��A�$nuR4=B������F���-�g˓f+T~���G�<�7��O��̅}jm�����Щ�+��0�JJ�r�D�W�hI��h�΀�:��lm(��*�R�f 1WtI�����#��uc��(~X�ƺq�}~�7i�@]���xrƘ�&�̽:���h�~/�����iZ�0������$άX���T>��+
B��8���e��U��� 83}PӜ�V��5@�s�C�'\������/�L���ι@������m8g��Xs�u{��@��P��]��Of;�Ȭ�����R쁷�l���	9\/��gy	�3�>�;k4����v��b��s�j��G��7y.Н�>�2xI��rH0(v�!�M<V>�Ӏ����Q��)x�I�2��lk]�X��gr�u`~nI����v�9���j[�"+Ϻ�)l�v[T�$H$�� �LZ"�'�+=��KP=CH�E�&v
��W\Sg؂�9+_����e����Rd���G�:zk��lKA���c��v������7�4�H�x��6q.J�=�z���Z>?a��V�K]bѼ�W���K҃J�ǹfkXVf��T�5�܀���ݡ�A�2�&�cZ��!^<%���c��@��Z=2^U6+?z���g0
��=�+�\D�o5�R?͂���YR69� 8R�m�5я����`�P�eQ�Fg)R��I�}��梦v��V	�Cg���H�R�>Rr��uZ
�Q<:�zgky���ɑ�|�i�[a+����+O��k��e4���@�'[3�G���c?s���v�/�����b�v��t!��z������H�:�N�����|�
���}�vm15���� ��*���Fio6)"2����.��C�W�e��jXt���'L���� ��5�Q�8�l��hY�?]��2�g͝xeIp��2�LN����*�ƙU�C�W8�9���)�ŲQ'UWi7 ���������d�T��d���i��2��F ��t�8���l(��s�3^@�O`U�T����~��O �v��q6�4�L��	��O7�cg��!�h�aW�S��>��-��!��d�:����4�LL�tLBL
��HCY���!��&�f5���I�foŀv49�1�l������"$΅��6c�e����;5[m������ ����p��o'�7h�yܷ��K;w��81-�!ŧM���H|��QJA(��u�j�V|��߈P��6q�*f�c$�a�2�*����3��2��N������&Z(,�����-���A��=߱=�S�b����r��G=�m'Y_>+mp7�\zN��Uo_��Fi�,�=	O���bY�s�tW�Q�R|?��$?��ǣ�0<@�~#�saI�;Jth'�;���D�����W �LB9�9��T^�E�݀��
^7@�5,s�%+�L�&��1Fvd�:̦	CbC���|!����/����i�j{jņx���+2[�

�k9�_�zBdn]�����h,k�,����ӘRO�����y��Nw���D� ��⎔����g�箂Q��'�<�	������6H��v��Y'���,���Ь)��E����z�i%	���lx�hԕ*O��߇S�ų��5x]j�[�j6���A�e����b�O�b���`_߼)5�<wHp<��I?8y׆�xIH.B��,C��9�q�^���cwːL��()X�wWF��ѿ �FUө�N�U"��P����}s3|�0~��O(�e{��~Y�=��:>Tt8]���G[&;.H>�}��.Dog���K�Sw?v������	��oLT/�C�NB�:r��t�m��ܫ���,7��J�< �C*�P������1k�ߣ��z��+e��}EG����W�ɨ��������\��!B���@,��4�+��;��� �����a҅"C0�*#�[-�5ԛ��*p�H����} �R�}@���H��#μV��O��7�G�9<�w�:lX!y7�Z���y�E�T�a�4�p���$���2�>V�u"�WM�u�ұ�'1�� N
5�H�Hb�a}0w��c .>99�b��k��.H�e�_�3�H���y�� m`��Yp@��T�'9p̄Գ��f��0�M�s�	��o��/AE����r�55א�|��ݴo��� ������T�o5�e��]��"��]_��p�����H�=dl&�J�DsH|M4ʶZ�8�=��R�,�Z\@LJ6�Q�.��&���~�[�̊��b9\>���)Q�6Rp�u|Cɔl�E��LG��J6�	1�3X�f�P-l�]���x�A�<F�a��@��{�x����������iiaB����QU଀�)�yѰ;!-#�{�Hy��o
�������j7��䭘�>k��z�]7K� �
�A{�p�V��K,�L��hl�{YeN����`5*�B=�NLM�V$�͙EI�*@���|�M��9>@!�������(��;���{ƧV�i��S�`���Ȏ���� \5ߥMZ�2��>���ؐ�`4�f��*+B�[NU��JS��G�u�I�&"�E���Yaԣ���sTr������Q������7�Da���)�k��{,Oᜏ>%5�U�c�x�琉��X���J1޲m�������"�i�p=�s.������}5���x��G����4r� ,bĳG�6uV��l79nau�X��\D�.A9�/fq�3������d$��@��L�:\T�*D�C˕�� O��퇬�,�=�Y� ��c�l�7Îp;3��>B��y�2����m�"{O/��&�#TmW[�Q����s2V�;"|�6J ȳQ2�DsM*H��	5�l`������{�	�Xh&~
(������!��˛��0�U��3;=��'w���/��r���YwCvB��t��:ǎZb���&м������KY�͏b�����`��s� �M����;�����Y͹*�������I[Q%�Ny0��5�����.�.�P��WJ�Sڌ���ﾭ�t]w��o��WQB�0=�& 5WyP���AA�ʣ!�����Z�fb�� ���p�ظ�n��벧N\��kR�L0��U~u��M˚኱��E�ޜD� ����W9@��_����|P&�-6�ţ��&p,_}zIdv��?�����_������Bd�4�n�;Z	�	��E�Fo�B�O���D�o��L#:f��nq*��e^4�)�_��
姵s���5:��A�.��+�SUJ�Φ��9>Fz���N0�ߚ�O.�}YS�g��L�`;N����$��_@�1��~���0�Q��?+�t1�w��Tl�ZP0G�1^���Km�DmfQn�¡t�0T.�����u/R�UL� 5�.����y�"�^��e�e���0u���{LV;F�ȯkm��^o�V;�RƜS��ԙQ8��^&��l��M�`@��.�<�we�LQ���h8�Z�U��Q��hlO�:ǭG*��*�-d��K����؇b�2��W0E,��@Ԥtw+����Ul9$��@���0�K6I�.ݺw}Ng_m�:|z�-n��s���#��eÜ��/��;�׎�I^Mew��g�n�3X��ɘ���:��/9��*/����2s 2���Ou�͍]�������P�	��H ��X+M�a'Y���^��V��$g�eseC�K^6%f&&l��
�N�".d�i� ج�  ���x���8Y�7^ Qi@P� f�v
��g���k"�GM��{t:�����mmB+�����W���Y��w�KY_���\JS`�6�!�sx^�|E�n���{�JGh����k6;㵔mߧU������tA3vJ�m������A'�p�@%�D2_N�`��`e���.}B��A�=�Q��e��m��	���t���ڔ�녓-C��^4��RVH|cIo���jq��F��JL�@H�>�P�{��l���\zi׵�y��t1CĐ���fm���������f�����C>��±pN�BB�-9?As�9f�%j[�Ms�K��1��de�Jv�L�9g�[^�W��j���[ ?���fed�Qe}�����a�/@ﻅ��.�\Chk%����~b��?w���'Kd�x�$C���@���wh���>�!�=ִ!=y*��X^$�rCR$q����S�{�1c�'�PG�	)���,��QP����p�e�����R2� �������ٜi>\��u�m��[}���T5-���l(���������li��u5�F�a��<؍��>����P���6�w�?���>��r+��_P��֚�V��1ֿh�-�C�D�K��ϥ"����~7*207|/�2�hAG��F�濆���~+r7���P���l,<tx�̳'��95�k���ܿ.�T�T2�l�Ɩ����*T�ܷ(�8Kb���{�;H3K��SD8,s�(���+��HΥe2(��nG&{)b�$��+ࢫuJ�<����L����iS�$�2.�� D�FL����~�]�D��Ϩ�� �L[��DE&S"P��bem�xe#e����p��9��D�e��[dmH��n��[h��f�����y�\%���pJvYDl�v���������S��3������E��I�]O���ၔlB�1�*r)�#޵�����\'��a[���"���.D����FQ,�y���,���a�x�*��Zh.�VC��7o�����%�͑��j6Z��p����L���<p��Z�8@~�jH.y��GQ%����?����q�]�����D:C;�+�S��_0,�]dp���e��oY�B'T����6�oݲ:m
cݼ�{�����ڏ��_���G�:	�.Ϻ�4��%��q_�m&�: F>/��r4^��3�2����;�"�@�g��\� ���8�Y���@}V&�� �#����)K��!j���∄�_ף@77��
U�}y��!L^n�3i'A�y�_8 @2&�qL����{�</��4�o*# �Y0*#=������:�&���\{⇡�πvnM_YTIi���s��3o�O�{�q̚��k�XK���KC�=��0Nᔑf@�p��7�Ix/��Ƈ��5��8(��=N�]�%�㨭'����	�����)��e�K`����K��Bӛ����I�7ņ����QV�0�U�xZ>�I����}��Ӹ}��d��1gm��E��^�W�ǝm�����yh�]�a�c��,)P�x���k��Ӑ�$��i�Cwӆ��&�<	���t3�eu�Nk����r�K$f�й��6�փ�!�Q�z�}�F6s��U>�$��w3A��}�~3|����b��!h~@�m��y+�1���F�L��� fx�r��l����XE\��;Ee�O���[&�- �F�*�������o��uor�q����G$��>�� �XrȸOa��{f�$`�{2���q��^:�n;�u6�nfH��frd=�<��r��]�ϭ�*��	�2<��9�%��`�����	��AG��w�� ����b����5K�� i�s�i�W���m��nJ��|94)e����5z2��v�Q@�n�)M :�k��)z�����K��}#�����m'A��[WV܉��b�j��~�͊����W�
�18�2�����|�n-�o�]�����B��GN}7q�1��(Vq��{�<��7e�
�a���	���C���r���w� �M�@�v*�X?_�"�v;#޲� .j� ���Ui�8	a:�Z��&`U�F5z���1��e�8 `OVj����;��͚n�B(��=�u���8��&��Kd�t����zR�Q��а9���0 [}צ�������߾�4�M���N��2Y�o�{�,�����(��r�Su��O\8��h ̯��H�m��+���~SJ3�?��s���� �!s���i��F������/4�1E�v�Ǵ%�<�`�J�OhODo	4T����}�����i���~�\����U�LdS�����F����YQ����#��zs�w`�|»�#�[&T�վ{ӱI�]1�<����U�"OP�� �C��������,?!���g&�̭�5��j�-��`CZ.-x�u�^
��g7�`QC!'��A�:�������kZ0�k4K�"����Ǉ(�{eĤv��{!Y���O�.���t�,V��*�w5\�����6hO������@ob�zo#4dLm��k��]� %b4PD`-Vd`0��{�g1l�IL±a3����������M�,F��?2Cg�&Y3)+P�J��.8�0���f�(�'e_٠�3D�V��Ɛx��e@:K�A�k	��}�����a�袈Z�&q�OV��)fM�m45�.�����hU\�=�����7/5�)��B�Y�yG_M�����M::�M�E���/�6ZÞ1�9�]����W���S�~%H!���n���_�����a��׸k>��i�{�hy��I�����-"0���޼��{�\�������Ѐ�y�U;��M��@�/�Nю��#W�q1"����%P��Ԡe#jBࢇ��/�}T�cr���� }�j��޻a-	����a~jys��"ν4z��1��Qt
N|����06Ckϛ!�G��ё��F4�R��Ss���4V�7z?�gooŏ����mI���6W�F�L�묆���D}�2
�QGt}_����6�)�	!@Xc�j���s�~��l0�!Bb��68���� �	#X~��@�{�3+q,�X�K�ˑ�S��j�}�{.��R2�������/��T�ܭ���-7ő|�js4���ie�V�11z�YGE���Xg��Й��s��=H���a�M�A�<��es�ѕ��!_�	��*�0��7��V+�J�Okw���n�I೉fT��#�șQ)�E���vla�a��5��:5�&|/x�s+bP�?u�e�y1�G2E3����h�O��X��-��O~��^3⭈2�J��X���g#X�)0�>���K���NQ�6^[�j#F�+AI&l_/q#��q�Jo6�z3���0��^V�"��X/s�8|�̎�w��"�m�� �H����(��mȠ��-���xE�M�����|�	~����P�3����˪Q@ac�3��tۥvJ28��\pW���ɂJ�q�����}o�֚��X��q
��e/t�.��6�h�N�`>i��C���J��]��@5�X2����e�pU�-vM �(��&R2M�Q?I���<����b������9�u���1F�u�p�C:�3�ը��.8�巯�7Ökm)?sS���>W���uD�2�1f�B1��� �8�ΏD�����v��Ϗ浰P�0z�%r��^�]W�P�Ɍ��h��<.y`�4_g�y���+��#4��+Bߏ0�U`�m��w�h�*�U*uh�W��8�YZ?~�Z��42��ZԖ��h���N���:c�|��l^H�-32���fB��H~\�{9+�x��Rv��"���g]H�[��f'jب��+8;�*��6����U��;�M-�0K/��w��=t�mU#�����o�_�I��4i�G(��ň�&㳋:�Pc�aF�с�9鞄�}W����*�2�1~�W��b�ɲS���?���1�38��)�E#_��z:�yE�zB�&����3�T60�����ezy*��j�W������S�6ÏmL��L�G01&ݵJ '�͡wx��*$8`����Sd�O�|V���
>'P��<*J|n��8�(-�@u����MW�=|��v���uLN��>vH�h{lz������<�yc���B0�8�횹fCb�ӊe��iũ������K�>����Q#��B�E��LU�$ �H7k�(�����|���i�ވ�=��u���KI���GcG�U�����/E����&y~X�V�^�S�%LrE�f��b�^c����x���p {����,������P�	�?XY��-R����*�ezqh|��I������8��zX*�T�fW]�iElHz4.Q[J<کɌo����g��X�P�Ş^J#����2��y�Q�5�_o��ύ��K�� �r)�YSa�a&�����zsi��m���!N�O�Y�2�+l�p�o*��+�[L�i��8��m��������Hο��{$?��|�y.F>��b��"L�_�g�ιm�wլ!��#�Tg'�T��9���/��<�C�'��^hK�l���vt��5-�S)=3K9X��Fl1�-ˊ1�����Q���?dq��eI�t=/�&�Q4�ӥV	�098ej6G:���1�=��l@���ew8BU.!�zv(.�B�֟7�-���m��B�<Γ-=�}���wʵ
�$ͣA��f!l��Q�6X�U�{Fw{	~�ٰO��ނ<���m*����������4@���DE��pp�̹pk�6���.����'8�'a.�#��ink����p9�j�ԘJB.*>�Uk��TU��hz\;d���.��	�j�%�غMԀ��mg�J̦��̑rY� Yl�%.�7F�)0']�jF�cc%r&��F��2"{��鎊�0S,����/�<�%�7�I�x`�Y�6[p�"�3�aT_�	T.����W�D���pk�y�|/�ZR����r���w�G��"p\yٿ��^�6>f�]��Y�tS�2 �	}g�o����iQ���_Ǡ�w��K�o�P�%�����..����`�T
��l�1�;<�Bٗ�wbɃ����ʻ7���^|Л|B��_�����xE�_cL
�:/7�.����篨��.Жɭn�a�%�����D<�a���m^�>qL�b����H�qZjͨ�_6M���ZP4�/���s��6��Xn.Dl����(��W'  \�|�/��tU���L� ��̀��_6����ιhtq���%��C�|�L\7�� >9���ct��m��	��X���:��4�Y�s��&y�ة�z��Ys�c-
|��
��K6'Oˠ?�yօWD�����èJ���ɤ� |�㨓ZLpr������3�2��^6�{~LB'�A^��#!��������\�g�����`���*�YA�2�-"Ư�(аb
]���x��&S;��i�Kr��x����Eۇ��熎;�T挪Z���f�CK��xW^��Q��O�`-�5�׉�$�����~��,�fy,��d���a�v��Pn#Ѭ����<�{e�:�:�C
�b_:$E�%�������lz�sXh0V����E�����.l�f�����o�V �,zo��c��O��I�ۻ�e�12K"�����Q��fڭ�|P<ҹ3z�H��ܧ�q�|��Vh�]�d���U�)��P}0Y�!������L�������|�I��5.�����:C�{���eP�,���N���\W�!���z�gPn$�p:����4�E�|�HT��%��vhH�C�
�`���+�
D2��P<�&�1gS���(�_8R�^��R�{0ib{\+����Ej��qQ!Iܜ&^���n �VcAna��V�W�o�c퟾Η���)��Y���h7-A�
�.���\�#?��#��̓x&y��9��!�0�u��J�*�\|l���2 n=� =!���+�t�ւJ���A��f��`���7��k���eaG�{Y�X]���U�a�X]���4#�޾ {��}`�ŧ�A2/r��%`��͂���f`@��/w���r#i_5��䪿9�\I�r�k}Y��^���LP	y���R�B\*x���[z1ʂ�����݉���Ӹ��3�ř���In �.f{�F	{#�UӤ��4���9/R�"F�e�˥k�-�&����6����������4EإQ j,{卥�*�3��B��B�HL�ڌOM����i�5Z�=��|����a�����e&��c�a�ʶ�ΒW�!��7#�������~���"����ڨu®���*}��}��*A�.���9�Q]t̛����r&�"$k�Y8���:�Ԡtyt~��,�n��#W����^r�`�7��}0#�v�ۿ�Y��L��;7�u�������g9�.���o�
އ�me	�bj6z?�'�T&?5TrC,�g�s|*9�p�1��2�5��UN�����p�#�N�y[զI���BE���\RJ��wg�@~�;�)��Q���!�|<9O���{1�9L8���y�)��/u�5;�+�q���U�5@��Uo�0ТP�<�S(��� ;��pj*�"�M��}4�JNx��0��ZKLΔq��++<mQy��������t1���b!��3�3��L����c d�,j��dVA'�f��H3Vl�Y����(|8��C�D����C�p�\a�(�a}e���1ѤR����{��]m;"�2�H��ZGR=���̽xtd�̊�OHk�����l
-�|�V��W��wTmQ�:q'�uC1)H!q������M[���}6H����t�ܩ�~��-x>C�Q���
�8����#��N�X�Vu�0�����G�#��6q�l�C������<��L@f��v�x�ۂ2�KRoQ�xθ�ڿ�8�M��,��_����8���j�qk���Q�ـ�
�[��&�lC@�qo��ه���R$���6�����w)�t@^�,�HK�P�v;�I���+q��A$�y߉'�/ۂ͞+R�����lFO�8(��6L���b��Diwm�U��Ȅg` ���^I�W<�;`U�z��i3
�����L�?���z�U����>�!�y�_.WP�;i���l������ �9���^�0,���Q����)H���/i��>HZ��6��c��|#�&��˹���^8�k��T��P�q�L��j���MJ/�H��V�^�w�S^zF�N�W=�~�� �1��,V��-#������� 64�c۔K��}W��V���`�#2 �U$���I���h)3L�A~�����.������b��H�&��5|P��t�	vt7^���P%#�z3׊���F�x�-�S񉵌#�D��,IBs�E����~�}o�i!�j�1�a�|���{NG�4�L^d�?T+2��u�F�'���ƽL�T�MTW
ԫȅJ���3{.�^����Zud���9�݈^�>c8�$"�>�5,��-���,�EW�D��%8.�2k����ܑ+r:D�pZ�m���"�t��,P�P��Ы������%��7�DV�>{�yX~�LX���������?͎�g�J�fL�<AXEH?�jP)�-W�Fu�(� ���M�w��~*G'|���/+M����������e��z�P��dᶟh7qy=���@����;��h�
�Ì?Z?Z h�`����77.y;�����>�ʹ4mu&�x��GX	������g.�?PA���'3��е�{W�A93�+�.�2�:�] ŧ>r��
P�R�B�U2
��}&���2�Nɠ-���U,L�����~В��2�+���-�{��@M���>g�MO�����W��2�]s���M�>�׭��+CL�8��6.�lُzq��4S#z����x��=u��@d����T�fІ/q��jo�_]$��[rd�ϋn��������oO7	���T�͵��x��|@d�r@�5�K��GXU��������8׊"K+vWSo��p	w���Ւ�JìrYE]�����vsX`�vu��-����K{F��/Ba,���6;��F�|��(4�?1u���)̟�<'����5U�1�w�8G��7��oLY�N���ؼQGS�Lڌ9��A���I���.6+֣��'�M���yY�4
��{�O���-�υT�o41l�"R��Kd]���B��Z�;����b����\��"`W�f�w������ҳ�N�,�*O��Z��Xӷ�� y~�@r՞�I�-�s^��Tp@�Ƀ@�u�|']q�u�#9T�M�G�2�J��M�M���:��-��p���n��1�n���`�JR*�'��Ю*x�*'�Y��bf�m���7�г]�ć�A�+�cp��~E	��NF�U~�5�p��I�q�aLRU�0	~��lKn�[3��i�Qq4✚4�=W��9{W��I~Z��;.:)v}���+�dP&�v��OA!�no��p��<��'X��s�A�3����:���R`���|��j��%�����6��z]qL� ���ؚ3�<J*�7{ڴ�J8Fr#�YȴS�:�^&l�)����1��Q��~��9g��l�N	�"mIz�-��3��,�	�y��l �q#��2�M���� �q�y;��_�`�?"�����i+����
��EG��(�^�sE�γ\�(��/�>5%�)%�2�n?_tn|�����:Y0�"v����2�X�����QOn�8C����־�׬ ��Mr���L�0ffZ?֦qW�7M=�~�H�T�`0U5괔�e�a�WF��~/�����XŚ;�� �c����_5u��6PD��}���EO�U+#�	p���NG(��(*��N<�����	��2�5��+j���%��Fl"�?�;e2Y��Ô?���-B���#���p�\��>�g�m(�r���`��p�� X�5�s���K�Δ�nG����Svw�|C$�l�/,�❌�P�D��28���O���Rhm)ψ�!a��)K�,`�����f�`����@Xv��E��>^ܢ*��d�`�����Xˌ�DNAy�%�p��&��q������$�Ee����ޱܠ����ײ�E���^Y��h�
B�l���}�������b�wm�xB����f/�u��u�y�q��y[xR��<v���Y���6��L�<�ى:�fB�b���'�N�H���D�(���)A%��W�G�}����l�����מn���Ϲ������)հ�in��.ä[{�}<��04�S؄�K�n4�_��9�ʉ��c�ҍB#��H��턴�^�g0���ul��ãX�I_����S;P}�lY�ŭ���fp63���X�bN�k+DŰ,��?�0�E���p�Z��(�b�es��]�L�O��q/�b����񙶽!-7��׳���͝vL�u�v�3YlcԳ'�}�-hcY�:����R:]!P��{�!*^ � �yy���eS+��1>���C��g�f/St�U��'��|��澕�Q�Q���rS��:�df4�. ��¢���SNBge�f_"_v��/��".K�m}W,���7����W"X�c�Z><���)��:^F�{�]Oz���b�]����r3>g ���D�mX�S�/��ܾ�}xl'��)�o����3���ݮ�������O�i;k�sUf�� � J)N��c�N6�
u����)$R���F���$��H���V_�yn*�,��,��a�#-��`�%�˺��}��;;����(���2����B
���u�k!'�"�:�����E�����@/�!}Ѐa�*�كKz���rT���Д+Z���Zg)��M˗�R���;�1�s�}X��u{ih�'����W?��	�����o��0�_%����� �;�}���lF�3�:*ժN:M��d��ȁ,�2�X��h��jr�"
/�#jfp��/^�5�6���[y3�|<ݑ_�p�Z�$8kD��9����#{��!ķ��i✎B�Rê�ˎ>~�Ǳ�r,F@�o1�z�=�u�����������Nl�؃�9�<A[h�9�����y�ҩʛ�2۾�GQGV��,z5Me�� �h���|u8<�H�������@���U:���4}�E�"�4��_u���<���6h���yJkT��=]S���WO��&�g�s>�H
qs�7�%,FXچe�k���z��jg�П�} d��W��y��`���!��;.�th�������1�j�rzO��ɱمm�>l���ڙ������:��%B�,M��"J$�N(�~�/z�zF�֫I��T�h����^�����v�o�g�k��Ɩ��`�/"=(�ѵE�kPZ���s(�X=t9�(�C��%�N� P�cif�A냟�՟����?5Xea���N�I�H�
���1*�ڛ����>���+�h��Y\>J��d[^K&��P���z��"�"�;�\H��x�>(�f��G#�\�_,��:v�/a�1�ngBV��s{��JM�q�%�}�7�]k�����Ek<���;,w�&W��)�ރ�Mԇg9@�����C�w����R�p�6$��S|�� .D�1�j�F��L�c��1��'�֑�U)��t#��]���*�
� � D+f14�ug���a1-:��'e
駠����G��L�V�i�u�Ni�	(��:rӇa�=1jB�tWa��I��!S"'�5��j�zi6�¶]S�����t�9�G��7�:�r6�`�4�@�ÿ�_�9.Ґ,?��?"�K�:P
@�蚊��/sBXM��9��9kX3�ű�E�GE��YK���*ue1e���$�Q؞�L�q�T��N+���w��+���o�ڬ�����#�3,8x�]��19���)�;�q&N!Ηv�i��7d*H����:�Tn3o�Bv#/Ƣ���?�	�(��ޟ�^�{#�� `�H�G�:Af�����ws�`�8�wM�tP���$����\ө�I�r���i�ߛ��9+$7-_<�3��a(�un�s�d� �\�j���M�">�	���a���	�z����m�����v͠�3�,�N��4՜�R�;{��ٸ�,�6E��,�X����o�6j��$<�U���
�<�9� �J?�2�M��2+G\���5q�������vl�T�ȝ,\_�F��O�%,ӹ4�%`�Ɨ��ay�m�ڱS���llD��R*����Z����+�(�˿G����A�f���5W��Tb~��nSWI���7����L���K.����#�*�zQ-��Og��J������UʾZ��T�x��b�Ql0A|]��%�S�xb�da�W��B-��d�?��*a̬�h�6S�x�����1�a�#I�i�>��Ί��������*��P������^��lW	��8�,�	JI�%z,�����%2�T��� B�A�
^$�I�Wo2�����a�N�{r�g/�yN9�5C�tP��fL�;^�����}Ѱ�ϑ$h%h�G�\�>3k���� 6&"�O >�d�O����-�5�?�k�N|ɻ\�
�"�L�Ix���9\^��l��~�����	��i����Ӆ���hI�>L�U׀�v�<4��B L�t��B����&:'Jң9�Z��nz�Ҍ���^��3˨�)�������`)�cܫ�,]�o�r�<�v#`f��nڙ���Ǌ�j�$'`��:֤�{�ZlŨV��'ߥ��|��ˡ]�&��ֹ0�E��-W�����ޭ����
p�Z��5�~U"�fi֪������:ԗT���rhM�v�w�/���\aҮ"�\������sS2{�$�ʂ(����$�?(�q��c�5d=��"^Ô��n.@�|�W�L�����̀/�>t�r��2If����)\�����L��O',�ʁΎSK�M�#
n^X����)�	��
�!�@_c�L#X�Л��5et��*� �W@��h[X����_�/j���YA��,'�����Dۄ;�kd�W}@���[ͱ���~��7wґ5jk2xYRD�����܆/o����/�6�v*G�$�X�M`��	u_����P�6�#��sK��1�$շ͏#�MT	�B�0�~�Od��G��i�㲡)M���y�Z:������Ψuq�P�fz��E6�X�o,V����ֳ�C��)��
�2j5��㲊���(hSH�u��μr��.�y��p���K�9���֫��4.�"��p���!#�.Fd1Ծ��\��I���j�&�p^N�nBs��R
�ڜ�^ƺ|��UZu�ǝnZ(<�8l�׋`c7x�tD�D��twa!
~�Z�zR�/��I>�/���,\`z
OӉD�c윮��9�e�$����X�Ć���^40�9đ�>��0	���i�͘����Z��;b�&��Fc	�*CvEJ�উLtإ�C,�a�m+��F���Gd�Qe��r���^ #���p�3�r�׽RtA�
�zT.M`pu-Ƃ�ѽ���o<c.�T�>���t����,�I`5j��M�[e��㻷���O���i��C���Q��g85�EP��n)��!QU&�/۴ql�y������_����jd��h%�-��4�w�?� �9�?�F��C�AK�ɢ��Y���'@3�Iv׷R��6��`D��N�W�M���b�bt1�[�,]�[��1��@���rP�q|����/T�kK�zz������QTv��q87����lv�}����<��}SAiA��D�_�
G-4��9� 4#W���K�Г3q�͇]�,O��9"�<۹|�!j֨p:� _���5C��*��h�?W+f<<�)s���e���� 2�`�U���zվ?ֹ֬�{�^ӥ���Ie�i���u�����T�&�s��,��5+����:߀&i�6n?�9R��(�n	$m��]�I��J/q�jg�R�O0>�(���H���J�>%=�x���[C_���ޏ	AT�3���iY�W�}\#��}�}�i �ݏ�:7��̔n*j��FJ/wC=چ 50������wiTX�w	W�ϟ����(6.�֨+`��'�瞎�HF�S+�9����S؂C���Y�_[�h�O�1^�2�D��[���`P-~�d�Z�,��V�pkؙfQ>_��b�"��Nx�s0�x�M_ȴ��j��������T�Q���uU�M������美f�әem���UVK�h�"�����0����u��Kdf�J�O�>�|7q����/�hZ6��e�b�~|BL����0JS���'�Ըn�6����܀���%
�'?=�vV���ԓ� =�Qx�{y�'@��.�qtJ�%ə;�ҷ�O$�6PX��O���I�߾�ncTh��%�%e�Jdi
����@H� @�?=�䮢^���ݽ�XW#��&�ǵY�s~�\���9.��.�A����� "_m	��v����	|��'s���<P��a$�̫��\GDo�̃ �?����9���[lBz�3��m'TO��M'��n��4�21�6�Ű���'�A�k�j|C`�o�ݢ�8�W[O�'P�*b$ѩ�>��#D�N��P2�g�S-��]j1ͧy�&m�@��'�NGE�r����V�O�=@�6z�T�H�D��4/������V����SQ�c�y��\�*�m��#�#�Y�Y����o�S����8�7�~�wWWX�@�q\"!����}�0�d���u%�!.ۙ�I�(���r�Y_�P��oT��u�(�kG�<VzId�G�!z�W��63l=�@�tf{TF������I�xPlЧ�����:�ӓr�} ����К�vX
j�[��.�6D���g�u+��S�#���N\� ��XF;��m8����	�� �<�p�<��G�Mc0���ؾ~ȴTL�+�,��5h"� ��t:GY�hN����>�@�L�B�~�򼱇�S>:AY�Qk�Y�Ǒ�U��]��%�[o\�#��x�7�+?���mٺ�%80�g�G.�O�^5����A��:þ�� �MrN^~��z����9u�X���h��yn��������oW7���g�M�(u'm��h�T���8�>D�l���%�G����<҂^��dBu�؎�{���l�.z����UXR��F7��ǫ�d����I�ѥ4�����j�4�ps�cRp���YHr;��z��q�^/U �u��v������_變+�P���Ur6ɜ������k���9f2���0Q�hu�Fk�/9��^�����\38�o|���==0�U�I��2���G~Z6l���$�6��Q���ʗɥ��S�|�i������0Q���=�4Q�&-S���-^�8'���Qj���+���L��;4���6\� �d��N0ۊ����aP,I�^��l2��A��k�'��*MH�����!R{�PڱM/*��6#(͙�t���S���"�n��Ohe����^|�-Q&:\]��<�p(����R ���U)�qB/d�ma���P,�	*��ٷ"�?[r�Hk��D�335������c�����ٚe��rd,�ռ�T�>n<QLP��!��l���^�.��&���7�nv�����7��>"X�O4c��%['��g�A����U��?m����Li�슺h`��<F���̗��p6�n �����2Kd	%޼2HQ�G��瞧v��'ǁ
�𚪒����|b�wO����/nX��O)Q��ZA}�S"�.g�<gاik�����3w۫$?�����ƫ��'7D��Gp�eVv��(c���Kg�42V��&ؾ�5��#����/� ��^-~��kv����m�uJ���s�S�Wv�Q�W�1��ጎu�y�A�h��^r��i�J?l�Em�}2gz]�p�L!�8f1U��&z�oYW���&�F��Ԣv����uE����iυ�}A�W���b]��@ݘ�!Q�O a|_V�G�ۼ�G��:�d�. ��>8F��1���L`w��?��P=�'�8���΍�Z�>��e��n��9�L7�.��HM� �m�>gs)��[�-	�"IlZ���{hA��-ħl��{y��a�sr��\I�U����iᢄ
:?��򈊪$	�*�OjT��~`(;כQ���}h��3��Ֆ���\}X���{w�(����K?��E	�E�H��h�=�R}kz�x@�2��v�Ԋ�k��^9��|VJ8[o�� 4��Y�OP�CZ0��M8��Zbq��ӿZǹƬ3��	�K$��!IH�5yT��[[!Ȥ��V���i�E9�ı̵ɒs��!���"��p�&�`�R�u�C��&sVx)�������kYV�a�9r���;1`Caf��7G}�o5�0R�G���(���^.� �$V�X�ir�3�J�
��=p�e8�aϓ�T�	�,>��Aĭ3.�$�|�����l
y22W�a9mk�+� n�NFY�,���\w��[�_�p���/��c�`�?(��j<�[T(
���]����sb���qE]����#�<���-y9Hm� >���Ar�j4���#�@�
j���h�`�{��a{�%g@��/�K��J��M�6�5�����,�C*���\���J�2V(OPb��KӨaGv4&���n���fd,����~p:{;�6�J���'_�xiC���
�P���S�AWBO�+�p����U�-m�1�;��[�σ�Z*L�<p7�������fz[�v~�ig �_$xʭg��2���9rFK"~�lIj]m_:��[�3�S_�-@�)4td@F����I��]`@(�`�M��K�2���o�gr�m�'��#7�n�(�d���ڮ�/n�j@��^Ec%��;�5'��Fd�}�K\
� ;���`�
R�Ce�sV���`.��Ͻ~�����T-�����'H��e��!�3ŉR��>6ۨgJV��zo2�]�{���/��<o0B�^��|��os��SQ,�4�u�����}�>nM���6A���}��čh1{I�DW���GX2�̎S`W�u��c|#:X����F��H�#{`�uo�ؘs<��~ߙ����qـs�}�/&����\�滌�+��?b�q��ͅL+�9��R��MC�Y�7��'��*�^��rI��Z/nF�~� ���J�o4~s��@l�B%�ъf�ʦ ��dl\p5��{[�J�3,���P���A�b�	�k,a"Qm��JF�k*�Y��沲X��qn��-�����1+�Ah�9Iq\�����fo��9yS��n�BQ�A&�d��m��mte��{x�A,[ ��V�a��j�Φ���;b���eG!o�,��ؽ:0a�wA:K}��g�m�[d0�	L������D�v�	�ņ��s��X���?,������.��Ŕ5�L��|�d@LZ{��'fB��r�0-GM_�t��6�K��;#�Ϡ���/q�U��h-M�����N����qN��?�5i���o��bK�j�+�S��<�����At=n�N�p|�xE�xx��ۚ�A�͋�K=B�Cl���@n�6�֑�	_��NޒY!E)b�#$�VL#����V��-ݯ4�UX���T+��4��'��Zd��/� �b��1j�e�߷Rmj�ERՍ0�Хz�V�
�?�
�8�����h�%�i$j��Xu�Ӎ�Rw8C��.�$(~�ub`X�6�6%᫝����U�fT�9�p,�����{�l�A�s�����Śt&ݛq�b�{ӥ�I�-�;�ݮd��x�Mҍ�L|E#����"l��tHb�w�)�n�}1��y���1A�8l�C׳���ln����8ġc,l@u9����p�ԥ�](T2��\��e��hў\x�9�4M�e|-��s��,A7h��bE��������rB@�L�!T�Z?���!�R�ٟn�_�wn�����<O<�Ѡl��4����!�0y��"oX%�X�\Ц��W�LŅ��Zj�W�z<���� >�.�ZAjБu[�o��-c�����%ᾸT_`�s̤?�xu4NҪ-ǝu��";_���Ң��]P7�*��"� Pd���p�%(D�2b���8=F�J���Y�0g�_�����oeL�စ1x�&��1ד�T�d�÷#V-?�;AH�AV��E{D ���{���r�T�����.AN�X/6�g۹����O\��GB̍�@J2�!���M84���hS�/�M��*�:��W����DqOCO4��<���Q��G����z��C�cӟ�P��.0�$�è��Jp��^�j��.0������K6�OI麫�_yT.�M$��8�c�)_�li�"5���]%��u	?8��(V �g�.A~��`��v�#��*�����O�\�����O��
�OА�<oc�bXF��Ek��l�QQyS���V�M<=�F�
P�뮐��b����-���E���Q���7���w�T���`���@�5�K�����fi�����<?�V�J&�+�������qp`��hWd����;|A ����	���yb3}���*f�
x�\YRQ��#`n�V�Y?�|�ާ#�k�o�앒E��>�ql@�P����w��EP9�O͗�k_��%���Z�r�`��R���?৛�A�n�W��;��f'��,&�W�% l�qN����2���駞U�k\�dK�n�y}3�Y����{�s+�-�+�7u��D6h}�����8�Ҏ�m���TC��*���~�.� BI
h��g.M227nJ�%�o�/�&M�c���
����A�/��~GtZ���|p	]����6�)!���o��s��Z]���&b%Y�u�L]���Ggg���ڳ|z�I߰ ���0�%�^W/��&�Y'�Yr��1�DC]��<9%��	�K�9e�dt�h�	�j���ȕ	 ��E�##�H����D�}���Cx(�J5�wڗ�A	�Qu���!�J~���.bO�s߳G�Q�Ħ�T��+l���5�8�ƅlcA�{�z"����6��we�I�_��,�j�h�~/ɐt�ln���4b��T�8�L:�`\ݮ����u%�?Q���$T��;	4�����ҭޔ�����T��5z�T7E:na脩m�>O����ao�K�R���A��YM�[hH7�ch
N��\iw��Υ׈�����^���4+�l٘��&9cj���6����W�v����n�T�6Lݦ)�����֝���`[[����p�� ������2R��XI���\|M�[Lw~�� 2{|ҽ�0%�50�Lzv�]�|QԤ��?�J�����O�r�Ia���Fѓrw�f�F�x�]ٰ>�)4<��p���E*ˎRh]��؎ޕ����&�K��n�p��H{֙]ƌf� oW�%e\;����(�����U��m�?��������޽��@r��l�B6U�d�y(#d�_k��A�=��j�ngn��FLz���Z�y��u�1X��6,Ğq���q2�u�Pq�Z(�L[M�z���iis�e/oz0���f�D�k����	���G�&G��t����;]2�!��L%i���2k��H��2(<6+r�bW�k_�����
��X�1��+ 7� 1��Nب1u+����I�@����^c�U:��=z��3�Q6�\�rKA���R���M�R�j�ǟ5c�װ
�V�]�~ˌ:S0������Q�~M���|��q�@W�q͹�;��<�����Qm���I��!+���� ��դ�mX��<��T����4��;��f7���G�~ vh�g��'�~���O��+����u}�(Z<'F��Y[F������x�1-�&? ��Ճ}\�>@���.����Xa` �,r������j�7�^�k&��-"\�-����|[����^�6<I!�?���m�tmaY�z�&U��{)q-X(��w���r¥�^��Ѳb;j��8��L�/l]�v�ċW��Mr���C��p �6��r�47�k�7�(q�� !�go{�Q
LXc���_���yw�vB�����q��N�J?F"r�~Hn�l29����n��tȌ�\��	�e��0�)���&�V6��?U���M��z���!��be�@޼<�j��y�r����:B��y֢s�N�cK;m�뙳}�=����W��F���<J4Ai<��5�D���%�"6j4'���ф<*�w|*�Q��4fÆpIQV�r���a�&X�A������/��PQl�U���d��rvL����%�����nT«��K��Ǽ�j\4#k&�`�w�^ቃ���A�;�s��g����G�C)[�i$� &3s����%���L~�txLM>�l�	!�l����yx���30�I�)&�w�?���cm��A����Z'?<�d�X	���{x;��y��k�KX,�@<f�Z��iV�D�uCp��Mߤ=��A�H��a�X�
�N ��2mHD5s*��i�v�gV�K9K�ONTogV�����L�Y�R��O���9� O�q�jZ��;�dEJ���թbOL�ފ����P�E&�w�+؉��{O����%�2y#&s
�<v/�}LJ�۽�
X��=Ǣ�^i��9�8&s-�u�^��[�/�eNZR��M�k:�MD���
�U� �B���8Qw\�b�Q�<�ݥ@�������C����������e�w7������(�3m��
@�h�.^:��e��ΔBbZ54�rx����Q@�+�@��w�������\�#�e4_�&@���_U�Z��SXV�e�:�v�n"��l����r���	B����$kUU���-;�僤+ej�*<����'��Q�;Jت��mM���!>�i�(&���um�tb�T^(u�ܔA(���$ΛVJi;���	C,5[���3�χ��Eсm��0d������n�w����?Ǭ\�\���=U��qS�[���M0">x����>�E��a�c����Sm�/f(Ч���j����F���D\I���ȏ~�B)^��α꾀Uy��\�>�65�~�1���\���8dM����hϵO�2̢X3v�K��$�#aB*��܈>�����#��4A��M��3Z��1� 2�U7YwP�Қ��MΌ��6�p����a(�/^.#�[�2��6a�kf%�Ϧ�K0�D��	)�1i�f� �-Ac�P�4�o��ߍְ�����u6�4l��Y�H9�0}N�@��h=��:WN9�]�!��&����X 3�C���6���o~� ����xk x��a\zY5����:��٘��y��-�Q�*�T��PT�d�]�]�*��G� O�p�Y>����D��^Ɓ�;�U�b8[1`ju���(NfgR�.(Ꚓ�u�و��tm�&��6rc�^�d���9>��Y��ګq�����($Њ�<�A���6�c_�1�v�_,��.��{���*��;?�J���s3���:�(����>=�E�N�u�`r�_�*W>�n���F��1t�3C��B�z҂P��Fh����Y�$�0D�( �0­Ub�H�2�l��h�>|�?3@ԣqQ+8��i��6�u�@a�K1)��[n�
�˴Q\��V(�u���'�g��ܷ��s�-�W��J�W6y�G*��(VP`g�,�P�Z�T �wT�ظ0򏪸UV�&�
F[Q�T �˄4u�!zO�!�G��q����9������P�j��gb��;��7���.��CF�M9:\n�ť.	�Q|Tmѧx�,~*��i4��� �Z5�e���MYF���P�5)O�����\�"ˣ�����+0��x���ĿØA�uP���/�$�q�`y�7	q�O��Yږ�2l�L�( ����'O�D���?`��S�q����A0��6W�'�q}�S�1��:1cv~/�>R��el��t�L�^�����&�*����pUI���z��Vqt��t$&Ƥ�@��i� �sĘy(�!�r?����>�=S:-��?�H��D=9&͐��6��Q�N-��!�[Ք���n���pJ�[U�9�����0D���5���l G��.Ov�lã>�����R̼?a��&i����G�)���Ǌ	���Ae�x���g��n���,�:���r,�mJJ dN�	N0�em@�r2g�E�i9GQ��r.���f#j�lxib�zh&;�\���O��w���ט��犙�3s�i�+L<nW���k�w����7\�A�_G鄍1�����ܢp��֭4[�\���S��qŲ"�A�ܾ��nA���i[tF#5$�E[���>G�:ߙ��|�z/�:+�Ҟ�|:~��`�P
��4(*�Y��J�t��B���@��6�bm����ͳ���v��r��!��E�gSi |I�AEBsS�'9C��/��ǖ�g �+�U��E�ϗJ%J5�k�$}�3��T\��S�C��&k������R���Y���t����K�,�Id��x�`x����F%�"+I� ����m��1ڝ�0��,\]�G$���&3v�@�NC�R��8]�;���Dx��x�@l߾:;U�Ԕ���\��ć�����۴�v��7��"��$f�Z~RކĿ�"����J%�/,�Ed]ut�{��7[d�ܶ�MH	�H"�0[/�?�N�V1���z�/L�s}b�t��k�����f�e8=��!`(�C5��w@������	��X�Zj� %����oñ�|~l��T���^^�uΆ��Gr{_ZȄ�_r�#����;QKb���֒9�\~M��!,s.� ��M��Ў4�~ x�S(ZA[�/��-�&Ƙ`����3�;�Tztw�4c�c���#��w���=�������_�Vݒܤ������$�o`�����x��<��0m_��,8�_�7�\�d(s�o�a��kq��)zb�M�|�w���(�5�w�oQ�!Y�37U�Nt�{����4-�I�S�Nl�l�k�q��h"6��J�� �����q�C�<z�[@��]��	�����<=j�9�އ������YrV~0����!1��4^�b�s�0��u~�����/��|��5�l�p��~<q�a��}Ӹ1�Ûu���������=����\:y�N����Tp:M
]3����<�Zt:^h�-�_�BnyO�'5��uH=�޽��aU�I��v��5���&u"��j�CT����z��J1zT�;צ���K~��I��
MS�y�89���9�A���0v����q�>��*OP�_���Z%I������=�yy�S Uwe5ع�k4m��(�UP*Ʒ�k3���-��5]4�ёa~��a�䢄1c;�DJ�9KLl�@W�R���䊷�۷?�1��3�C���BQJd]:������_���b���]�C�>���C���W98sc�<�X��7}k!]�t��F���͌�)��y�)��Y����<\y��?;���m����pV%���^^����2S���ؖ@(e7�?*�p��<IUS�o"_	���,5V\2�}S�^L�
�ã��Fq
������)+hT�ӋogLL=YuKJRS3�<fcR���Z�U!;��s���x�5%y5�f�d���;��=�Z"��D���xjc��4��PC%�;v��d(^���MV��b���ǫ[$��CT	+I��y�\��	�L�%�A�P�ZR�Զ��d�	�]�`���ٷ7�u#��Y�t}�Z���1�vx�FgP��7*�n��J��[���(�nk�%��ȭ70�w�j��x~K��:��ȠP��������gwl6���&a�=�.@@E�Jk���$�� 7������k���zi�~0��A��e���ǀ��y��5�f�~�Hn��0��Ǟcm:��"����a��5E�?`s���}y�Q�j���)��
���;��@�v�|[�1Ӯ�_e�'}��RU4���m��)m0�t��-� �j͐�Yn;��uD�I�O���
��f!C͝����u��\m97,�g��1�2m&������L��p���Tg��C[�*��H��6������/
ƀ�y+�͹�
��d�<�(��2k��	*�0*(��

B�j��M���gfciCk������#�z����"6�{�j���So::�.�Y��o����0+8�oẬ�Nz�YM�D�r�(��+k�����?��9�#�,t���.�
J�G��E�0"~�ƪ1�?���-�W7\�+�~>2~)JU��k<;��R*h%o���$�ơLΆ�ꁢ�(P@w'm?�մ^v���*1nܫW����_��׊�}��[��i�� {�Y�i���Ē;��Y��+|{�|c��l�0f���-�V��Vr��g*��F��J��~L�!�i�AE-�q/�o���jb|���zRV��ks��O��,��O�cؽ�"�6� �G�f�_� �<�Q����x��?m���1���crO��lK�5 N���^��6��*rԘat$`�_aP�	��E�$��@\����!NB�\y���&� +��Q�OV#�@�_!�T��#p��=O��%��)5�Y���p:�# ��?,�D�U@��]9+���P
Kid��z��˻¶��2V�'̢l��~?�&,������}��N]-��la#帆�q��A?	�E�T��%��!G,S�-���Ȥy����y���90��a7YS��rnC�����Y��qiE�b�!?�?��i����q`��(wCv6ٽ+�ޙ�Z��+=N�C���^e���J��fɛ�����랪�}�T� @���\��'q�\��	�7��	� �//w���F99�5�GS�����G#W��=�V���=ZgJ� l��Xa���8�E����_��Q9��TK�*�`G�0���8���(�R|�yhk��9
sׇ�sss�O{ьF��Yit��s%��h�HܷCo��J���*��yC8�nWޑ��훜v��i׋����!�%:@%r�w}�T;@�,�f>[��	GT��B�\u�v�I�'���Kih5do��+��`��@�mp���iC�I�;9n��^��7�$�4�RnS�)���=�T�e�r��Đ!xA0�O��6l����<���{���A,�_��Ӿ��L�����酰�8�dXȫv�9�ź��V����;Z�G�-K':���ÀLH�=����~�t�k�V���=0����%��3���=�����=⏩w��evH"è`�9����VKT���<�+���|y�k���+�/��g�@��f�ݭ<7��z�y1ׂ��Tw7`��t@�J�)�Ά��Od��z��n��WZ+�P�
�+��$��{�rs�f	]�	�P��a�&1���;�ku�	7æf����SZ�놀jf>�*�x 8��p|@����e�.�[y���-�,G@�M�8���i�IO�(�[�� �fA��),�!���F�k��4�
���AeM�1Q�1����B{�n�[���TD��9�i�"�П���%���mG����$Nz�(R�1E|��'Rix�4���'�!��=���+�Y��$�Z�yn?�G�ϭU`]e��� 7�yJYdi7eڽ����b�F�b�)V��o�����#?0+U�WR��I��-�ثG`���%���|��B�Nm�����I+���h�S���߮�܀�lt�fWٛo|>z3r���at��`���LI1J;aC�n*��ݜǳ�9��)��O�)���Fn^�1�'�U�獌��3��{B^�
���d�( �Ys ����%#��?p���{4V1�_��l!�B����}˧l֗ڧw�	;���C,Q��t1�W�/�!�?&(�
�J�zm�R*!m��#��,9�~���A�F��ԑ�{!�����y������5����3��,}���֑�kAL�=�uN{M��"��{�BH�1v�^?���P���Ô��&e�zq��q�Kpa��\���af�8
�|n�xhf.����hz�R�`5ZP��-�݉-��}�����P���}��2B�eʦ0����a
u]��Ş��꓈[�K��(��ƙ�� �)8a��������6�JNԫΨe^�ִ0IW�M\(t��{��j���FA�p|$�ʟ�S��ɮZ1U��4,��[#.��~��ȇ-vNGl�n|����#��'3�^h�O���
�{�@�������8��|�*m�%̄6Y�
5�������w'c��Sp&����fMPo�GX�Ɵ]+>B�8���M��)[.�M��~$%~�^���J@�7ǯ�!�؋/du����+G��t��Y�}���EB�~�����p0d#n@Vr��ˣe��~��x���n�,� iwQLe֕		��Q�dP����p���-�H�${ў��@|�u�Z��/�Ħy���+�������҄v�g��$��P���j^ Q�
���^���u�5����-w�#m?ه+G3D�P�	 ���R �]��VwN��Ł���.�T���|D5�_��wP=��l<��$R��E�9��+�w�`$6�ه�6�4� 4 X��뽃�0�:f��7'z���q0�~�2����~�1�)Ƃ��h=����Y�[xZ9�'�^��u�Ԝ|r0 &�y|�j6���S��hy����4�4xFlv+�������>	��Ͽ�Q!��2W��^Gb!�S!ӗ��|��o%��"�<>�YIA$��.�Ҟ\��,����4�&6������fsѸk�����]���u&XH�S���
�L�d��J3%�]
͆�ZHb<����;ͥ
�[)�ޔ�{Y�9|�_G��F�'����iy+ʥ�(�3���0�dO�WvS̀@jg��t "��Sv�~�g|�)���^q�Y'cj��,�������ݏCLO��f���M�|bO�D���ެ���+j}�ȟ��+�^�R6�*pb2H�P���Q�������F�@+��'=uA5�	�fK��zs�8	�i0�0/�3'�wl��վՋ�����!���(Ԉʑ��b_xG+���o�l�r�0Wt מ.ݠ�=���v�}��h�
 J�ܺ�����dX���-$�XQq�7SƆ�x2
���r��,����"O��:��?��N��a�mSF���i����ɖ�a#a�WQ��+�]���Ps��}^y�Q��B���᧕�$AlV[�}��r�<�.?�$�<�����*�!�E��0M��8��)��ٗ�4@G��6��B޿_W���~b�����3��gC�0 S�m���z�<�r�x1�� �vu#�$K�D�+Q,�^��`,@`��L��B2��ȓ5���?���N
S���cz#>,/��d����6;Rk�v�W��7��}6^ߧDu��6��x�n�bQCڥ��2i�%tfo�;�qW��%GM/�gQ��l��_P�++���YD(i�,3h���������+Q�k�	_�AJJi[�~fNc)і����Y�vi�VkɥSÉ�`|��"c�5�;QW���I����\��L�?oRB�x|�;��F�'����KCOjP�e{��D9o%��[jY�$����\���q��{�j�&6��04FI��Du7��W���.�9����z�2ڮ���i�@R�ekq�����t�ȹ��`L��I$@��9���B�ޙ�%$l�H?a�%�?�(��o�m�����K�s�M̗4�0a���}b��BJ�Z��E�I�$9	յ痸�Z��QM�����[tN�}�Z��/�F�C	«�7����K���G\���:f�����jv��V���U@l[�Z�������Xv6_MF��pGŀ�-WX�4�����Z��M�2�n��ה�����|B�[Y�v��w�]��¯���5����4�fPԛ �R���L���Y���<�'�|��~�,�]�5G�]��n�W�`���Ӡ-Ê�ɂ�J�w��J��r�G�|���ڙ/�W%����r��w@4�s�qI�"����!���S�
y�F �ԉ�=
���	-�Z��&8�98�{�����q��5��3�ZNa���~�k�;�2��4����)���+~�� /@y�^v��"�����%k��`ʕ�8�xD%-�����A�����6f,����#��I]F���F_	��w����_�8�j��L�4���n;_��%���9./g,��ST�_�j�j���9��L���OO	}7�-�u=W�h>$L����.}yT�/ᾱ2N>���K3�����t��y~B "Vz`U6ۈq�0��L��c�:��3��r�៹Ҫ�5%�7���*U�c��y�y�n�ej���ˡ�� � 0��(b�lw�nU��dԱO�[�G�${�� T��D��W���̦�fO�k��W�k��F��ܢ}����_�O���.�`piQ��;IYH��C��'z�{�1���[sDV�Z����p)3� ꧤ�Q
+nQ����D��[�h�oM� �X��3cZl�s��-�����V�)5�!������
��e<����&��a%t~"����4��[�>.א��Z�aeݱVg���o�.��s���eTs��2'��@��A��a���
Hx>�Ơ�CR�]�V(o������+��U��y Ӝkʂ�t,�̞B�������G�	qn^�9qr�$��B0$p��%q�\j�Qy��#�[�������Y�؛f�T��j}}P�Zh���$�N�Y����'l�'�m[I�0�����^�*)�r�ӕO[����A[H<��]������>���<}� Q	�m�C�zET�u"s[�^2��`�~�x�37�i&z%?:���.������8Y�z���q\��>�Ģ����/`��n���&�~�BJ2��؂4����t�^ޟ�&ZN?���p-�?y��o�U�5wX}��>s#̓\4�ܶ��;[�x�uH�@|�z�o�w�0����ߒ!M"~�� �c��Nc���t�a�n��ɀ�� �9�ٙ�s���xO:���Fz�� `t��J��)�H�=-�AE����[�B�7/����AopY���1�gɄ,�.��1�~��'(^�ٺ軺]�9� >&?��A"dz��/���q_��3كs�P&���:�=�BDw�_k���ll��ԯ�~Xf����6v�v�s0�\&�ԭy���oHᚯm�u���%��4���i����������m@ׅ0��nvy�*��}������_璋�N�B8�y2�tG�+���å��SZ��ڢ��E[O�ߎ�RYB:�0����2ʲ������2���;Z,{��!f�)�wP�E�n	]�۹�K]���8�K�f���X@��84���3YC�Ċ��:�4x��]��T�zL��ȩ.�آ�0&�U���&*�x����h��a�=:-�h���_�]eH�E�NЉ��|nн�hW�z��w'x$��5��Y����[��0��U{_���o�8o�}3t�p4O��o�p��х5�c8����>���F>�nwI�0ϰ�m�\/J��oU��OS��QW�YÆ{E���7zg�_]�@a��Xu;*ĄS][]��a�wo-�ch݃^�l�y�9+��\=�2Z�b�"^i��w:���	u��7t�U�i})}�W�x .@%3F�3���L��V��"�ܝ:ρ�f��&E��G�D�X�i��[���A�+#�� ���rȱW@6�CF����ˍUT�^��+_|�69��.z��|�Tr놈7���-"Wpt���}� []�I����Β����>��O/(1<���F�l�U�uN�.8���q�u�n����W�\�1��5hԈ���o�&|*�<�-~2dOM*���1����	����Ioq�J����3�*�Cb-�#w����A]s
�U���M�W���Un�7����5_?�I��l�q�yWas�"+�2oŎr���2w���?�X%��m����\5�k��y�V��L�#���)r�q޸Yw�aϫ�)��W@�[�"<�1w?�{&��c���lл�����``�cֶ\�G2<���Sy�,>�=D�S-�"kʐ1�pm��H��.'����.�h�^"A~�9��4\�~!��f�e���r���;��<����dSX@-���K##'�Sn���1�7���,��0��I���]�Ps9ܖnj���>��R�̛U�D�C�U�*�H�,xN��#�H�Y�jr-�(�(��"5�؟�2iq�y*�A~ނ]�7�7�L���L�}?Y��lF;�<5EP���x��
����Ęb�#�AV dpQ��i���?﹆��	��@�d�ot���t7�$�ձ�\F]~��Bs��g6�\�����Ȗ������L�^�?}q�<���(H������E?��N����H,�wQ�d�ٽ=����kSY-����6�|^;�� )�+B9��P٬H<��c����(�F@&	m�{���H�Y�K��V8Ҁ�4�3>��כ����W�H�Q��Ƶ�6�T��Ƴ��qzUW!���\�,��D�ΒګG�����%CS��~X����c�y����d�D�QV����`4$"ɬjz
��� ��Ez�:XWz��w:	��ߗY	3{=�{����Q����,�9&n'��Ě�v�H���&��/���MD�I��s
�Mńa�����./��`��A!Nef�GD' d�%X5)h~�s���^0�Qy�m<cmU�2y��,)fr�(�(�eE� DM"E	���6�F���*}{I˙@��zx3=&�8��}�7�#DC	%��;�F����K�/���6�z�xS�Z��!�:���v m�}L��Qp@J�s��� �.~�>9�kY�l�>�+܊XS�(Y�?�P��'眬�.�7u!��7&Y�ayRS�SIj|���&�AH�5lZ!y�p�:��~�bn�V��/�8�����v�ɊW�C�g�M'���o3�Q�h�|�U�Խư��T*P�����j 3Y�h���;?��S{���8�҆)�Skz�����b�0��{�V�X�A���?�ُz�����Ej�A`Ђt���GN��|c_�m!����x�V;a�^Fm=��q���98q{,u"���7���Z�[}#���ǡ���Se��2�����̑5S�����7H��7t�]�w�:���q�%a?@���~���W!��[�5�}#��D�0�L�͝Ԗi)�������plfȳ
�dk�e�֋�g��N7p�?M6��gY�����`�o�t�zQ��y�\ۨP��:jO;T�B�n������ķ�8e8}���K��{��G���ؚW�t쀭���_��p	
	6�������F��4TT,�d�ٚ�!�����	�/��"�dt�����OzOK�Y��Dױ�΃K�UnN�o��փdn�1�E/�^&j�vE �X���,h�+��
H��Q��FA��sB0�#{���g�V�~eϔh�3�N�(������Rke�6��MVhG?O�Mȷ��]�s��y�U1�iسqc�]�\Fm<���\L]�B�1�2d	�ٟA�ձ�����˛�`�ه�e�5@��o��~ԭ���f)Q��v�Tc�$`��_H���W�s�GG/\�J4�mpsL�:���q��{�[�|S��s���	���$�������KL���v7X�>+�Z�d�_A��Q�L���� ��x�D@&+?r"y��D5��&*�{Z���h�d�%�\O��r8�?B�u]M�z��҅��8u����D'<8�"-~�u>���(���.�xz?!�[�b9�����A$�XX'lF�C�/< �VS|��� n>E,�nJ�L����h^S\=��^���ϧ�{�ީ�+t����^8�xc��x�o���Fy!P\Nz	}���5�d���(�<����=�Y���U���g̊����Z��J��%��!���*���x���(@f��!V�c7��9CP'����љ���i��^��t�\��T�����;7�1��B�DU�T��>9~������J�0Fg�P'��vz���THvcx��J��)�qX^��QUn�E�*��8�n��Υ����/�I	�������#�tK�ȹ�WL7��ˍ}͇O�r.p�-�莅,�mp���A�j���γ��+|�Xl�����~���!62
Dqt��R�w�� �V�Vz($1SqT/,|%�c�T�.CY�:�L��+�N%V�����1g��{��h�����X)$U��keJ=�(��Gz����RP��bF�+MlcOH�[X<(��$���\�Q�e�}U�Na5�����=8�+���:U!����.@s����̓:�s7z���?����ږ��$oi�Z���uB���W�ȁ'�
�b@A���{������������[jԁ��ؕړ��m����lbw4�aN�C�6l*���
9Gv�����h^�m�B=�0�X�6��Z%J;pz+��A����G�r���z����8r����ɎOX(�\� 'x�9�����U�ZB	��#�G2V�Hb �x�	���_.,���k�0�D�ZK⪀���Kf�V8�?�e��T�݋2�fwI�x����|�A� Ϭ�U��I�e�|�A��*�,�e� ~w�)��o9��N��d���6X6Y�KA��7��$m�>C��C�]�Q�`	���L��vFX�@��e�_��	P��h����3�H ̘�40�}�ݿ
�.y�J��AphL�j l��xu��}#�T�u�3���+�����2�l��&�6�=���)������iQ�Qm�����O�A����a>������L�+1؆��4GW���:���>���%�56�J�hq���	�T50�U�;���h��`�X�hܗ�a6�ǖ�Ha�P��ƚ�,|�J~��8Wb�H�׃'xR���t�- ƫ��])�q��&m��J��cd�
�z2���]̎��Uhs���װC��ļ]�$���ٕ���6l�7��e�m?�e���}#{R�p~�x�N@V���*/5�Uγ�W�Yy�j��1Q�������^��ȷw�R?�v�r�!��Q��L��1h,�Vi�Q� Fɋsz��q@F�O�W�]0��6�K*���^iU[��Qd�A�ԥ���|�7��V�_�;n��
AC~�Ĉ=���Ҿ�cW	����|G���	�Lhw����X�6攫�����"�6{���v���� ��,+Ԣv�Eb��P�`�8bG[H�&\�����Xqn��o��Vep4z�<� x���Ǹ�J5U�*% d�C�E@�<�)�Q3H�S�`K� 0��� ��T���t�Yik����r=t+&�ZY⌖��D"��7��5ERD�!��b�̎\c��ؕw��3&3c��X~��:¹ڸx���[���3�kVa�ξ_N��Ju�Y�|�{yXd����A�+�?�,�pG�����*'��5[���
�kbXx��̖8v�)Q���j:�RG87� ��s/e}M
�p�:^��7�X;3~'x��Qn� �%{��dt:/�gO���
��T�K��N���1��Cm����h�U���#4�z�%�$~�R�kO��Lg^E�1`�8�h�J�O/+	x'p �k!^�VCs���=�V;u��ӟ$�1n<�&��s3�=ں�^{�Ym<\xۅJ��`��6A�g�U!\�J#�kl7>ſ�2�7���?�2�ݢ�`A�7S� �|�Yi'�ڣ���Shi{%,�Αr�ߋ,N��xи��-���9���Sh��]��3B�8��C�W���U0�s�v�P��6�r�	�eZ�y�.ɟ�a�����&��#Eڍ������u�#������\��|�&Pe=+�E���P��/P3�Zs�]�`HL�1�>i�$���hht��/�h�/�Fܜ�8���f�Y��L-,o�6\�nI������!i��s�hY�1ا��~�o>�����=Cv���뵶�wʯ��G~<�En�[�=OKn���!��z�- (z;�����)uD";�	:9����}6]���n!H':[��*��BN�ո��f�᜕�2\r|�#��,�ѥ��5�it����`��J"�3�y���8>H�e~���@!���#�|�q�t����eId�����~�$_�v��Vs�	�8�^c��FnXh�=4����ƭX�VU���,�w�\�	t��?=��%���|m`��L���w�t��P��n��g'�V��c��Vs��^+j��I��+)e���@�����w��h�QHUv����%���� 3�p��w1+u�~��Cz4]��׺�eY3`L�<�� ҺV��r�{Ro�����(��4�c:���K�#��w+9�="xp}����P,jt�7��!�31�	�����]�XCu\���½��K#'�F/�J]\�(S�w���.S�Z[ʤ�1�Z�GQ�\E�L;%���QU�9���AA`�����gȊf��
:��������5"`�U�І�N�'�s���:�-�;^��mW�r�����W�(E��?�[kxA/�����V��ެeP�5L�/��I�*�!9���:��_ _�Q��X�F4��%ş��	�B��� *�7�r�;��z�N���x��̻E���n�I��w��j��ɠ���W�M�TEm �DA���m������>��ŀ�]�8�!i�a���􈝛B��7X,��X.n�i~[�ce\F�����g�sEى��b���Fu�pkܥ��F*T[w�<*:�Q�V������� v��B�����H	<Nt֊N�@�$	*w��X1L� 0��*f��z�O'�>���G��0Ȯv����C��K��z�*!��%>.���:vP��V�� 
P��^Fr�A���R*�f�,m����h��r$j�G����JQp���4Ǧ�0�����(���T����Xwyh�~8���	�'TpJx��%z>3?�T��X	�)�\q�̬�_��k���
�����6�/�J|�n^~��ǭK��~���SXX摁R�I�O���O����H G�"��V��8�-���P��ƌI/+e�Dř���Qr�,)Y��Ɣ3+�Y�w�"�S�_g���KJ�=��k��WĢ`dI�� 	<XU�M"�7�^������.uN?[y}X�<���٬7&d[�-Ϝ�Mcxe4��k&��%�JV���S��&wxohiK�u�����1��!]M�՝Xy�,�F8D*��a#��Yx��@?"��Qz��6*����:G��r^2�����u�jZ��c��-Ӎ�ӡ�����c���[����N��'����*D�EA�����}�Y!���aAz�&1�\����7��hpgLR���͉�B\��a�D�,Ȕ������)SZR�~�b��<'Y%S��lM���jm+[S��w�|�o	t���,A�^�!�ڭh��[�"��t�b�Le��hk{o��ff?�%�f�U�Ix�$P%��0�����^�<�26�	մ��]qi;�I�J��6ZȄ`~{VY���o�,u%�C����{�1��Y���>PXS�h�d󤔀b���ܲ4Q	��>�����3�*:Ɔot�n�Q��4"�bw�~f���y#�e�j�
�E�:�����L�Q�H��Sz��R1f�l\�$}��|\�vy� s�2�M���Q�r*�o��>��BD�I@1�˽�B�0,���?�,w?V�/` ��ܪ,!Ó��-}Cg�]@��H�wN�NT1LZ`�V	�η�!m �o�{&,f^1�eO^�@$�CE�]����F�½\����1�(�$Ҧ��ms�(�Yd �A���O��\��Y~f�8qϊ��A�Z&��-<�� ���N�y��uL0_b�U�U�x���N����'�`�2�_�I�;�&���,و��P��SW
"��А"GY���x�j�_z�9+�w3�)x�y��k�.�&a�j�7f�X;6,ʅ+��t�goj�W�8�i�p>?b`?�@&�Is&+�e��;������{ӫ �T	!U�5Cú,�ʜ3�%���@0T��Ա~�s���|��%ﺔ�裲�0���vF!��6SNi)|{ku��.ݡ���W�"��(�|l��@���S;^o�A����f;�,���@b���j�i�M�`Mav��� �Ś��>5����=_\%��O�k�(���p�^d ���!�1I�pc4+AV��V.{?~0?!L������K0����ುX�{�p��E�̨��J<�W�!p����m�Q�:�߿42�@ܗ��e�ôY���S����
�DN@� Km� ����3)�:�����'ȓ�>O�u�/͇]���M�KC/LI@����U����䦒�ҟ���Ź��zx�1�m�h�S�ӴH�Ja"�J�W�@dso��cW���xw���{#"y�H��\3ר^������5Ѳ�d9��Ti��q="7�}3�9b>��.iH{+(s�,C�$cpp�X����Px��۵�J�����8X����9��k�~ma���\��-�������^rn�"J�֑��ƥX��;!��?].���.F�kf�ݸ��wV��ҁ����o�?jxP�%ä�-D�Cw#x�b����A��W�����,W� [����K~ߞ���C+�+␖�:
I����AzP:����n
�%=���6�Ә��k�`� �]�\J�/�<-s�U�SS$娕�Z ���q~ܝ� ��`��bl���������:�+�7_�G%�w�p
��֜S�^����鬸>�	wS��z�mߥ�����	�DE�ܐ/�S��0,	�c���r��68|ќ����t'�{�j�
���f�vg��z*˂����3�VB��p���Q j�z�#8�+Cl�̲�|����IS)�� D�K�Ҡ����9[C!�Z��
vtM��YU�dJ4.�%�A����u��V[`���)� >��C&�3N/~�zM��OG[��?����@D8�]����#Y<��ιw9\�̸�h}���Y\�Hx��o!��%a*F?�J�d�L��W������K�?a37��LIKO���OJ�ZM�[� ����ʩ�8UK_.�A��	G?����J@u��GU���K��3*ۺD6�.�j�����w2�L"3�bLcړ��r�}��G@jXo9pM[&�!i����� x�M��m�K-'cgJ�����E�[�kq$X��9Nu��UC .(�	���T�0��0��g;S�9|��E�QE�l�<�5�/*F��;��`�Ӡ=K��'�Z �MI�b�R.��1��X��1��!�WPK$8���x$��7�B nQLR�o�4�A\\�����w���GJ���t��^�e}�X�9h�D�/�.3 l~ɀ���B6���B�fE�'o똶>��cH=5�-��Z�A�HL����!��(d�����C���t:�l�Ck�l��C�
�+'AAJ��`����Mj0�&�=N &Fx��@�a�M��ٙ�?٬=�erV��i#���(>iE|��%�/��j��6?6/ɯ{�zx1Zŷ���ܶk>�@��{
��;����z���A�*�W췿��D;�X��P>��Y��Qu ��-�cz�;;n��{�WzZ	�.>�w��(��cL\e�.,��I١7G}�fj��_�I�������_��$�8eV)*�����g�h�G�L63{|�N��~v1�Y�I�;8q�bq��ʁc�z�s:ml{b:��8	j�����Q�Q�]�G�aӊO�$J���*1 -� ��F��b8�����ꑶT���Ƌ�-��K����D��v6!�|�ǲo�L��7˲0�۪�n�^��=��Q�$��.����菎ir�]���.q��NnK�S�2�meꨟ\ʗLX;)Y�Hb;G���|�8�a�8��\���z��=>����F�.�Vch3��A:0�Ht�=�s��eSA���I�=��H�aI�9���a����c��N?{#�_F�+3e2{��P������7�^W�p�5����������F+M�ק�XiG#��{a 2jp;�0XE`W�������C�LS�й]�h�r���X3�F"9�1�#F%$��(Y�#�V�AK.<�ޝ��t$b�llO�ن����4,���]�~2�NBF��bd��^՞�zf'�R4�(��|����.U�7̛�zH%�*m�����@%Y�n���~8�Ё";��0@�y!���%ŝ�]-"�s.j%�\�
�M��C|ǫUHP���ΛȄ������4���jUI͖���i-�Bm�C4H7d��(����8�K:��;��y��V�c�B���M�2z��g>�!�sw��#��Znq&,����p 0���2�3�p����gd9z�3�a[z�&����X$!��۫ ���h.ԓ\�
"�Cn��/s�;3���VQ����< S+�`C�/��Gà?�ҝ�N�}?H�B.p����*I�r>6j
��WI�� [���~x���Ο9+��R�����c#���↿�z�Y�D'��R���"q�� ��=+80�/{1�M�)w��.��,�a��0A�@i'����.�!�Ć�����++��s��la�����	�LߦflZ]�·X��}3T���bp�U��[���M�p�Ŧ�|?� ��m�)�>�Զ�}˞;�ߠ��8j��,�����'`�����#G?mZ�l:��~{Q��B��� TWe�\���N^�R;�]���`t�PLB����"��D	�t;�.�B��	1[m�t��Q�2��K�ٮ�_s~�?fO�P7�R
�ÞL=!Z��AWS��:��7�.bғ;�B8s+��$vcE�-y)î�wb����q��9����6�=�P��&�1��!m7������H �����$1��5�B BY���fB�3�N���]�.jl�z�t��Eq>�"*;uE�(H�I��*Y L��̯9����I���/n5�6�s�-����I��p#c-[&_7_����K�QY͓�K�!ex���ЇYO��yJ�~���`�cg��Q�j|5����ԡ�Ly翹�W֞�#W�>%���[¤����c�f��㶷�w�0|k��6���m�%^���%�h%�#�4��p�W	a���~���1;�U�`s2'�z�M*��67���j;-�t���T$�=]h`v�G�Td���3�1O����Jr��~WZ)�9��#��S��� �օCSf��~A�7`=�3#%f�gcp����v8��"���%��A�E�(u�!�d&�������H����	U�(�r�<�#�.,y�}�J�������f"�oc��)���N~������E��B��$
B�P뵓L��.����j��6�Ѱ�7kHU�'�S��c��Yy��n��S['�Gy,N��Ck�p������<k)�0�o�|���QgU_
����9C��I53GWLI�؛�|�2��\�G�BMa�G�Q�\��C}�+N=�iu�&�u��=FS���7+K�0.�0E1+���-b͘���]$a+�z:�®��J"���ll\%d� ���C��N��~�Փ}�V��{��Ê� ���Kc� Le��ī����U�@NLI�P<���L������A!���r�t���vu���K5�J�PKӵ|�.�2�吷��V��B4c�R_F�	"i,�>x�.���iȁ��X��V",��7L�U����V����  OT�{�q#4�/tK�d?�Æ�;��9����R��[��Gy!�۝7�d��z9�?�X]��/}o5�E���C�M�_Ա��P����f/ A{]MyJ�ˏ��Ƒ8sI��~�^v���R_�J��	<=ia��;3s6?�}0^r�3,"6���P�����,��J�e��Ә\�rWd�<�{
�A�p�}��h	&և��A�82R�q2��Ԥ]�����>�Cޘ��T�7��.�hB_��%��Dh�R��WB�Z;��g��5�7��o�b��Vp��'r8Rhpb@�Y�nK����{8���H����:k��u�H{:S��	��"��)����,B;bE,V��,0�}҃��!�=?9;]�h�ϺE�f�}X��f��S\�,����G1��� \I'�?T��ׇ�Q�! ��FyJdֲ}O �HI0����mx�-\c2���B'������
ܿ����"�-�zU:��n;��e�>D�!�C�.�a		��G�w a�F���@��I�N܈�����Z=������W?���S�*�x��C���k�����H�ђ����C#������� ����,��DvU��kI^�1�y��;�gR�n����~]Ţ��q}�q����MJn.^��t2�ڎ�����3�^��J�<�����Ɵq!=�Rǽ��|���х9�a<SX4�c֌8�Ұb�@�4W�y��c�µV�(�}�^�<��Q��dQ�n��{i���9��ͻ5�#0t'(��'�%"�$5`BS�/T懓U�������X�Vu׋��z��]J��K��C��"A/�A�kX���ci���m"�-b���':U�&68$^E������;��8n��G�t\>�3. �;�4u��cV^]W��S;��c����j�c��.i�3�|i��'{�)y�ߒ<gu��2s>�p��h����9'CBA�5�x��e,��r�*�N�����^b�c��JW��=zf���ɿYٔ�)�����k��f;cw��Q3 ��8��8������[3[+�E�Fx\r��g<~��X�Z{����B޺\���x,�'ͼ}�k&�􇷃e����P"r�<̮��l� �\iS4�ƅN,T�+R���\*�'%���s�~{����	2B���|��O�*ӓ
�vҾ�8�� �^ϕ�퓹����R���U;9%�&!�Ӊ2�iy���f����,m����xS��I�g�-����WC7߮8sx����/:��*�z�:����8d���X(����he(ô;ǚkb!���j�_�=hX�i9���+ۄb�܀�@�j�
�k1Jo��K�_%Z��_���C�].�)�]����Q^�>
�.�GW'��"���]޿�U} �C����3MW<6�&��e���5M7h��!���ǻ����ժYH�BNߝ�
;y=�1�:�)��yf�]me)�E�=�o��	+D}ѯ}�3Ī_ �k����O�l��CD�rsUͥ�-n�|�R��L������6h%��!���� j��R� 2�3�:t7���9�h��Մq�M��:N}��o� ҈g�_�p���>��u{��9���LL��������f��"!��J��78��&���4�';/>�QL
!Y���Y	�g��Q-�휰��#)����������.[���v�%�+AŏG��>�b��^��	Z1����h��XG�G�F����+�z���NR�8U�3u)�/�����9�
�JL�tQ��7V����p�]�f���o��@�v�������6.Q�� Q�ڑϯ>��;	�(B��`�o�N�|�ci��Ѹr�W�Z)���ߤ����h�}&���1#�u�?9��-����ٓ��>����E=9kf%���p�iU���]_�'�1�h<���;��(s�*���\��Q��+���~�O��#y��M`98�a���T4�u�VEa�` ��_y��UN�-���'H����m!=yi�ӑ<�T�`c/�,4Ӥc����F嵍��$��Q�=�g;ȿ�ڤ���� wWص�G�q����� \{�^[B���21���,IV���Rn�%���+B�`
,,Ʊ5(��	�.>���aϐ˪��O¬)��:�ZH)����8En������yQI��"��_��^� �;����"���$�U�z��W*�ӣ��0��l=��f���W����L{zXZߖ�����=0ͻ��:��	��,�ߜ�Λ��Tt�M�I2��Elc�ô�Þ�ۑEE��}�A��A3����Q��ȡ���Ύ��M'7���ᓍH�����S���:sAhڞ�5�Msb͐,\'�E�9���Ĉ�y�����Ycz4�Ц�=���ߍ�1ԻS��,��A�^]�@�����z	4lл��b{��SKN[d�ů_�x��}4�]��ܐz�z&�N�?=Dӏ��\����&�JYs@?$ĥV�8�M����]�xhSK�{��$6����9�#���joP���uU�9��5�;����^� щϾ
;�{�Ĳ/�;�AI���.)y�;y`��:��mLbaL~�J0��K4%N��%sX/�]Bܶ�.
h����mfJ�u��Y8�[��� �B6c��2:�w�v�x�ZKb<�K�f[(���>3�׫��3#��4��U	�'s�,a�`޽�͜��y�,D���22�K���Zs�<1����ǞB�'��3B�� .��k��l�F`�+���}��x��W�η13�դ������\F��V
lZ���Jp+��_h�ѓ�q���@I��)?��o�ziA�E���U�N)��0�)�1ʹ�f8��g��l��6���� :ʴkخ�͇9�X�	���ʬ֧q�;C鍡��~���r*�W�@��V����]�m��_�8@^K&�MXE"��]���.0J��0��@�Z�߫ь�/�#��J�E���� �yBN�j��"��|}��p�ߞ�L�����H$�{�L�����������X[Ԏߙ���]B��.�T���9]�$��Uе_����K�	�g���B��c>�6���PR�d<3��;��]�ɢ��a��v.(�h��j��Yg��w��84�I�S���Fd��b����G��溡��K��.�YDz��{��z^	�F3`�όɥ�8i��JO��5��,�D�Lq�����뚆VI�>`瀼��0�xC~}$��[S!�"[t�(jR�j%�a�N����\%�i��dGFS�\������Nxu�X�����ge."�3�%�Q��	pQ�`���x	�#1C��e�t�OQP��z3���=g��*Yҿ���!H�'��;��h��V�cQ>�YIN,:�\:0��z7���vz�R-�*$�!���O#3��i|:!�O������X*�D����t(�����'�?b���^o3��gܾ��]��5�Fb�4��
3���f-��J��	���tG����J��;i?/�o��c*�����d�<eҴ}��;0�J���<�T�+k%8
sm�������By1���8J���ݎ����[Y������X �(�Y��*�y@T�5nq[0�U
��:�ʩ�.��Ϊ�si���Ay�J��r`�����\�=��P��w$떳�=��X�Wr�������-��2��d<26	�U��(��A��Q)3��x�3�2�+�W���^y�WŌ���W^���_�@7{�y��H�%͒Q#�8����"�ܱ���'ʞ����H��>#|����^�2�'bְsl�_P�w�&v��y��i`T����[�W�?~����l�&�����A�ܷ'�Ek�e�T����Z	��B�nG���[!�Ŵ�!_ʭ�W�3f��Ώ�p�`Ҁ�����@IXDe�W������4N��C]Ҽ�_�{�W
_��A��M�W����!�S�)Vw@��zU�MT'X�Li�W���j��u i��N����h���E4D�_B��7�
����W����dZ�o��X�������0����gC�Q"#Iĺ=�n�����{ �G�~�r�D1@��(f�������:������2;�l�ˣ���b	���z�=�`\Ђ�8I���3��ӭ�y-9E'��]��c~�8��K����b�X^dZ���L�"��"$���!��:Sfr�"|���(`��Ě�OdRʝ?!��E�����:˂96��_=y.h�c��ؖcM�Hp�<�r�ހD-�<��ȇXX��7�a{���Р���7�x>�����MH��u���kV�0N��C"�Y�Y�dAX>y�������ݶ���5'+�ewsߴ\�L�.��H􃉂!<d<X��RL�J�n?c�-�r�V�3Z��s4\�?�;$>�8��d���!��$ڢ���������kg\��~Z���P�̓�H6"����~j�bټs! WϪDŴ����׬���@S���H�t��,�����JD�n�U��	�	��6$�0ܚh[����b�����+����8��0Mi *酰���N�~+;��W�m��P繧N����3���A���z-ݷ�}�s�%O����eH�t�>�WL���^�7m/��p��y�'Vf�l(�t��(�&/A�pJ�]D1���~r��?P�8 <|#K�ܗb4�?�Lɳ`w��1�5��4�ib�_-N���?�ϓ-w���)'0��k��{A��b��~�?���]��
��Vd�n3���i�k�+Y�t��dif�k�n���C���5H}�/�JR��^��3XqI8�&/�=޸��Ω����z�jYO��r_[���xRE��Q��0�Y�BvB���$.�m�ϭ��/V���ï���_=�Eä���ʡ�u���S���ڔ����Ů�c��5�2�Q��(�n��#��D^����!%���A+@���_������Hr,w����n���!'������������xl��
O��P|�9:�ߵ<����*���'{I<
��^��������0�I��
 a�5��O����Az���ے���������[���ܧ㝳\����(��%Ķ�R�>���m�E:�2Φ�}���!|� ����k�{���'��-c��\o�Ў�:c�V�x�o�q#bK{���.�y2�ہc�9�?�#x��~ͲǍ�;4�^���D^hI|�����V9�B�0C��DO��]u�r����H�m���#��;�.��u�_D?��$ %�;�pz`�b�3i	)[�oW�E6j���ա��Y>��ɩ q��y|I3qDfY�M�J��N�PF�v/րU��B��s��~��R�	�7�ʬ�SOp]��?���>�/;�2�U�)/����'rr�X��z�&`�{���N�% �o)h���-0ݡ�;���X��v�b;:u���fلj�Ւ��T��\�Xm�K�b�ο�ɺ����Fb��^UN{���x�#a7�YsuzN0UtHGQ=6��R< /s��k�K��űZG;%x�ܣ���=���J,��]��6,M�'1���-��\P<w�g��G��y�S��s>+����%a0z� >�	�5���ٞPt^���6�hc��i(2!��t�:|��h�f������Z��Jhw��"b�[����#��7<��fDt��xL��S�lƘ =*^��Z�g���G
�GD?m��>:tf��l2A a�~�Thi�AB�	��;�l�g�=G�(�H��^�	G�H(������FL*�J�j0��ǔ`��lR��3�w�S�6Q�+��a�6�Mi�n�.ډ�U��tt�	5��������=�!^��������r=��b0��NBן��<�-�8��㮒]��,.�hb�i��uJ���jvOi-���XfM]�Q���{��E��q 5�Z[:���L�z���s�OdK ����A>�t�q2b!M��G�X������D�(H���O�_���-���	g��h�x-㥃F=YU#�oBv��^@��� ��2�g�S���9�<�����uŪ��xiS�3�)nTdq���}�qIH����O�-��mƺ�vk��Ĵ߯�c���cbv���K���C��j�� 7O���ܺn-E��ќ
Wǋ+t��ݷ�B}'��f��:�ߕ��[�rp�����\�dz@�9�C�A�/0�f���־�z}�:���H�5�4D�j����qg
�so�M�^���L����8��R䝡D�t�dg�YN��kh�TJ�.4�k�<0�|�9xȌX{>��G��ϭT�q��4R�!�E���
l�J�0֓1߫.�]�)TR��ڸ�-�$i��a�T���'��֧��tp.>�
CdX}��s�w�����g$k������"ӟ]"����N�H��Ft@�������]�s�� ):]�nm.%Q�Oj�0�7��A��@ɩdq�h{�+�Hf�\��l6>6" �ձ��D��@2�J�dg<�B�f�5������}����M$���˗Q$g�uJ��ׁ�&�)��YA�,v���KD�v�&��	ڶ�����p@l��W��z�4x�'+@}
x�$~���'%��,0#֓t;�[�Uu �mG8H�%���(B6�oO�'4��e$�q��r˽Vj5��^�fX��,
n�����Sy�9�F��]�24� 2��� )�$c���0X��s����^w�"��3��x�)&=I�)��c� C`��aM��4Ns����j�V�ħy2G��?r�\�5��%z0~,�W��
W�Ҝ�5�˪�Ԃ�`�R���)ƣ_��>��W<��J3)+��z��T�2�N���K2Cʷ�{*�=ִ���� S�;���X�#uQ�G�� ��i��_�����(G����
��4]��H��������7���m�#� ��UP|)��C��@�&��sj�F^/�:r���[�p�x���|R�ۋ��h$ZA���bu1$E�^x���SϠثXa 0E�k��i]k���7���s�M'mz���H�,�~��sb��ϚE�>���M޶G�]�y_z�ރF�r��G�����l�R��G�ӢQ��'m��ot�,X��)�7��S� ��[�H�뜙ﱋ�����~�y<�B�(�X��"�@�ǝ�O�ϕ�\�������8�и�?}e�3/�Q��=X������֥՗.q���x��n��9�/��vHi������݉��mt1�N��RE��Oɓ��u�y�Ƈ�tBD���J����d�5R��y��OL�m�{���P��W��ۚ?Ew��b�R�ƌq�9l�$j���B�<C
.5�@az/����=�ܖ�W�j*^��,��@��b��K�iG�����b �Ƌ�3��s3M3�#@2�G�EK��H����3$J��3K�8	z8�w�^;{h4���9����>7\���)䩽�p��g�F;l�_~�,�(ʜ1WD��D$$`ܛ%�0��C�Ap����0���+c��<J�~�]�{�[$���`z}��������[�ؽ�oRl���U`�ea7�`�3���
HC�O��U*q�
6F���q)�f��I�2QY`�S uYP�\�sBw�)nts��ّ#ii��;�@G�ܟ�w�Zv��|��'�SS�o����<�8!Lr�����ۜ����4���	���.��Z��K�@Q�Y��O���Ҭ]7��=���Jd���ǘH�H�m��3�����	��0��.;�a�2楂*��y/f��B���̎/i^B�ḣ�h��,���(i��6���|�]Y�C�ͭ߶0E/i0�#\}���(.пU����aw9�
ۺ���9UA�^F�7G��nm�_�}b1u�24����"�_X�'
Igj��N�)g��L�Q�+���隇4�#����H��,
������f����99�̾�{]����]�oAF��1P ����i|����`')��L��#�s:Οa%�Pc��O�F��0Q���2"��'��l�����5W��0x�b��9L3Z?,Vorh���D
���b�.�:{؇nY>�����V�n��,f����Iᇲ�X�j��L�o\�/3���	V�zۃey+�U/M$E��b��4��Ò.���T�P�ö�i�v�;�4���[0�3���̭+D��k�R_mdK'\t�B���^A�w�����jr����(��SW~׳��^�{D_�&��ӗe��x�͋��SV��}V|��� >�( �y|�]n�p���n��;��ܪ�᫫'�t��%ł:g �S�}gX�-F�F�X#&�ʵ���	
���;1�����@mZ�yA���P�|�2��bSg���l���>j�tà��E�#�
J�z~
p���5	���"ۮ��+�����f"δV��#�$�zP��͘y[�y�t�F/8mv@�NA�z���9_��D�ɕ�ᯍ�%����]�d�e�߭�}�����,v�l<�\�Կ>���h�Ff�i��;p�Y�M�ӽZ�O2{x����nʤ��F#���0Ũ��dT\n�yF9�cd�.׭���콀xNAyv^`%o+^�g@c��ɓ�v0�FkGd�[�nzs7"\�8uѿ�'��,��F@s�6���e4��9>�UeJ[E�J���[B,���:{5w���E�^-��%!��{�6�\��1��7�+��$1Q��N��!�F�+! x�%T(�(d4$_#�U�����ܬlx��c��bAT�4�x���MItM�'�d�/j���匧��D�x�9�F����tM�=�����_Ӿ����������AӨ�������n�jP�W��=$6hg�P�=QM��L��^���Z�oOs%c�������я�Z���<q���ߋ:���镋[�q�>^��:�_����)�B0�V��R!�1)H�t�j��^$��6^�Z��y�:��nB#Dg��F��b����˲��1���o�-�6i�~����9Z�+�A�5�$��U�}�XWQ��!���ū(��ˍ�I�x��_�Z'�t��5�7I3Kg�_�I8ʑ=Ч��c&Yg�(_�j�1�a��ħ�'��Z"w~����)� �,o�p}�.H_r2'��o��e�dny	�������y��̨l�L�TԳ��ԡm�Dn���@m��c.m2eO���N�c��r�#������6����߂Bx̴��gb����UI��n����C�oxb.�j~��
�m�gU>�[_�>������jU/�9����1���JbX��V���Q���!Nû$+�h���C�cg0ʠxC�BY��	�����k� �z�a��ċk�s}1uS Q�]*c
6�N����Ǒ��m��QQ]�ѹ��_n�E�]� c��#Cpv_�]�̧�R� r�ʼ[�pF����O�3=O���75����sb��߄�m�'*m�k����Y���i�a+��Xk���w1��sV9>->���o�0M�a�G:hٳ��W�F�\�s���U����'�V�����"C���'@ �|����K�*L�A�x������5�B9VE��	�>�fV6p%���<�1=�!dRNI�_�$���X&S��D�!�m�<�h4JBv�����Nqs8�.	uv(5a��u��`ةGƬ��g��-���k�Q��/�fgz�,����ܨ+� 7��U�p3p2S|{��n�pס����L��w�a<p{ǶP��.�H�e�<����_�K�p�sg���|r�Ky�Ȯ��9�K�Ь�-�Z{ ��D��2�4H��t�`*O��5<��5 )�r�u�EP4��ik~���@�����C�gV��o�Dc�����d�R��T8E�'�g����oJ������W\��A��2��a�e��wû�6P�| M�պ 4ǬY/ɸ�t����A��	��DR��F���#N���x�4��U$d?�E͕��d���[�V�)%�&�W�4�L��6�YӁ�3��;9���W�r{�I{��e�y�ca���2�:�I�Y��è���x�\rJ䥅8�_�.uq�x0���(\Ι������Ԑ1���+[��\+���w�A���Urӣ4��n�)�|}�1�s��G-˳���.�鞜A�"7>]��BV36ObMVo�c6X�a�*F�C��}�2pY)Q��ꦪ,�u�z��c��PpWĭp����Kq '�_�E?O����Ć2˲��{+.o���0��X��mN����%�>җ�Æʳ���#�^%b3)����B�d�i�6�p]'}',\9X�R!����W����i�J��vBE�������[�c��`��8w�Fs��د��dG
eZ�Q��ԟʹ�tG�&����ń*-���5E��8�
��1Ӳz'���mnu�4`Qb0�|��
KZsᗷE�҈�'�����9W���1��e���W}�7����8�K�.����m����cF��~��֤�����'�}�.�Q�7�������vԝ�s?B�\�d�קL��~_�*�A?��F�(~(��TS�^hI1e�b�p�^i��ܰ�JЭ,�ΨV��m7vb|4�t%D�|T���b��;"�����~��Ӻ��h��;�*
�'�I����� m��L7D�j�t�'������\�]���٘��L�#`�
�vw�&Ÿ����"rO��"�B�홋V�H�����_�d��|�y_��2C�;��}�� C��� `���q�x�g�\��H�'�T_�)n�I�\)d,ʹg����Y��We
ːs�|:;�sSq��%B��������d]�޴K6��c��	:�ߌ�=��aM��{�t	:"NX%\�$%�*Bu�Uـ��P��ָ�^�)6MJ�ބ�q��ӅX���� �� ��� �5yȺMi֑�p������-r65�\?W��;r
��Ɂ3�87E*u�"ꔅ�¾�� �<>ȯK���K���%����`��&2���4$���N�0B%;��Oc!$���7܌�QdW���d���1�C��ۈy���wM�;��a򯵼\e.bZ��~Jey���{��f��Y�D�1�X
3�B�&.��w�{�D�ʩ��I�Gi=ؓ�৴J"?.�>��O�UҘA�v?r����8�^
�Q~�ͯ�C[���1�g�]oE��}�ё�5M�M�	�v[�b��sp�E��m,L ~� �k��B�n�X"N�O�COYo�Gi���u]����z���mk�m�Ǜ���Qw��B���C��6��Q�
K����d}��$޳�};������.U��2��E5}u�`1G�?��O�������vG&%q����dZ�7F���$bYkmBJ��,�O����l�;nn|	a���xj��H�0�ÇG�Eќ�<���,���ۼvk� ��G�����eģf�Ɩ��*5^|
mS"�cɾ���}���(K�2G:��o�U
�3_8~���ڊ����(�>�@e�q��t=��|�5�k��R��Ţ)S?����M��,��N�2������Tط�l����[�+�'�1�u�r"���.���W��d�R]|','H��! B���.�D�L�-�
K�J�5e~��n�Ӣ�e��l���Ȅ4ؕ-�;��e������H��~S��7�9�r�a�y	1�؉�������M�I�������E��l��cf�Hk������=L�����ueHG4��_��J^C(��'���k����[�f���);�y�#���i�����	�W��u���=��}��VJ@�� ���k��7q�S��-��[�c�M�d��
D 9�0�����%i[�|L9?"ScW�9BěSƗ��
��b�����Ҿacx���')��B\Q$��<9>�ٿ=�:���7��"\��1լ�e�Q�t�@��I���<
�P��V �OlK�|Ǝ��0F� q�1�b>�'�;�G�u�� �j�t6�3�t�tC3>Yh�Dr'����Z "�h[X[��@q*��>�ýQ�Zr`��u.X�voR4�vwݕӨl�7�zI��B3�1�Y�_��:)�ȁ;��\~�V��"��oRNQ��������Va��ׇ>��vH��A�(��Ѻ�AVb
���K���fʞ.��omv�U�Ynf-�;?KH�?}������4;�ܙ��1c<큟�s�w�@8����"�V�)���JYӁO2<�8`[�3|������]=��@�|�����;DԸ}���1��ͫ���fZu��Lv��A=�C��j�0�$�����tW�+�a�Z�e��[��`_٩AX;F�̏;�(��ڭ�~�%O�ma$��~�
V&��"�#cٳ�j䩋e#-���B�Il��,"�f}��?��ݤbY���sr'}U�%�>rɒ��5@�SG�?��i|�85���\eGG�{6$"�vY�#�t��o7#Gn��b�!�S$�Ż�L�x��tS�7����.�Ϲ6��ь��ct��Z��>�)��d"@!��N?=r��ԅ@&�=���^GX�~�z��� !����!Ղ\�v���O=���Q�\���䀢Bȼ�9l9|E��낖����<Z�CT�8�Ɋ��-�'\�k��Xp�*N`|�n�n0���0�Q�7������9�帝<�}W�� (��.�er����U��	b�)����t����B���P�k���QxL�տ?r�:ʋ��tbVI,��S��B�t��&e!L��Fh��QO��B�E0�� Z5�;��#�ߍMX���Qh0�����e��Mee�,�8�̱+���Ҿ��E���v�@��a�9�$ ��=�L�+�] l���e�
jMW���6F�+,����uE�tS�)
�
�Ax$����p'pl5�eY7L@8k�eJ蕄6�	���.�%a�cV���U���9����3�S�Ϊ�P5���:W��C�@1{���0cd�g%���ǹ��J�Oۛic���u'\� ���2w{c{u��Μ��gUf����o(9зcUhf�Cr^����9�f4G���|``^'������Ia�3�T�,L��D����׮�C����;�y��"�*�Yo�DM_�D�E(0�o�gJ�"��鬄v����F���8L_�H�Z�["�u�'H|�k�i�X^#�A���r�7dF]��>����t����j	�ȐyOjS��ėa�pPC��>��J6�4�VZ�!�SC{J�����Ѻ��T8߃�1�/cE/��V�OЕ�7[��o��"¦��}�Ct8�m �.���FR�	�0FK\�6��4���w����5�`o��}�M�g[����!����!��O�p~�E.�	�Z�-j��:�W~R��>���o��X�1@��0�_�#��d��Q(H�a��:��:�BZ�|Kk�md"Ϻ��4�g�y]�9��P�gx�aK�**?�d���2��(AuK��3T/g�3~&��./� �C-��C�9���W��=����ܟ�1:�h뚑\�*�磛��U�K1C7K3�}�Ѿ?h�:U��堵�I�.�	�%��bT�h���1^�>���<$9�s���ĠS8�����~ߠ�x��1'e��v�ܩ��A���L��*����V�ע����3��ǝ`�[ǉ7S����;�A��꛿���ժ%L��:�>'����
��Ƌ?W�;�2ʯ8��T�$�a��tp�;%��R�嶊�R�
U]�>	���Uu�+*%�I�4]�$��)�|�:9\'�ۧD�c�����	j�d�}~`��f�Q��t�I�.ǧ3��!T�.�,���M�������60iu�U���1�~�*�Uw�M;-��F�%~�ԺB��w"�A&>�Ӝ4�T�35a��>�٬��o ��곤h6���|Ө����Ѫ��e���HKl��9�7r��s�Z�뜌��� ����e�7�#�\�+6ٻ����ĥ\�MʙF�Q?Hh���"�E>��g�V�4��v6���g�U�!T6���b���4���N� )99�F��md��\�/\��yG۫n�c���A�8�d�� �;��y�L����5�$:�#IH.�� L�(i���Hji��*Z2$ݦ�Jlt�F�
�wC�� p������ٽPni���3��4O����w�%Kgl[�b�WZ@��L =�J�p��6l�〵���7���?h�f��9R���qT-���|݉Z����Ͷ@������x��?]���:R+�I2��:&횜�L2���=�l��32'I�#��d�Hk�����I9T�&�Vg~2��Q�.LU^�`� �:��6�;F�d��r6�K�^ɦG�?����-�����:_~�?�5娥:��Z����z#�=R���w|�@L��DKSa���:#S��E\��y,��4���k&w}��.��R���FM.Su%i7�������X��e�S�~�����?S�|6M'm��r���pJYLpb;��00�v9]��FO���Oa](Az���4��=s�(sO�&zK�X�z��59�?��Y�7]OR6�U[~��`���t.�{m�rD�qm��ί�)�=���(i��W���C�td!
���~�b����B֜�.����U�y��BmU��2<b�x��5�0O��[NE���1�ӎD��2��b6)�Sm��PTUq��/@4�dq�>&���W�\�:�O���1u̱^f�w(ZP1fto�e�pjw�K`�a4�K���!�*�/�,�4u:�R�� �H,�cH��Y��6���{N��^��LxA��R(�>W!5*���XA�bYƯ^�J���RԜ���hx�����z�4Z�C�Ȭ�E�n�C��F����ke�Wв\JY��j��Y`��s�*A�Da������3u�:�h>�!ӟǭ��+�f��~!0��Z�{�rc
���]E&�DEA
/'M��.����o,���G�x�uV���%o���q'艱M�f6D��f�Ti},�>G�VM�i�P [DB{<`��"��UJ	ق��64a�`-r&���!�QV�2pC$�B���W�>�I��Ȁ�4A�Ŭ��Ba��e�ie+�it]�;�XK�$4�}s��u�k��Uz�4��dk�]���D(��-b��q'�>ן�G5��7����R�*���޷2����Aú�1;w2V�*�}�JSCpmi޷ �.Ҕ����ߜx���*z
}iV�@[�L^*_��~�0�nF�'�M��G��ѿ]m��N�����#�b/�y{h!��*"5�Gt�d.\	��ٲ��jM��M(w�+�y�����I���Md���
Xq���5Q �_ ��њ�Ț�[q��$�Y������P�42������yu.�ڑ��C I5�1�*��}~	tQ����=��;�7:��.s#2��I)��/�vT��[^A��u�W=��z~�O&�961��O��P���	���A��t���e ��LM�����Zې�_ѻ(˒��*Τ���/���=Y�.[d;���Ԑ�p^�����{$�v�8fĔ�W�O$1qOU#��6�<�,3�!7n��\�_�JU�Y��×����(�>f�yP!&vUd��ύ�|���~�c#��Tq��}�Jf��N׭k�f�P�0���fbrH���[B�-�i	�c@����u��Gf��̓e��?w60��(�w�G�������%�9�C�h�wu0?�0D�'�̨6|<�
G��I�$]�Ϭ�wt�Wvf��}O5�E_���9R�ډ�·�n�s��p[��� <u��G�*�=�2���)9�ÛK��h%{M7C�$���XI,X<U{P!�),�кP�"@ͣ�%��/�:&�E����Y���j���;���%�v�/�ߍ.�$|�ռ"���C�; T9�+Ƴ����D%�ε�MN1�m��w�񗘼��ⰺ�D��m�[�;aE�K��C>0-$��C5b���P������i`-a�㰉�$\P�a$yI1s�.���s��{"i/`� �]���/A�R*�_���(�����������#��j�T$/����r%;7Ō�� �8�6=a_� 9��u�^��:�5��j���<���'Ӭ�rwz�m��[c<��`��Ynq��v1C����a}��N|?�� ���c;T�{;��H?��䒻b*`u�W�毓�N�G]R�t���e@�b����]ds�nnJBw�E3�?uB˖ŪU��6]�FЄ$Ma�;w�2e�,��],�o��kc_+��X?u�72�R8���ΰ�p��K��/�ݺ�`�`����
�Y����
{�p
��Y��@U���17���Ly�/k� ��y���}�ĳ�l�?�����ƥ���p�ܶ����ΒZ���E���K?�}⺝��k����W�h��,:��1T�"�QB�6K�����`ț>�YB��ǀc1�#l�b~�~��������v�2O��Ӎ���ZVŝ1�@7�k-zכ�RlHC���f	e��"�oI肖ȿ�Ԛ+��yRzz��q����4�(��1�t�%�D��2�챸�о���㑋�(;7�7N��\���wǏ��f2%�V}n�;_3�hL�����fxxl=��y�k�<���is��Vb�YGΈ�g��I1��l����]���v�w�	�h-����h(e�.�+Ǽk�	=o�_��T�ŀ��2�p����s���J�48-�vA��0��8K/x�r��Z��T�W�[6'����d�L��T�wP'3�m���D���8�6��?���'���V'��N`��J#ı�D�3i/���b�*�qF���_C�������[-�v4�@����ox����a�0z�5|���/]4f[]�X�:W��
��z4N�"�o"mٶ�O<m����G�p9���Y_Oy���)^�+˕=@�{�����z�v ��|*h,���7���n��K;�S@捥;Sp0����&��ɸ��+�����u� x��9$Q�����4���V�H�����k,����D柴�;q�\�eӡETc�΀�#0�6w�������]�s�5��w�Y�$�%����J�3	m�rwBg�k�)w�(|��бK�j:�wׯE���u�^n8R��snB�����D�:��%���RGL�P"�#a�Gn��VV�9s����h2��R���%��c�1���Ϲ3k
X����)�ɜ3߂��#�d�E�iY�k��J_�)�u�Ҭ���e�¼�k�&�R	s'����E�;0xQx���,4�i5#{�C��v��γC�|�x��n�P�O�3?)�=O�@�C?�̬�:�;�`/}-\uV�M8�i"����rJ��@�m�N�A����� �:#k����!�{%�Ǳ��)x����%ן3��4F�v$��Z�cE'*�+LRܓ��|��U��_=�2�sRa���ВOur¢�x�_���ò���`��=2�xM�/RWՍ�\ �(ԄMg"�{2���l��>�Hn��O�����$�-����r�D��h��Lf>,h?�:���ާ���*���|�XA)�<�"�Q�yÌ'�k$*=t[5�r���ڤ�p�B6�������q{	K�Y_ｧ�q��O��fMm��Y����X#��'�G&#����d�I�f�t;����ć�W"��	�d�47���dW�2s�A�l����F�����聠M�:GԃG�O߆:�"�)
��b&��!�w>�w�A���[o�2�NJ�a�b�᤬	����AK��
������+R��������s�ͯ�G�\�!�b���ps�N�C�ٰ�vl&�."��9b�W"xWZ���������F�3dq�	��x2�Q�)�bxj#w>[��\Je��^:@A��{Z�
%�Ƈ�{hq%���M���B�l<�NJ^f���"��<��d�9�R��=u��D�_���%;x�>O�OE�˥e��ՙ����*�L�L�:�έA'?���̓҂�_h�t��5Ox�����Q
i�ʮj{������2T��ĉ�R̸][7L	�T���oX|����OӍ/�B>�ҧ�"��(���aKNz��lY�,�'�"��xr��@�儤yG��Z�d4�F\�צ�׍|PY�|"�]=�����F��x�X,=I�C����3;�:��T��7r�;9¤�W)�I�f��=xo�0�`	�?�ud�1!0�{[��@�ƹ��0E��	t ��$���Z�5=֩;)�/�-%�L�{	vC���5h_��O��c�6,_�,����;�?�b�l���nX���A�X�e�9\��z9H��]��{�����̨��͞7
���2��۬�W��t9�ʣ��m%}�;�/@���e{u��ks
Dq�ӹl�(^���H�m���d	*��tަ7����A\3�*�3�Rk^��Q��'���f։G��|�)�3�OD�X�`E��(k�����q9�ĦT?��DfH�^6gd<;�;{���e#�����%G�6ʪ��"҃z;0,5P�"��=��4��> �3vc�b��n���}�<�m�uG���K
����x�96'�>�	��|�ܜ��{!PSc(I� {��N7_�?f���J�������F�O �����,O���A���x��)����^��`��N�4�YҪ�N:F��wh��`bb�7�*(�m&����!2꫞?�0��,܍�0*E7�&>�5����e'7�&�����W��\������l�k�w��������r��}���F����}�����������,S��nl�I%hX��q�۔�v	Dֺ��g�	=��y>��
�o�6 h��	8�QKu�6c�U��i�!jcj|W��#z>͸�(�8�R��p��41T@�`����Xk$����4,�����z�t>2�x�1�����3G��Լ�6B�?;d.����L�� %����a'+3Al.���3��bt�Og���[�BƐ1M"��sy����ghJ�8��w%�}����zځx	`��'���;"�W{�}��4��4N��]���B�������!�ҍ�@sn��q�i��C��C�gzo!(���C.��LM�|^~���Ek�/�o?g-�� DKyDִ��y��A�P<�����BAs�d���}��Ul�����Ww�|m,��G&)��ؖ(F�sg~jI �oeֈ~��R=)�SIŤ{9��P�^`�(2���h~��I}�U��K;��X|�� ����V�gփS%K�+�S���;D�]=�F{<��	+_�{��y@l������A�V��5�d ^�Y:��66����(�^�b�W�,XY�ח�}��kL��k�O�;k��5�����oX���P��Ӑ�����z�'1dW��j{������<�t.�"J)��9��o{k.;B����YT���q{x�l+P��9Y���}���'攆h?�(э>٦�[	_�� ���(�Nף��ܮ_�hw����W.A���=y?k��(	]~7�.I]fq��C�7���J]�U�J�n�����m��g���ςK4���K���gƚ�<�z?����,VD��J-�F��F裂ɇ�����<0+�,��a/�	�j����f1{�l��1Z�����l�iх탞+�ۂ����A]v�NK�hVڰaky�XA�x�%$!m��p"�j�K�?3���6Г�N��:�6G΅����&�WWG�2L<����	���ޱ@|1��:8�I���W���{f���ϫ�j8wvu|��²$����%��D.����݉���
�1���(��Szdځ��r0�(��s�"Xb&D�7v�K5m����=�AFM����H���r�s�;�t1o��������%�L�p�L(�,t�A��ᣩ�@K-^�+E�d>�Q��^O�Klں��	LU�k�������{����f1���N�̖`�|4AZsRw�9�|�$
��H7ϛLᘬ���<M��.�mQw<�v��/uF�@�y�#FE�+�8�^q;:A��˥�ȏNc콢*�e0��aB�K��K�F������@_�C��/�����b�7#9�G@2�R@���%s
r�$��;����r��>Vw��Q�� I�C���-�%E,�:�/����hQ����[�`ǫ�bK0���0z���ֈI�������N֎�&q>;w�XJ?ΣLtZ\��4=H�jd�����J���N,n�LTj��E+f�*��I"��_Q-9=�q{@��]Fk�b��rO��at^­ {_�%��i/�aZ��T�͠G��dB%c��cGFA{cO�a�AN��Ǿ�r��ub�V�}��q�:��q'���q�(a3W�>y�ǌ<wlvk ����-o��4�D�{1�5G���ů�/�M'Y:7eۨ�h.lH5r�bWC�9�nώ�]	9�q�p���5��	�Y�;64�w�����5oFnlE{�`���޼�V6�-����?27,gI��u�=�5��Nv��y�
�zЈ���?��\�y]�HG�S����+�u�Y��y:k~� 6���D4"�8Mi�Dl"~�d���2�nvrl�I5���H��lQi���.m��znX�n��Oč�}���%�]<^,���0���[�_<'��t�5l\O�'A��Q�k�9:QI�im���F�P�F6�~��}�U����������8jU�����o�q�����f"���?*L���p%�^����~�P����z�����W�vֳ��i �Y�۽9��a������k������՝��4�����t���ȇ*��yR%��U,��J�Q��b�J?B��+�O~��H���w;x��~���g�a�	}�M��ߋԼ��t��+ m֑':��5ػk)����9��?I�`AT�nY������4�:�y�U����õ�~��ᡦ� 	�^ƆJKx!	:�ֳ�M����랿���I�Ӱ���=i.�]G�+���̛��|UAI��w>�JH)��MOU\R�Q4�)M���7ǹʷ�2���o��|�*�QO���n���$ySg�jP���"/��l�g���A�J��MN9�V�c��)�=efi)��8��!����J[�[��d��d�&�9��O�׸� ��Ѿ�S��0���]2Z]]���nŝ>�#n'�'�����,�S���h��(×�=k���w���Y([W2K S�$4/��\_WV�ҹ������~lLWXE��E�A��HN�C���6�����V$h�뗙�v�l�A���u?�+���?r�G��~1+�>��>�� �2{y�M_ޤ[s���)��* �.�10I�Ak��}���X?k�`�Y��Z����E��� L��Q�_��*r��;V���T�����#�v(�\�+#��7`/>��ɻ�}�d�F�?(��8�[!h���"�ɖ3��???[�yqi�5-ck�iGQ����#\Kfrݠ�m-�nB��sr}^Nr y���έ=�[�O �˷�{��n5uқOx�CC�M6@�ǍI�LT����.�Ti!�l�ƙJ"�N�aK$�!0��zLq�3�!�|�PM����LDF;뢔؉g�rC	���ʦu< 9FA:�0{N"��4@�����Ψ�$��%�##1;Z�6'�(i�t��V&�fM����v���];�ٓW$	{�j.�Av"���r�A��d�m�v�h������w.�(6��{�A|߶���6	�#I�BmQ��麏{(�az���|0��E�u�H�&��?�E�.�y(��?!�Ɗ'G��ai�Xͯ�B?v5� G���%b�=�_���I��ᐏA�������������$��0�J��1�U2��� X�
~�ܟOȟ�Ӝ(� P�!�o�c���ɣ�TBX�����Y ����2�ՍE��!f|s4Hrʋ!Ꭰy�u�&��4���5���h	}cOG�*�W�U:�k5�Xo���Yz ��Ƒ��	�	#6�+��E�q��<_q�֫�>״q��9�k�Z�[N��@ݸ��L���zBn؎��`1JbG�å����N�%ch>I�g6#�c^݆R&��p�p{Ie��C�
�9:c��*�ݹ �X�vY�0��"
,��F���#��2Ja��l�	�+�̲�ܕ˶�]wM#(�'n4��ő�No�����>�B���{�L@�A��U�o8lK�o���o��E�f���K�J���l�û�K7Ф�\][11��Pb�������Vڞ�Y�N���|�ʶ�@<��(��v��-��|����ɀ���S�.�ȱ_��9.ĕ���I,��kMb��y�F=�@Ѳr��z��dA�s�`K�Z����ʚ��M'@yܿ�����/,�1�[#w������+�v}� ŷ$�[�P��|(~ �Oa�qWɲ~�4Cq��v�A�F8��e��≆�!n,>L����6)
j"�B���_����6P�����%s�Wy��wu�1Qz�����A�[RP�W����m#��j�.��7�?�'�����*�xw�|�ĆQE��w'�U�Iٸ�=�t������{�9��S�9����t����p�yH�I�>8p��B@Tj�E!/�Pݴ�S�����p�^v���h7qs�y�OE3
������$�(�o�Ñ�o3��և�R�C��֬*�1�!Ο"lT�{r��=; /O�L�~T��\����!�
�X�	T����W~<�B:-R9̙ �˰f��\O�9ϋ�i�*sLeQ���N�
hȳn��a���7�.Eg���Im,u$<&��y���cV�tP�%�_���0f>�PXޭ�p�k��Vy��s��p]�y�z��������c�y�Xpu� hk��F��y�sҭI��� ���Y���a@>2�zZ�Ʀ����S��9���L�@.A�G�
H<41X:#�	cI��LΑB���L�e����@�/�FB)ƕ_��D���ׇ���%�1'5�$ұ"��e1�N%�Zre������4^MSr��#)�;��ml��祃b�O
@�B�xZ��ʙ�|EJ,�eԕ���Ł[�,ПR�)/�y.�t|��:ʺ}s�8���}:�J�JZ3���pklHKe�u̖b��F���U��X�A^7����_FY��}G)ġ�J��$-�_�m�Vnf.Nc�ɽk���0��z:En�AV��F��bO���i�rS���ъ̱�F�;��% �EQRF]��*@�������ƴ�.�b7��ެ�G:��	���0\�'��V5��A>d�W�Y��Wj�9";V[AP�~8���v�CtF܌/3�q��[F�I�&X�c��z����[���]��w�_$��y܁k��2pl��۰��0lc)��Ow��JߡLW}�h�Ȅ	]4|����+��Nv{Q�k��
-�J�|d	�[������\E�TN/�bʖeoF�8O�PlOؿʵT�����6��p6~I~��<���y�)����n�����w��*��M�aI7	����V�	)����^���~B�>af�&�$V"u��t\'*�B�$A}��p�܄��%Z8��7Q����Oo�sc�n���]ݽ�ȁ/�}1ۺ	ENnu��X$��v��M�*�o>�1iZ	�j�fR�2����a0n����q=Ĺfݲ;���3xW�F��� �يb�OT��.��%&<o�1�
d�a�7|f���r��!�RT�1
RA��RM���i�Z7����ʓ�{Yv�f�9/�!(G&�nE���k��E5�}5)i��SK8>h��hɈ�.��Aug)��5���'"d���Ǵ�`���t"&&�v7�%Ū��i�_��5�@�f�a��-��st�0�_ņ";�Q=��#G�ЉAF�r�:#�t����3ە>I�����>h%�P�K��(�\�ǖ����_�˿����3_�2$��V?A��51$��R�4�LE�����D� +�U��4��������;��97�z�ǯ��`�}��n\P�@M��������5�N�&$m�eΝd͚�U����td�{����<�g���ym��� ,�ݞ��|�:�9I08Ʒa�T��j�q�����W��{��Q�ZN�,a]���x�^��61����M�r�U/)_��ߒ��+��|"C>r�-�QU䓑;f�%��`@4>��>���
�M�u(O�ѫl��p;��U`34�Ӄԇ/YKP8	r��H\<�J}�$�*��>�C+k�u���B�\W��F�b�X�(�`E��{)�c����3kȥ~��9�;�[��z�v(ă��t��jJ3�.�o��|�]�,X⣲d��ht���T�,���#�σߴ(R�<�^�rNh��Y��d"҂������ *\��lO�!�>f�#"�榑I������z�y��ں����A �p�˳$8�7?1as�����)�Q|�!5���ɺ�S������3�w��a�`����sȞ�"O;T�m��xS���7�R�HFW�L�,��䟝�0�N��J�m�j�����D`���ٻۈ���:#U��J՗�'�����m���:^��Z��gZ3?��3��nyT�߾����#�J<\����<4һ�^W��!rÍ}=	��E]�cK�'�O�N[���t�g��;2Dl̔�j���Oq�+l��x��Ɇx�l��d(J{���#jI��\
�~WG�ȭ���bq��P �����B�$rdB�|�>��z{��[.�>~�^�9������$���?����G�]��%���A��)k��
���PP��~����Q��Wm�͆4��BO}�����OaD�?vko��@��MK�u��D*W���tB�Ko�������О'� Z!.��<����S��ZRu嶍 �j�{�x��_?��lc���u�)��M�K��Ś�����
:�(�W�
%�Ӧ�"�['�#G����V�0�ґB*"�]�c��<���1���S�Cђ�ܡ~���t��7>�_۟�s����l��{��'(!��ݘ�c"�H�Լ- ���=��|��� [��:�9BDa���v��}Q`��I�ɶ<�썇���P�Hp��:o7��t <r�:�[�$ŧ٩G�x���bC�j�ף�9�(��@^��c�ŒB���A^ίxM� �*4o����p�L�ٌf���(5|H�:W�4�4Ye_��Тa$�M႟Ӏ����'�W���p���NaX���Y���ᛃ�!qG)�>�]hG��p;�y �,W���5j��6�nxyN}�A�]x��2�$��%�S���[	���B������7�G9ȵ�(6�Z��a�0>�S{���-���_Vˁ4���#���B�q���t_}ޙu��ez�)��G���g���?�E<+�q������x@2�C��/���7$��U:Jz礼��ק�|�h����1�*I���(A}�����1\���F�\��ղ��	���e�{-���jL5IU�k]������H%�ҝ�˦�����}�ˬ���	�-�
�}n����z%�t�E�<����%�u���&>:��9�%���v�/-�#\e
����=k�40mzH"|�*��X���x�;H��aZ奕���D�A>�������W���.!�NA��̋���$��@���	�cx��4��|;��pm��C����%�����M��O2�~j�N��z�"�3���&Z �f@�
�ڐ����U,Z��������m�7x�/n6=��:�S~,���g����Lx��_7�*��UW���o%���X�L����<[~� ߲�@_mK ��VNf;Y�9�N�*7�I�=�k�A�b���fl0�w"y>�)�̱�I[�,L�q)�j�3pV)�^BzK�I��i~@�E�?�~���7}f��\�_o��$���7��ET&���7Ӣ>��*�ؙ'D�8y��y��_�C���������v+s���	�Z��Q��Le�GOǍ]��_m�oh�ߎR+��S�QvӁ��#��ĸ')��.�}<>̳D�<8��nJ̾�3�sW����B����{(���Rf/�� �ђtw'g�)�,����@W��M��_#�!�W�ݐs��	BM�;���}T	�$`�W�A@=$�Ft���3�u����z��8s%	:VE�����p��5�f��,'EǊ�P}T��M�Y���`{	"l�V;�Ή�d+�Ø��\+E ��79��	�_��@�H%�~h�۪��4�_��=�֢�5w_<O���2V�������J��'q��\�z���E!ˈ#m�H1$���:���;��D���(�Dm8S>��끽rKLg�H���QZ%<V!�#+�`��Y-��
�!y�8��*��k�L!�#�$�?�ÕZS_�3�lPt*��D-����ז�	0��ɂ�oG� W"P��8P�PD���˖0�*`�����1,�n��V�~�X���Mi��,�wYa小ܿ��HW�pGB(�@	�|f�V��Y�d���y���|��879u0��YS��Q����d�F�Z�:�o�qq�oS^��mfF&bPqxc�PeyỔ��&u6��BQ���U�2.�����1�_����Z2sc��"�s�/�n��l�P0�ԃ�,6��M �d���y��%���JMh�H��Hp_
ŵs�����k��O��z4Csr�鎕e->�N#ͮ{�h�fra
`���1ʅi�����|*7�Fb1ͳ�6��4_�u��WI�����ui+��w�J�L��H�WB������o{��lW���=��}��=�Pے�"5q\�{w�w��v�����w������in��D
�2||-���m�\O�9�P��6:3�;�\�1�_C��?9��6����,*�:�>�}�%���0�0��H��
�s{.�ȁY
�b,�Wp�s��ڬ�C�n�L���1 G����)בgFl��!Rc`���"Lp]��׆f�R+?}��
V
�L�~/���Wf���uѪ٭��Y���!���SrX�W<����*S��0K���7U�	LӚ�)QY'�@l��Y��<kn�[��L�m�r���[$7�>�w���7Xyt�o���Y��?t�s�[l�/�#ˑ��%hpz!���:nڏ�(+�}K���޹ݙ�a:h���
!�h��Q��t�'`�#R�g�%#�풅r\7�� Kg���-|����n'R��HL��r[ �*c�~�n�l�=��)G6���2����:�|k������S��g�/�&������U8�c^�;��g�ʐ	����1��YJ��B~���DYB$S��Ђ{j��*�B3{�u��b圏08B�F�:j794�d����+�+�U�K�]�ں� 7�Vv'���#�Q�]5qA�r@�9w�	�P�ß@�#��6���|T��dx��U=���eW�m3i���l�j��?X�l�5u��*�*�_�%�黈ĭxDvy��Ԑ;@�Jl�$�St�H��@{c�wsS�/Tw�h�|C�n����N�q�v���L�D��C?�%!f���{�A�۬�\ l�lt߷�O��-vnk��3W�:������K*��.�ˊq����7?�oi0+��'M��AJJ�X�[�?Z]��3��*�����p>?���p�N�>�=C��.�X�D�p[TUi|��rL��+]����S�����o��ԧ��z��b���斏�5��E|�����F�NU�O�n��v[8�JG1�\b�a�0lD�K~���0�p���M�����$�^����>2��9j�K�q�g�j,
��mJ֙1��^g�!8�[~�+�J�vI�$>����y��S�l������$���j܍�IG�܈5�{5���G�3E��Ze_��|E��1�Q_aF��q�(���D��io��OBO���(�XFMP������m�}�i�t�'�fT��V[�$K�@@�r[�w
�C�-i���vO�C���|b�]�d���Ta��JV@��f��3��R��/�\�Q��3��	����h��=�3�l����m� 2�5�Ē���{^������#�S���+��&���/~Q�i�i��1���!MeS�����O�>y�C��ʹ�4����p��Oޝ\�7�6��-�����Y3,��F�?�ٕ<��8w���TLx��w_ ��*N��͋q�2����"��##E2H�Yπ(lPΫ��n�(x5��kjْQJ�&��B�
|pb�����m;ψJ:��:�Y���\��k��z��
"|�Jhd�~9��'��{?�0�����Z&LZ������zI�^h�P|T�G��ו��V*� 6{�-��/�3ϝM|�����J�=�L��`|�T�?�C��x��(�����+Ra\�6dBa{�\z+��G,�,���T�U��N�ȫA�f��4��|�+�n�ݲ^R&��e�"�׭V��D����W98�֓����A�rcc�А@���f;Y�.�N1��Jx7�HG����#���\]����,b�8�l�N{=���� !]��͙��Z
��d��H ���zS�S��X�dăy!���"3�h��I���n��1su��� �|*A�uو��\0�d�M1��b��^F�Ԑ�|NA<�5��E%F����E�m�����o�ka����e��F�ڬR����w1�a�ʎA H��eq�x��v��$L�����mp��	�ֆ��	;�PU�6^�5%��h�毿�*�B;�D���./�dT�����JF�|�T�2~�%�B�Y�-�lj��L:)�h�)�9q�6��0�R���|�P~�,�z��KfXqw��F^����5��	���^#�����bU��9�d��
fv,^��(����7;������f��r֧wM����o����ي�:+���]���}�[q�֨a7!�(����[˳0K���zNc�	���5fK�e!��,����Dr��)�ɗs�u�_P�uT�<A�wJ��a��@L7fn�V@�)V���{�\��Ʒ+�� �@�� ��<f)
[JԪzo8�lP�p����+�Q��@�W���%%��(�r;v�6�V:�m�ʙt% �W��[Z�s�^�Wn��쁪�"���֑�"U��l�HgcV4��
��9��s���Ȱ{,g��x R��哂s��%��ٴ@��پ�������d6����9ݺ�w?��id�����:Y�ս�A��OYlW7�?h�f���W)��+dF�B.�DgX�K�m<@�pP��jN����CՑ\]�=G�7��,�`Fnmc��m0jF.�S4o������)�z*��R!�>�LJ0���� �QD9�m�M)"p�M��+��&��:g��bq"��e����0�8��ל�Z*�y]0ς��B^�a��1�Q��85<xQE>b$4�Yof�
�DY�v�3�ث�i]�XL�/�q=�����=�ݨ7�f�H��&�(�n��J��Z����A�3��Ǔ��+V�#�Ũ
)���J�o����#�m\������A��S/�� 2��SEt�T�l�Clh���Ђ�Ș�8W�K���JE�q٘�Y�����&���<!K*��t�-eλ����V��b|��6z�b4��p�
=�ߝk���VF #��A/7���A�Ԟ��+7�޹V5K������ �E�R~E2�m�.��G��@��|g�C��!��n� ���o��h�����N�0��Ӳ��$���@n��Q��v=d����&��;��!���&�z��K���&x�~�탾�ّ�!G6n�G�Qӂ�~
�p�p���I=��*l`�q��v������N���o�:Ԟ��Ɏ��E��W���'���,�c���3k`:������IJ%��nF�$$0�[*}$�,S6�bp��c��	(H�>�{ij����W$��z�����(�Z�����-Z
Շv!���'7�.%m[/�ud�`�=��O�is���T:s-s˂&/^l0�*�)�OO׬��B8�'��q�|���z�w��Y9���PP����R{G`	�8��g,���9~i����u_�%�{Ls�&��*���f����t�c��~��|���o�d�y���{`+�s�(��)2�Y����(�*v�s߫v����w��9-B�X�oBf�Q�v�/e�^��[�a��!���H3o�As��o��B[�?�����^y�Jf7�!Ӕ�c��뉉^�)���>��G0��\J�f1H�_�>�uG�y7���T�T�,ȹ�W��\�e��Q΢��V �A��R��-��Ӹ�E,B�=�p�92��������w4���<Ek���]C�6�aJ�_�**�i�g`���8� )m���@�n��L����T�#y�R��^���F;����{�C|L�
�}��y�^W�)�`s8Kf�����)J�}���9�&��d���Ӊ�IW���z^��b��a�M�%�n���{K�z�z�@+|k�ȉ��t�����V�t���& ��Xb
���F���'-8U��#�Npt<xw�)����=7�dE����.=!��)�g�������O^����X����� l�X%��O4Ԡ(zJUi�5Įv���oK߷��rH��Y�a�]�p[q�<�{&O�C��h�A�FZ���Q�h�]���d4����iV2�g��7a�3�B��ٴH2J���fuF��cQ��-䠡)$���0�F��gs���	°wj{���:"㷔��)cl�u ��iq�*1��>΋���E=�a'�a���h�i_�(Em<b��+|��\C�0���@��mO������]R��\����f%5�Ȣ����F�ս�&��W��'��W6��|�m�3`ŕx�Zn��ful5�fS�@b2�Z��C�&B�@�8���<��Jr,-�o0	�}��8�?�N,�I��t�滓]�ʶMs�ف���J���Iw6L�j@�='7�w� �o7t������'*FgK"W��;�w�r���g�����O(��OHV~�xh��ܤC�Z6혫$1⼕���w4<A�����]��k
+����������_���F��,#��|H"�Ԙ/�Dit�UM�F��a�taW���
/�۝F��n\S
}rP�H�M��L�Y* v�Vj�N��������`s=�|	�`\����U�7PNzZ���ܛ",JRb.r!�ֿ<G��N�շ��(l���='�9�n�-��&6��,���e}�;�:�/��xMf �!C�|���=&�EE��g4~�em�Q�X�~ySC2�@�oGLD<7��\j�G��M��n�4K�#��wl�r���)tX�쒭��ʢ4��~#�d��c��D�U�u��+��j�D��)G4Y�]w�����g6/]�OɅ0=����U �O c��z��{=���<���t"IEp��&P�]^��8ӎ�!Q"�����{��g�l�1P�zTۥ�P7uC�s��^r[� IE&;l��j1��AJ|��|����s�\<��+�(,��]���{s��h���c�,�r�" ���448�uXK�)�0\WSu�s���ֿ�1IB0��$��� ���f��_�#ާ��m�uF�N�֐7`�K�Dl��x	��7��?��[�����y��M5�� �"�>r3iq�h��Y�"���D)#o�0T'z������h�L�G��[�r,�ʸ|t[񡔊ꁣ9A�"�`�gc�B� {a��?(�ػ��~hjK��cK��"�Z�oi�(��D
/�h���F�vI��m�w����5����A�UdY�{����G���z��!�	5��1�,ͭ~Q� %�������Q�^���ml��ul={S��0r'��}+�R�1"�Z�N����=(�dx���"�E��|��X��R
��o=u�u�?��O����z�҆�,��t4z5�ʋ�.�l��2*���������D\N�g7�I$y:
u�!u�3���R\쥳�"0���"m�<E��:QD|EY�<^�9�;;�f�DY��7�+Eb�f�-�ɻ�O?GG�N�V\p�k�PZn8�c�ↁ� Od��I�{�g�0�P��
���k���Z��7�vi�VȺefG�3!1�s[���ͺ��ÔS3�q�Y�\�w6���j��
�3N�Vc��aݰ��#���	�$����n���W����=�[�X����^K���	L��\l��0[���A�����RO>��"�O�jH��	F�����)��V'y�1�I(��!V�$�fE���v)ܝsY����YoFcS��3E7��_��s����y�a6 �G�ϾX�(IÎ�Jou�_`
��-�E��WD����{j�#����)1�$��]zh-@J�'�rg��
̆�Z�{�V����O��|۝(��,�� �^�u���28�����H"hI`�E��h��i�m�o"e��_++@=�^f��Eh��b��!��|D�A��.0�ˋ�2R��김��9؛r���yV��n:mC����["�uZ`7���e�yb�
F�v��_Do����@G�}�����!��h6{�60��.��P��Es��� 4؟�>?�kbAw��ƚjU)1jw�5BC(�轺�W��4*z�4����׈��I���e�C�
��]h�f�K��,�u5M6��R��M*���P��~���r�^x�L_$���7�TF��tJ|�_h`YH���������G.ښ�(�|�
��C��P�R�V�#1CZ[M/��ߧ#��E��ңR�$���a��pl��U� �xF�؛��(q0@m�O0����-w��􉙙#�`IrGuL#�A(�%���`�G|�H�4����2��X��2�u^��cяYb9ؔ��=(��йh<�e
V�-�8�V	_������}r�	=�������b�ho��C-�.S�x�%��}-t����o0~���QJ]�j�X��۱_<8�c��Dư��9�H�`��;��;PX�?;
���_�H��_3n�����f�W��u��Ł�܄�:�~T�f�;�k��x��(��0܌���61}y����A�J�˫=iδF��&�K�.I�4��|��އ���Ɦ�F `"��f�Ip�L��תM��;�#��t�
h<գ��#|���p�E�M�F�3�#�Nϳ���/��x��� �q̀_��!�W�Ӎ�}��:�!yq���%�&��M��6`�/Xل��]�~�}�7����6��	��P�!����t�������`���d�̡l��|�V���}�,����'=��Z�+N�����k���2�.nO���
�}��U�lu/\=b��P�d)�RK�;�f������a>I��3v��A+��r��~��%��m8�	��4�ՙMIB� ��9z�š\�)A�d�A8����y	jR�Ka]���)��p%��AY��s�ˠAM����]ǜ-��W�[���+�/%Yz"��Ӊ��3��"#����l���$���*p�� w�1Y�����6���`eB �#(zI�!�q)�g$z8\v���	��hb5���e��~ӻq�8��B�3�yM�H����J1�:�\�18+��r)�]�l��L�n:��+7C�Z~X�� �{�P�m���A��u)g򗕸�6���-N͉��b-�*�L�?��ѩI���h�E'P�;��z�q=n>�+�2�%��&���<�r*�Q���Sm�i�G"�#�c��X	�z�I�5q�f��|$a�^Xͮ)�P�����/HR���>���i)�#�I#�C��>ov�%|!*��l������tg�����qn�3r:��J5𰝪��(�W�)�D9�\���%�^Q羛�$��8�i���4��Ph�� ��]�J&`YX���&�B!;'DL0~�>r�uB;�aM��{�H��'���L��h�ÝQ���0�B�i����O�Dmd��r?�	�A��]�z�Z�{�mJ}����>D�z{�����f�h;��#K,��L>��B�l1;+�2,{3{�J��#��=[���_K���c6�s%1;�X��A+ҳ����f_���{��8�6�-�'�����T�"��&���#=�hF)��Hn?�����2�2���r5_�1{��k��5�_C�~9���eH-(?� D�L��-vN gx�L��ǂrH�nN���+��k�ɹh����;G+*U��HBMŘ�@��L0aƕ*�5W�bۄd�����(���IX}L+�Q�6�5��1lՓ�z}�܆!�7b����8yg�Xa��/v�]����pPlM���-�.�H>��
f5`Y���@�2vA�)���$�k�Ig���
�񊂸aX�Ǫim;@����'��<���~Y-FL��Z��F���"B�v���t�ؤd�q�Gqu��� ����t�(�k]1�/-�ן'�@�-��-��%w$7�`1�wo�l^{5F+C�e'?�ϯ0���_��A_A鐄�Te�y+�{])��b9>�V�AU@������ .SƑ򉾰�+̩M���>Lqv8���Uzl,�H�,�הr��JW���W��a#��s����2�T�����
KDCH�F�%q���T�3�̟7�<��tɚ,�}c����C�ǡ'(��`�ފ��,68u�����#�)�	</�pJ����;��8j��sѡ��a\�@ZJ���y���U�B(ېV t��̚[,�E5z�׃0��=@^���"l L^��e.�巸TG�(�v����(u��d��f�O��+�RZ�r�;J��R!HjĊt89~���J~���8ת�f0��-���'���4Ģ�����`~b4%�� ���C��	@i-@Y1?���[s.gMBIH�`�r>' _<��(g���N˵�`Tז6[x�,:!Р�+���Ṳ�g���5YGh8�0�{av�	E[S���y�x7>��7���D�;���%_��C�E����{
��SiߵV�%��nּ��3�m�����]���{4;��hDږ�����N��vԚ�Ӝܮ-�Y[�wjM|!?��_�W�z�:�^8?"��tD�Wc�� g�(�f7Tm,�Gi(��Z�&mnc[��і]�
�ي��i+��pNڏ��Ꮯ{�����o��ti}D5^Vb����~�.���jq���P�]���4����<�`=b4�-����-2�VI�'j�6�tG�f�(����U��`=�}��Vl��[���v9���j����V$A��4l�Px�4#����Z�u1M��E�"���.SկA���R�97�v� y'(γ�я�\u��y�五����D����o[��%ܪ*���i�$h5,Yd�Ϙ��j�%m�]�Z����G�{��oB)���ce�ͯL-��j]R�L�~��[��\;�P�6�p��l�� s"��/�(�\\���t�w�0���Tx;x��c`�o�m�OMÛe���G?���2��ss�2Z��� U{'���������� 9�T�Uw��$7��&�a����TS6��o�8}���o�R���O����8G�rG[�O,�����v0�r3F����������p���M�֨�Q�\���N-��7\<�Nq�Q�8R�e��I��Ҳ��悉������B7H?���6 .8+�b�R�W���c��1O��1s��ƍ�����|� �B�h�6F���~K�z7~Oj}��Z� AI�#���uV��P�a�;����c��iMw��ZЋ`̎�x
b����d�(�#l>UbKzz|y���C+�P(/uc	��ɸ�5
��^�����8L�7���0���COud�Ճ������Э�iA��8д0Q#/����q�'�_1:
��)!���E?߼�~���Dr+
��T#f���$������̽�cVĴ9 ����R�AUi��%����<���H𯗾�Cv&���\yu/��2�b�š;��K�;�a�D��*��\��܋���`��T&r�
��q��`�9V̌m�:����P����z���#v�i�*��t!*c��z����B���d�l�ܷ#�Ի3l��x>�~����.Ht��dx��,7�5�2�:6�,+�C�\E��Z 9|�]  0�7c���I;	�?t3����Cw�?���3���7��e!�Dӭ�y|>Ba���;�6k:6$d��&��=�hX���E��^���2/T ��u.�E�\&��gō�K�-��ؗ��� bW���G8g�IB�M���G`�4@zR���ḑ7���$u�F���-�j߭�$���;�ׄI��?�	�Jc��ǫ�ZU�TC<,�;kO}�R���D��!;�5^dduc����-���W��������cI�a�A��=��V��W��F�|��Km�����f��p%�=h>�_��o�ĎQ�|
8"׌yj�H9��T<d�|U<��8�e�72��z9z�'}�b�od�)����1�C���=B�W��Iҗd�� ��vU�3���
�B��@���~Dkp�(��g��4�#��&�N��.��nẇ�`�/=7�!㑹�E�~�q���{�6K��v�*�C,v�[�����r�^�\�g��H�E }���s�U��Q�#�1���@���κ�iy'���t�"E;H�?�T�.4��lr��^���'$#$ŉ����ꆫ��E�lV�.�淑 0��&�oO��|��L�ֵo��SI]4��eo��7_�TZ4�'(��n>�.q�P��g칆�v�M
Y���;D�]ci�A���VM��{�4@�`U�!�GP��p�r�H���o�t�D��ꂷ_wf��Y4? �1�cl�e��zx�����B��U���b#̍���|����}^�x�b��y�7��|e���Y���߷3��&�RK���Z��W�`Ӹ3Jִ��R�%�@$�.�gX���]4���=$݂h�_J���/����s��͕��&��9��r�-/�kk����Y��5���ʑ�9��5ϰ,IY�A�F��0�w�jUj�`�F���o�k=E�/Yݏ9(���]���'9����i�5"��4@�4�S��2�>���:�o��Hv8:�
:Vw78&��Tf:ʗ�Y �%B�_�6�q���Ȟ9��⧔��b(�����^��e'��C��D1�7:4���]_���n�Z��
����(��5�<uvh��T�(��)�'*���ڧƋrx�"f̴����r#�į�,��
�yOG�r�H��#�`���?��������TW�M��H߹Z���4�
Rk���-Ĝ�u�£
 �Y?�i�RLb�+[�t�2�O�4����N�H����z�{AM"Q����R��9�TB)�_Y�ɓ�f A��M��T��+f���<�3Wn3�JE�e�x\�����b�of��5�U�*^�;�����E�0�<��z�s�9��H5Ae�z�N�Zk�,~p��xs��P���!�������
ÑX3O�$����u��ȇn�zɷ���m�,���tH2����ҿA(�/��a��Sv�'�Sq�����.c�Edȸ�,9c!��v�IFU�O"ٰ�Կ`��*�A? �틀$P�x'S4��\��\�	2�ά�e�F���<љ;��ŅJ9�~7������w��@�尉Ў���7����8�׾�l����=�g�C2��8|��</%yJc����c+���ZL�4���f���'-��+��%o$G@=����V�x?R�0d����zˆ!!&:�Dd�u�hv���%�T`3�=Jq�r�xH���ӱ8�F&I�exw�������wpܡ4������SA$����̿����|�
��5:$��]�:;Y�>5?�Kd���H%]���b&ldޓ|Z8����N��į��33�U6�莼=eF3x7TbG��s~�/|�A�� ���,y>w��f�$�K����Ԁ�Þf�cF��D��C���0D�?�Rt�<9�@ ��;��\ڒ����z�6�J�&b�7^��Vc�H}-$q��e���ќ�h�̟k$�<g-����rPh�E�`����|,�/+�*�oBQs�r�m����	���+y���KC��)�3�hy�Ď�P�ē����i(�{�Ѿ6Ik����}s���=Wژ�@_��Χ��%�,��K�D���~�������nK0`y�V+����mw�@Oul�˲J��Y�u��S8j/�c�e���~�N�a�_)��Oi(���	!d0�cY�����Scض1��;��wn� � U=������2�X]\ �qHLi�K-��s�#�2$P<�g��*U;���P'��U���j(%���gs��k�(��]��������o�ڑtL;J(��eU�[��A=f�>�Q=�15�J�)��wq��_S_��ܿ�-/څD����;a�1K]�%�2aR�T��M��.Qy�yzz�:�z����5˓��=׆G����v�)2:*�vY��ur�ɤ����y^��LTt�����O ��PZnC���z�3��D�T����:)B}�v����Y'�$�����>a�g��p57Zޘ��U>`��h��%�I�̑[�Ԍ10I�x���A�&�Kk��j�V�ѿY��f� �|�6oa��{��ڔ��8c"8T��ٳ/*l�C�p������R� �d����:�Ń.lt� ��`�{�@�Z[S��)^gU���Գ)*��?6aei���?Pp�Ao
v��������x�#(:�Ϥ�����ſ ���~Z7����,�5r�K{WXCW�d�.��Nu��=��i�|i�*��65�g���F����"�_42 B3 ��*�lۊ��0�/C����S�hޙü;�7�6�{5�N�&���̑XX���4�^8� ���P�L��l�{�<�ک�\_���_-���X3%J7�5h�wl�S���yc�M�9�X}��:�z�[����f� % Y_�ڋ��CU�����6�+ uҨr��ІsT��k�Z��"����>¡��i#}�)�iUI��#o#+/�H��^,�a���f��:��J�`�"*K�Ж�����Q����B�l�b 8���2�s�2���a	<�r� W����%O5�E^):���QYɪ0k���P!s���N ��v93��W^Q/3$ ��u�>�%�gY\:im)ҷ��^Ti������������/ ���U��Ư6NPY�B��hB7f���o`���U�&1�ˎ�-�P��V����0WGN�T�h�g�u?D��fL.,z�/LE�&L�G��Xat���(�-�Q���J�����ƥ����L�kK[���;V��ز����}�Sm�4f�9�'��=Es����/F[��ªbc��5�<b#��yn�;(%�#�hZ_��:ͬI�bƅgp`L:�t�D�K��*�	c�][�ڥγ�`������ER�b��9����^�{MǪp��4�����A�[�H�!(ϳF�#�|5s$.c��g.��i�l��	Ni�ߊ=�Е�{c�Ѷ9��r�J�U��Xx�H1�=��"��J����dK���(��p�Q6Cj�L�X&���DV��p7��7�Gå�h 5�g�I򵵦&��ɫn�W,QG�t�#t�fY���A/|��F�VS�Fv r�Pm�
�vDB? "�4��\���f`\�m\H���0�9��
	����������9Wp��W��BB�f�x���v�CO���fp~9&G�.�G��'��?	"Lϴ�gL3΂�I��l��eY��v=j�w	��;YT����f0�0��b&脁���}�@�U�ْ����&	�3�a�i�w|3���ӹ�������m�ێ����(��rj*���	��GgҒ~�����5C�� xu$\���:}^����D��7���.��[U!�w���hy FOUj�b{[�4�%��G�F�+����$׊��Y}�.��֧RR]R.���cy���5�ax��0�Ѵ,f�������쐌#gwzr��ښ�-ф 7�xs�M�W_�p�@��P����z��ΌWR%�,�2΂ i,�J�ІE�������1Т����
](��vh���A�!8d�p�� �(�Z�����
{^�5-�N4iiA���gٯ������h\�jp:�`ճv�X.ȴ�܄�����C��D>�׊�H�'E���*�nq�g�����b;LXlb�e�a�8m����k��8t���O�!i��04�)�1�-��r7�F���[#��>��v�iZ�/Biop�z������^4-#����w��������z?��3�B �߈�l2#�U6y�a��T��5��x��8��[!Χf �D�7)=���2LJ�6��K~�J�{l��1TYcd���`}� �%{R)χdN�`���_]���m����h׏��Ly�l���,����%�K�ã;p/?*�L��j2W�n���fE�v�q�e���љ�\m@�+�q��Ĵe�:L_h`!����5v���+��yH�R~�~�F��~jir��}G���c�7y�}�����z ]"�D}<xB�}&3`Exv8`�P�����S�<{���|�0w�x�;�	)AS�%� �]�"�z �m2�]�b0�Q�~�ZFn�U&MF�	����CSt|'~�cJ����geVm�`���h��)XS�n��˿��g�r6����;7Uw������|@��_$��o�3���'"|�.��x<e	�(��*>iz��� ��ǵB��qNT�@���i��I���x�Ĉ�B=j��]$�������0���>��B����r�#�b�[_��GS��N�$���)��Ӭ�&;�4�,����v��Hk����;�<�E^�-X�'J�Hox�*U���o���S�ɾ� ���=�G��־��<�z���Ey3������(J�o�yZ�lWm.��7~��O�7��%{�#͚NH`A��높�6��u��z��viu��ٯ� �i�Ky� J�r�~�;�����o4=�=��/+���<��x��=b��g�ð�7ן�?�>i8�6Hh��Z��&���3/��G���j��'h��[��Ok�iS����ԶFEc|⠻m�blR�m��X��� 5M)�}Uo��ЇQ�oɔ�_�e@
c�t���.�(��~_)��("�z�����ښ98����|k�!.Cf8���/���!���X2J��ꗌls��s�B��n�Pg�/^��q�WTueO��aE���8>�(�3��ݙPV�Ir'�v&���H��3�;f3�p��z�R���fv��W&���xa#f�a�`�r�T�`u�P��S++�L�I�$�B���(0��w�Sf*��,e�v.�/9�DG�^��Q����������	��i�c�2�s<н!E��|��g-��䃟��DS#�?��}*L��2Ģ}��h��ť�+ȍ9P�����}�a��r?��z_I	���lT��0��U��~=r�<R�K�`W�y7�>�9� �O|Uh�@-������Å�pn��W���0_�<��Ñ9�Rwv|�A�� ��q,8K�b��� �BF�a�x���u�&��M�i�ʉEL�zoϱ����������_9��1�6�r}�WdM��6x ���$Z`"�h�FS��Ͻ�^�����ֈ5h��Ͻ��̻U�V�N�t�0�Uع=!����D�#�� ��}���/Ĝ��tEI >����f�wl�Ĳm��W}�S�#7a]�C�`0]��s�;ߨ�V�w�%;��u?���mP�
�5�p�7�F,\�\�R�a�g�y���9�j~)��MҔ�W�8
�ܦR�ND���TP�i�ى�(!S��F��7��#��i�Z�E�}C�_����	��2,�O$�($  �D-񅛂y$�N��p8q$ye��Z׵ӳ�M�Ɗ�����PN��WT�(�!�70E
��Rv`�$H��(�o��dj�|��[`^���F@?f�tS�vҽ!��6ѐD�S�Y{�1�媺OC�.�N�XI��#Su��2(�蹂���)�z�me!��2�F�{�"@Oj�96&����E}�û��BH-�&��<���z������u�Z����CQ��k������نl��#��]���_r;�ߘ茗P2v�$'Z���Z�����,��>>�&�������p���Nt�F̚X`��*	!Z��S��Z��b����_/jn�V�\3�����+~~�r�TD�a��'9�Mw��6��RC����A��,E�dO��oHV���|p��[�w��R��[G�� eaf��tm�c�E����z3�Ǚ��@zb��b��D��Mq�~��8��wl��p��Ly��\J���­�7������Á�J7�����¤h��{qF����w�J?�ɳ��(�-������ �m �q���k��nQO�&��z]�Ӗ��m��6��{���u�-��Ap7F��8����A�Ȓ7XcE�,_��3��N`�"�l�C,鰌��˞��b!MױD��נ�Ѣ��n�K\:R�G�l������Ȕ������_�Y���\˦y�S8m%�� O�Y]�Nұ���:!81���q����D����I!j&��r>-��	#��#:Om��<�}�xY&/Ds�H�9��$� 2����e��IcP���P$��p�.�����#|ږ���2{
�Ncї+)�]<:�NE����5�W�0_��g����{�2�.Z��Wҋ�F���ipl�R��A\��{S]���~#�m���p�{�@��l�Ԥ-WG�$����������ehjnW뫯I�v۹����D>[T�ա�?;=�bg��6[޺wM�T�[`��Rq>;����S�.�a�M~��4��M�*�~
@aN�:pD@�e������M�X�==Sqk��`�儙�ub���os܍�����C3�#
��ԘV����� �P4|���R=/�Tg#D�� �	Q���J7p��
�m<�=򨈉�o^���	�>���ԉY�@�%l��Ջ/�6��;"FM�]�ՠ��0~�_ۋ�3�qE寛����bB��b�M�z��ӹER�q��T5G��|�t����$nB�V� 0�x�I�	�n�$�݀�R�2���e�������`^(M=1S����������oVV/�D\���ײ.��	ߩc�ao�@��E�}�Y������9�U�}b0e��S�hJ<�U��!"��SA9E#&�L�5��N�א�y�L���8�"*OͲ�&��\U�ȫ�4K.ua�>��%����m�-b:� ڑY�����䲲���+3~�wOԯ��ٛ˴��@�]���g���9uG>�y!dC#�{0�M>�[�^.aK;L9����5[4Ӟk�'�:G���A����У�m'�h�S�N~S�K 5xG�M���?6n�	�b4HY�W�rֳw�o��JK�K�5h	p�x��-�j���yr9%����H
�IJk��:��,��牖'�J
S*r�ˎ��K)�#YQPY�?FHdρ|�5�u�Jlv�c�l�*v.�SXǭ�9ihzJ��Υ���ې�D�p����	=�?>�M�$��O���s#�;���	)�g{��ۨ��2-�s~i*3o>o��Q�Jiw/<��q��\�ɯ�>�w�-�vk������3�S~���6�Ք�i�9�x�����n?X�e��r�N?Zق+�nB��Y�-����E��Y'�Ѻ�P���5B�fߏ=2Õ1P�x٥�z]�1�@@h�X���L&���_��U�X�������V/�4zi��,L��I��ĭ$��^��e����虭z�$�5:����	c�Td�f|w�h��X51��%��
����#!�NԊ�D2�(67e��{
ط��R��� L���
1fs1��c�9s]�Z
��
w֐t餮F�ՅE�x°������
G�=(�!����ճ��g���`/��w����+4���w2%�	 �u���oQ�X�]n5Ʀ���$o�p	Y�}�`�k�>)52�C�ꦽ�bw?*�7��%L5Ey�rq�����i��/�6WDM�E�f�����}�b�#C)o2���
�	,�p /���&���R4�k�<��,��BO��?�uYUy��3���/���g��1a���Õ8}.�2N�T�g�L&�w�͓wm
.�Ϸ*PW1��h
�
�@�h����ݩ
e��L�L}�(�}�Z�b;gr�8���l��@g��F�ou�׍��8|����H�^{�o1�B�u���U?Z&��@R�^ȑD��Ng�8�%���";/�k���ڦG�D�w�Z?'{�A��!ܕN��6��a_T!��Xq��z~��v���.s�߷NT�H�z��D�|y1ID�Kgd��?8P���&�S��9!�dR)	|�Fơ��_���07�1'AXj�a�
�����7�Z���42M��'�I��P�}���q?������8_D�(�b�`P2]����}�j�64��mS�0NFb��{�M���� ��K��ԟB���떴~�:*J�S��8�2al�,���0��aF7=�ql�P�.���$\��`�� X�4�H��A�ǅB��|�)U���=�I>�l+���C��x��[�L4�/�Oƹ��^Z�(�7�J3o1��h���V>c��F��:}�\�qm���~�vY7�U�rӅo|�7bX�͋��,$O��x�p&#NoDJ�f���Q��|�R�ֽ��$��5�A3���>>0;�j�1=��c�U�L�9����Lu��nt
[W�?�du�9䩫6óP,�,�ZNi�%|~ �/0AO{4�p���rdz�?R�L<@���1~/�6xZ���@L��hp���G�����k��z����D�܌s�q'��я��%JPZ��fg����|���c��V� ��E�ּR^W<�hI��H�2F�|��"�둕�����0�`*3)A�`��o-JQ9�[�h%�hb���z������ڕ}k��r^�d��|.���t���7��o�`Y/��󤷘������mZc�tא� u��-ӊz?
=B*�1���x���Y�7�}H?
�����W] ��`0I��%:�n�q���swI<�^�&��"H#ڸUJ��1� a*��[�WJ̿��J
�ب�o�?�,�HW=��w�'D�������O[^���W�ٴ;
��PR־�*C�43Ezb�0�*����u� ��"��M�x!o=�W�8� ���L��<״W3��k��v>b�+a�$�L���.G���[�_L�b��^Oh��������
"q47��1y\c<N�OV2��J�]���������L�a_�����T�L���vN�F
S��3�J��@=�X��qݨw��S��k{ȱ�o�ȮO�������yv�#~������f��]~�?o�շ�xu�h{��T�`oO�WVuO��ꓛ'�sl"'��y[���7��p�����rm�^X���*��/���_�f��7+k��5Ta|��9�5k�!��O���T�������߷��yƮ���KB2,��6Ă/�P�W.a�٤|'���M;vys%��+�s`��M`��Qje��S�H�9�+)[W�����N]��9�9�{e)�k7�>�Yw�f�W�?��s!M�e��e�<�E�jV*R��1&|e��Э�Õ�M˩�؂�f���\X(_5�ֺ���������ZO������*i?B!���J7�fK�a.k@��$�F�u�τP|�Cm���F$�<]�IH����`%�f��T�l�\�WT��Sa��]e���1�]�)���$�ksOf��|r$����×��ű�@�{�����#�D�I�܉r	��e�ϴ$I�y��3���UT\_�A�Y_�Nnrsw�����/�qsAғr�)p�,9[��3�V�����3�;�#�dե �W���Q�(�-F�$a6�=�	C)"b���+��Mx>�X�˝�R�o���8��)�!���΢�Y��`k<	�l U�ǐmin�F*Ό��/rRJ[�TP��gy���x>p�:���<Zˣ�T�w��LQ��3��+�`�{=�Q��������[M-�F�j�H��+��(X�l[G�0��.O4�������?�a_�9�of*�0��	��p�3RЮ��(���)߾y��(��;0����������\�o�����8���-�Z3{?�'N����uO��Nv���:+P�������w��'MaȐ�z�Y�P�
�-I��5��;U�>�`j�=9����=����M�
 9s:�3L �����/�h�cZKU2���C���uF!ڃ���_��L1�>�q.�o�e/�w�L���]�l��!���Ɤ���g�
��%�p�mg�eb���"!j�h
a"�]��R~���"|𾁍��gQ�(��@���u�(l"�/��h��<��,�������V�n�Zd��i,��K6ό���n�o���(3@��6u�(A���Ѝ��m���@����֪E�&=9=K�J�]vK�O��^j��X���N�ʸ�_��p����[ʲ��57�SXQTz�ow������2��kX)w	��O�Y7��o(�����YﴽT�25��h��
z�N��d9}|�
�WD��Y�u𹼮��,�T��z<;��ğTw��%���eln��*�JW;xQ��v���sG��X�R#ĮZ�3�e��������- w{��kt�O���`�xK�Jp�[��m{p�Wp�?���t�eT�9�A�dL��÷p���q���:��C�7����T�d�|r�t���o���0��^z�)Q�M��_S�9�C�^n�J\$��q��]��M�W�'�����d�� ְz?�i�����W����KpJ��;�\ }>c�+"2�H<S�g�h�Kl�7�T�y������"��ѷ���~J�)��iuʙ�~TE���\'9�Q�ճ6g�k��O�5Sh��o��a�Ɠ�#W13�!a{ϐ �M7������ĝį�ٽjC(JB�;�z��S��������ꍛ��m��'�
j��S�.^1:�`5�e+���2�{MOl�?���]��a��9^��G��9^�m���Z�fw�y�1�K���]���D �e��X��2��%� fJv|l3Q����.ii�z2#q�MQ�KWr���;m��R�
7�ۏ�-k9Q���9\g�l��5��x}�[QÖ%Y�Lc6ƣ��r���Uq����e���k�*$R7E/s�t> .�`����k���յ�s�!��N��}}�����(���5�#�Ya+6��'n�H. V1�^����D�񻻧(�+�斝�C�-��U߿)�Z$꒣S�ʟ=2���c�����W��u"������ɭ���9���W̧l�C��JGU���s���N\�D���#6�o�x~=��Z[ �cdaG���_J��~��%	n,���f��~VD�F���Pͧ�GZN�H���F���3!QV�p�E�E'���t��7��"w���ʍ[�h]k��+C����D���O���<!a�{���=�E��`��+�!J��T�5��,\c7�~l'��I�ߐ_{}�,^!������ZF��8����냀�ג%�X��N�N�+.�
UZ�i�P�`�����|�A��u�?@y;�@���
����� Q�@�V�ڛ��g�k����p�@�D�ju�q+.�l���?3F����$�|I��O����(K����5N�̥@�.��!I���u�����8q*v���Ζ@�=��	/Yj�� �� A�!�tB���З�7Ǎ��B��D�U*�h/�ݝ����������юG��G�;�l�M ϶~1~���g8~��8-�(B$���Yߒ�	Ϝ���n]�p3�z_�_>�9f�W5�L����]Q�I(l�>_e	~Բ��� &���D�X�#��ߚ������G�����T�-��p%?+.|��éU'hj�8,���Yd�9�Z9�YD�������~��;�Z���(z��TùB��["��t��1���%�Q���^]w��^?eV}}�1|=*�?N�Cm��h�-�Z;����`}&tzK�o��:��ox�����{�G+������o��7_��9YW2q��aV��pS��ߏ L8,Z��z�b���Ȉ;�o>Ƒ��Q�}��>b&��� �����L\_�,�8m��y3��BSw��{�@����,%��`r�` ������_U{ѷԈr^�SU�MȮB���|����HCu��ܣ7�����*fs�R{E��5�4�7�G�z���mf���oCt��P��8" iG+���][F5x�Lk���,	z4w��6��gUO*ge�,	e�3?\\�{܃v����23���
�(�S���RW�1~�]�+�PS�����:�?\����_J �H��c�Z8�-��anpp9�;�2�:��

�d�����,Wx1sѰ�&�8j tbo�<��jv��t&'N�_uI�1�0S3A0�3��]���qj
�)g�So9�*?U�x�&aX�C�ʊ��u���z��"tC��JVw/��[���I/�o���Z�犭������Y0��dOXr�v߈a��������Iq�Xvq��W����0���������L<1E��I�(�I9_�d#B��#(d2&��������$J��C�˸ѓ�\?jP�!��>�`q�\��J����GO��jd��"�'(1i�ڶ���{�:�iW
�-�_i(����H�
_Ͱ��$)��D�EzbG��t�Q`"�+\�(��X�݅��!+~��#���b22>�$N*C�T�� �i��\�N {�	H��Om,��V_.�9�zq�e+�����i��Y���	4]W�i��ˆt��cKck21$x�j���m��o�����ƴc��6��;=�W����۬,"}� :ܰ�VY�����d�|MZl�����+����F� ҩ��)�ii׉��)�|L^�Y�W��7%�jHP�c�@�؁[W>ʅ�@����i9v*<S�� 	�H*Z�����0�y�g� ���D�*˻l8 R�u���P�a=���k��_@vrk��ֻc<-�'�&:	
{	��|׻k�N������x�		�������xK�0�3�YD-�q�AW%�Lp!���
j���Aa�3�W��ň]�ш��S��[Foh�uV�a��C�L5 ���S�?��W���j�P��)�coz�á��Ԏ�J�ݍ�+�����yow5�F"�E [<����r�����*�y|%�U6g�	���c�Q��,��к䠹IJ%ze�e���kː�Q�h����m�l���I�.W�Tgb� �U4b�e�ZQ��k����{2�q�_�`�P��^J��ߝh��p/'[���<��vn��"~�}��N�f\�J�ɵE�ٰ���k��'��q�����ɱ/a�揞�#�����)�t}��0j��B�-{����Y�b�xꮑ5��)m��~���u$���
�����&�>M&��g
����b�����64��곀����/A�������S����=Po��^�K<j�h{=���nm���:!�5�tfF�5�n�7uc"[��[�q4�{�s���ˬ��+������$S�����y-��gs�AϬ_��Ԣ�dNQ˶DR)N�Б�?Y���9��4���GS��jFnrD౻�)��l��'h�>�Ȳ
��o>��_Q��y��IO0v�����x�b8�'{g�5]ʡP��!�n&�g��R�4�(V��-j�w�7t���(_F�z�����"4p�ڻ����JFi�CYn�
�&}Q��7q�k++��ye��!S��
� ���&3��!5jbg�l,�M�t�L�J��k����+��'ܹCB�&ʺ��&n\�*�L���!q�� ���Z�\��������;+��Ƕr.i����8-��������� �{u�/"`���"	�߱4L |i��kM��oZ)���7�齙�p��e�*�Zޮr|�(Z��a��ڛ��@���wRآkv���P��{���5T�6��b,�c�m��A9���>��n���3�v�ġd�~�����5�x��=�O5���ȴ�����]V[�n��������P�|	�<��&r�;�.䫎�D��-���]�"��`��T"�x�G�f������ם�A����ҍZeX�s����oP1�E��Bl�
z)μ`ao|Y^w~p]\����I�)'��rv6�N=2�a�b���֕�pҾ��;^���9�O�Q�*dg�V��(@�!!�GI�_{`pЗ���X�cV������(h�֙�3��]4����o4�H&h�w��H�0�Q �� �
GN0����_�q3�s���]����aH%,��"d<�,us�|S����C␞��$�>!����Bs%�֩����LЂ�P�6����c"�YyQ�@���>�>��%1ڍ5���<�\{MK��K�"��a��ιP8��<��ᱏn�\��qJ���eb��QKS��&.�r1b]��UE�wBdU<�?bvTa_Z���W��&�htD;��:���sW��+����(�k�u��8Sܐ*�0S��w�woxF��ݨ(|�1@؊�ײ����̃������ٻ�e�����;�%��Q�	2<�Pc�{���Ѫ���o�c3a���H��*^�
44�Q
�?
��o-bz뒕��[�+
v�е�zݟ=�|����ڈ�L/pg.�S�-�V��!�*�3k���Eŵ�f���{��1�:���(V�2�x��ɞv�)-��~�M�Ѷ������l_ �(w ����[�rM�/ߖC2 ����n�0J�F7}�B�!�(�̗��Ø��>l\D!�n�W��5eG��l���Pd����Dq������yu��-�̦>f��l���α/����q�MT�Y��w����<yZ��o����V��#�lS��c�v�p�]��r�{fA`��qn��4v�P�
�k�S�8�5����FR��ݱ�&q�2닎����.�$L ��9�Հ�Օ����E�D��7h	���o�qD��n%Q]�\ҿ،$C�W嵛?�,�m�r�����[s˼8Ha;�F� RcG�}_��A%bj���ƈ�yῈ�n Z���ߺ^�D�י3Y�!\�.<�����P"3zQ��E캄�Jw��'�K��+��J��';@W,��>w�9;��#Y�%�B3ZiJ�s�(�T���x�Js�uNl��MC����L�D�r��D�~�4�`B��.A#2�
<e]M�7w�	���^2��Y���<G�U��$�l˾T$x/9'��x��p{}<�=w��_�d�+�Mt��!����@�d���'�����0^�T'�����L	�ګ�t�K���X�Qܥ3��qe���_�@��0uV+���p�s�lf���P�;�'X
�A�oM�7����A�����p�^&��0��ؿ��8R�问|_)�p�P/��Dg��'{B9Ǭ^�iI��#���Ԁk��Є���4x8�%iQ�-��P��/�?�A6�H�������H���}��I���{u3��$��ͫ@L�oF�Vh�Ii3��U��q�=�z�Fg�p�m��68���k`)�E����9�%�`�Qp��g�uvŸ���0���]�Y�[�Z/؉i�W�e��ٳݛ��M�����k�IE�|
�@z�5�f�m�o���~���l;z�R�}z�U��r_`:G�����iLxs�tm�Ԁ���O&nj��"p\�l1U2}�Km8��8�9oz�!jr�i���2�������o���٬�_�y|�k�����j��m����G~�,q�j��y����|Z��-�������Ď�#��4,��=�[dI�!u\��P��c�J�o���y�3A�n~	&�ԉT��A�}�k��w����Y�����!e3�!�M���&�f�TI������	�A�.�(k��+�@,
���P/&�$��^�V!�<�iV[V����b������\�����IDUW~�_�:�LsXb�i1K�?���xği����@��}[�A�ؙ��s��Ƈ	aaܰ�J���'MU�lu�G���t��XշhR֒7���
=2�5d������EV��É	гQ?������dJ-(#��*'�Ӻe��8%W��'v�۹��A�ZF��q�\+pq3���JeL��U���p�Gڽ(o^T,Kdަ��ʳ�^7�t<����'p��^�G,K*��\"��������{�a��+* �}��H�Bo`G�߮ןI^�N�f޼���v�K�Z�E�/hhX��ߓ�归�f�N��i4e=_���]g��a�U�>N6�'7G��YI0x]��Xi�c���r���-� C���^�ͬ�|��
f�q���9N���48��|��OWwn��h�=�X�R�)ٺŔ�G���|��,��>����}r��F!{8]A*9ͭnp��8�[�3��j�]�;!u�Ɯ<�֋\ԖL&�U� eh���`�!��z���J����N��^V��&lu����4%��<4�@��6�4K��nF*C{��;����{-d3�ǥ�l���l1��W'����K(��{����j� :�Ů)�E�Q��O|M�+J�[�O=�jգB�5��I�82��S�KD&\�p��|���~�[���`P6�;ֲ4�!�+�1M%��J*\F���LU�>WR�@W������P�/�8�q�S�xuL�=���	�1�%�:�ZE�:P$�\����m��T�����D5������48w�*�R�}��1g���G���΍�\�6�r䊩�,��Cf��N��&?Y�Q%�K:s,�*/�j��G5����ײ'���i$�x$M'�eD&�
d
YO�Ů�R�w�:{c՗;7�}v�e�eՇWp�9w�Г*������{ļ�Y����Fq�>-9>���&�M}��<��
g��ӡ�0W�R2gEi�1�m����T��zoK��.BJ�՗ǭM����	-��H@�ª���ϙ�d���i���w���jk�����{�>�*�2%N�F@IuU��`߲��Ɩ�%��n���'��d�_���߶�9��z����Y�gH����>�l�:A	�}⋤1kB��1i:\��z�k7(����H�z�����#�&���>�ٲ��lv����V�����H�Jy���	{� �����M׉s���j�	7'�"��{��<��j����y�t�:c�i�O�P��+�>ޮH��M�h~?-��NwIK�,`�'�Ye"ڱ�)��)}�0S��[�|���R�Z�U�N�T��ׄ�h�8�z���I�}��.��Z�Lg	�6=_1���$Y�D�Ɨ !������P�dY�yIR=܊����e��F�aj�����F��i\�B6P�B��A�f�US�����=��w)>�ِ{r�@O�,%E1�B��(d�����͍�����(�+��m\(��;�0���k�X�㬯ɓ�l9�'{|?6��W�����]�0	߮���F�ܷE���Ă�!�\�
�`Oz����?����\)��X�%M�0E���(�
��F�p@��,ODg��K~�G��\�Κ�[{���N��8�{m����*���a2���!e�x��]���ݤ�&��1��gYUE'����j"�/�� �8�Ǡ��>eq^�`�O�Ų�]u�r��?�"D[��2z.t\z�
� -$W�4ь�������(��?T�Bla�����-�ث�vnPq�h�l����_J�6&o�i�����tB�)�_!�� �j��prG��Y(M�4uԳ�a��@�P�tC�	硍���b!���4��&�?�/���y�(=86�-��̸�ao+��f�Z���>�����JB޿ȳ�@켑;�TH��Qn�.��c&�˼�;�o��IT*v�i�	��X{K�. 8bMd;�`��<��ђ��[����5֩]$��Qw�����pu;#U��$��A���ƭP������)�I�P�aF#a{d��c���6���,�����I��c	��Ը:SwI��9\�h�S��Y� !N�^"�7HIl%��$�0�!Ma�C�����O�z 9���Ӯ8Fd�H��~?��>؆k�%a�������Lo�@�@�\k��@,��Ŗ�P����c0�R�]�Ro�4#�n4��u�8�}T���-�-P�/F�♈F��M�XЦ��=p�H��<~����/��`���T�n:N]荵p���Z��g��L79^ӿY���\�@����x��/��eY0���ѷ�g�=����.3���_®e'���`#�F��_쿢���� �����Z=���ۛ�@�
�L7
�A]��3}�s;ղ�U�z��nKcļ�6;��'��$E�Z����7�������nX��o�]�
��5
F �[��h�y�SO�**g^ק�]A������ܩh�{���/_g̪��d�؞<�jL�$�,�����r�<A�������@/� ����JV�q�cy$�R��s_��3G)��؁L�	�~F=M�Z*�&�[�u�^��'�k�������H�fZ�=��ǿ��ٸ�p�-�>.�w$\9P� ��,g�񖂊��R~u`�X�SI�qA�-N�,f�M�)�Ĩq;ؾG��Ҿ792�{��;�kdu�~[0
�!�Ĥ���ΐ�����m�CZx����</�VSX6ǔf�����h[-�6b)�.K<�$Y5rS��#ſ~e�xr��c�hb/��X�3��Y�Z'Vqya�G�@�9�՟�x���q��b�QZ����g��@5%#��C��H��}�8dy��Ր�h��'��� �j�|�SQ����`�j�xt�\H0�^vz��տT!1�[C�A��A��ʴ�% x�JA=P� ����f��#?� �^t���?�M���!�V
�w��0��.��e��@p@��N��j���*��^�Em��ù�lH�YF�޽�A�.:��]�#8�jq���4]9�
��VFl�Z{��o���>�����j��1�s���(<����\@��8�e���.yZ��=1�I&�����s��.�K�)�.�wI\E0�d���Ճ�R��a��.�B� ��l"�-B��&��Ν�
��!�ef�~�wW%*{"�X6yg��J�S�G�Ӯ�������x����F(�����'�,�7`�Q��n)u�͌&U��w��2G���<�wL(m|/��w����/�Jo�H�u$67P�6��c�m=��͸���}.�#scޗDDt)�NjNwM.�J?$Ÿ��SW��s�����yɇ8l���1}��"� ��۱.��=^���}�	���1(f�?,�&�'����K`�	=޻��/�����.w�7g��q�'_ߴh�˶����M��K�I|q۾�5U��a�t�Fj`tD�[Zf'�i3 �b���
x�/.觖m���=����pd���tw='�M�:�"�a������r�(��x��i��C�߬K3��A-�`��~B*��L�چ����'�=�aK��\%��l@�.n�r%�}�f�K��҉�ae�*�e)il����H��6c�)�W�?��Tn*h�?�с�Q�<A{�{-��A��hW�����hR���[������G�Y���z��nwH��Y��3/��ӳYc�H�5��0\f�F�"ERG�����Xvm�г�%Z�
�g�r5�u�j���А���n�M	�!�+�PEI�Y7>��"�Q9"t
u[r�vn��g4���OjN��&1s�2��q�#������"�˥�(�������;3C]�s��'�A#CE�M����Ry�g����76��q���fꆮ�q=Y�*��אַ�T8+�����G��]a�J-H����AEr��^��|���V_r="���c64��J�^!D8��T���"3��6a:l*�$lVZ����Q��?s��jl��CT�צ�뇘�:�3Z�%C��Vb�C��Aw�Sw�'�y�W��V@X����t�Ms��VW�5�-	�ӋCd���i �r�[0̮\�V��G����V,�c��f}�Gq@+��J�y=��]�h
;��������jt��N�R[����.K���DA�$bJ	]֠����ΐ˚����4	�W�^l������N|�ꞽ�����b���80}o���0��߁�pP�,�* QQuGK	�ê���a�9�o�{kl4KE~��7�}ۺ;VH���������1ҿ7G��OF��X�vZ��d%c�K�J��x�MP�d�$Sg�@d��A�����5��6ǠSoBT.����&
� �r��:&�2�I̠��Ʊ��3����U���kT_��`wڞ�8Q;�s[
C���akh&�k��82l�yNK���Y׿61�mTk�jj�e��&�88N��"1{~�yKi1���k�����M�r�eC}�%�ʥ�	���)>_�1~�I�)�ߠw�_8:5�9Yo��GEPR��]S/	衟��f���gth���_�mN(Nq	�IF>E����<R--Z��Wk!d��4p� ZV�AS��<K�����¹PѢ[
f��BȞi R�����ع�1;㿡���<�Iͬh+�>��@:��3b{~��Kw�2\}p��%m ���B�0�Eٶ����!O�B�r%�l�o76H}l����=��սu�ѵY�v���<�<��j��_v�|S*�(�Ք�l�>I5ug���4�M��z�/j�w	 �! ў�g�G�bYi��I<���ԟ�9���zau��I���31,B�T�mu��H��ɞ�pjf(dl�Lv��ؕ�ه3
���� u=�ϥ�����k�����j扽LM�salqH���Im]�\�σ�D8�8y65����
��#�V�A� �)���n�V_D��b��#���e?���M7�ڼ��;�!�E��Ԓ@��H~ x��d]A]�Nɖ吹+[Pв=X�X��6ə�&����u���4�h'���d���6I�2q� ��O�Pt|�b!Nx�٣�����+<��+�%��L�G����k��I�� �����a���-'�?�7� ڈ�l���dU�7 =ߩ5��(b[ܣ��azP
(N|\���h�*��tCw���kԢ[��rXv+��Y�BZ2N�|*��!��c��?Bڛ|�����9^�+qھIj.Ak���<��"�������>V�P��kǻ�G��!���2a�T;��%{��ꟙ��@1C�A�S����Ŏ6�ĳ�>�o�J�g͊��Kch�2�aSk#ђ~�#ޤ��\0!�*��7a�^d%N7@o'w3��	Σ�����p܊rmva����k�zb������ kQ�w�b4#UA?�c���؋�7���?��;�:��ҧ}A1@=�#)�@���f���7s��E�
�m�4�Y�Su�w8T`�E����G�v�d����VuX��)Yt"y���u���C���/�v���~5td[=�t�W���[M��A��`�xVw��p�?����4EEH���	����Po�.E�B�o�&7���6s�A�q���TM�3��ff��2�#�����5� A��u��^�M����A�mD������){���m�g�
��8+��&����J<��ܳ`P��,gm���*�̃܌��S)����救#���á�ѐ8��3�s��k��>�\��#�� pF�0o��?-�@K�Ȯ=�
ǁk����L��'6ֆ���#��5�¼��@nt�W#MZ��n���`H�4uoqx1�&0�X���W�Y��$  ����)%a�}x|�p�7����F���*g��1�zZR|f��k%|LT�P]C^��$��}�''V��M'^��V�h5$�_b
}��L���*�A�h+�;�MZ1IY�e�n�pO����V�&�(�����}��ؘ����H���sg�a��]A�(5'̘Ҏ\6�[c##tX(y�,���)�C�s�;��n��D5������SB�x���ƶ����zp(�֋B� �����Q0^���S�T�f?�(�#��>�o����9����}j;rDǖH�y�)4z�'��̩,E9�F��I�s����=�`�,yu�ۺ�%8� O���p^ߌxCMYK�r������S���1���	�ށ$��J���Q���q%���ϒ���35���m��*V{q������I�51/�/x$��_��_���:�+��͞GTfw�2�0�択��$ �T��ƾG��\�r-Fv�o��7�i���<h���K���il��GFuB��.�Sn��I(hЈ���*/�i�1�k��r}�ڳO�{\�󞹇0i`�a1�A,��˩ ��l��v���_V0��c�[�*���t��R�k�7��p�R�V��i�3Z��Ph������vCa�X\0��y?y=5kL�"���w�@Ȧ�}� Tj ����hA�QF��!�%y����Xm����0D�L&��l��_�ɚ�_���`�	�B�5i��ּ�F�>ُ%�w����m�6��m����8F�a
����@�U!�6�TC彪n�žu���ư��o)x�����-ʁ�AX�'��QdM4�_���c4ǯ���9'Y��l����ܻ�3�'9H*��ޅ�5)뱕߀1d����*�5W$��2fa�'�S6ju���T��d�]��𑭲7�;u�������h���*�C��ޏq=]\�Ԯ,/x�d9; ~��|�]�@~�g��tW���<��_��@n�6�\8�*�J� �"+8/�qĒ8f��fQ���p���X�s%m�ː�<f©T�n I,�>b�Ö]x��i�)�D�ut�^oO�C�Y���
����	^�@�����s'��.�����]u	h`��Z�Og�P�#(Q�)�GvyN#�񟫼%qͯ��.�AW9{��]<}�I��1(-�7!q��};ɿ�2Pt��zO��>̥�_K.y$���z��xC�jJ���Z@~;ݯH��v)b���t���X��`G�7)vlLs�j�6P�;��>{�7����,���������_� �*X���2ntOX��B̗�� �'��ܔ��x^�� %Tʲt�=����\`@)9��G�F8�����MY7?��r=�܌�\շ�'I�}P�Mp0�}���2φ�7s�e1X t�(�9���(t� ���#ֈ��Ƃs}��|�p���k��X��X�f?Rr�P '#�ci�H �+fm���p@�a���ҙ���%� [|���Yw��-I���R�0��Tl����ʌ`������=�)L"iXvx�*���z�0aB�N�9J�%��n��w/�K����f�~�����v���Ef.5�)n��L`T�RO��͍p��g�&-'e��Z} ����q(��ϛ@x�k/|4*���9sq�5�1(��������f��Oؤo�9!8�5����H��x�S0:z���/�\�o����P��B-��ݎ�%�F��!��3���-�>}��i[-�n	H���0�0`��-X��W���{HI���˱���.xބ�}�2-i��: ߨ	L)~Y2F�@����m,qg�ŎN�J�B𗗡
��252����@�ϵݿ��Q���;oЗ�KLV��a�i�pBz�%��U�����#&�j[�!���5�P4P}����ڪSvo�UA ��:��9O�k�U���J�$��y)�@�_��WO.2����h�jg�D��>P�Wvҗ���0�j���+���X��{���>��H�U�G�m*N�b�N	�V=�b�`��	�=��}��r�w]�&J�m�i��� R���8�3i�&���:T���fD���aŎ��_�P��l��8s+д�Ϯ%) 0�KP�y��v�Ƒ�$��]x K��U�j�I�7NOU�h��12�7˯��l����e/�Q�J9��w(�V�~��d��?⍓׵\lZd���?`���sB�������(��K�E�A��JK8��}>�Y�^�!��B ��yʵD9_dd��ߊ4o�]դA,'w(���ྶ泫^*z�4�f����\�a�Y�5h�c0>w�V�5��yǈ�����~�cY���x��f��l�������ΖI����()g#� Z�M6����Eg�S��e
�İZtra歃�����6C���Y�a#�Ւ���	�}/�H������vl,���E��G�Av��h���K�e K�eI��(+��wљ���J/�߷�����ri�N��lX�����O������
p�w�@��� t������T����]��� Q��S��
��C7�RE5�Z�*Saҥ��/*d�<����ѕk�0���V��,�c�!85��>;��dV��o����X���a�����I��b�Lg������bM��1�	�o��6�\$Y)�ΫHɍ�,�G���U�X���	-��"&���53}KŎm��_�� m��d���
��1��"H�K\"[�T��/q��4�G4*i�������q��c?�|��8v��)�]0"��zZ�:W����'eB`!�y�<7�M~$SQ����pM���mV�ڒ��H�h"�u��Bl%��]�@]/o��-G����+�
�=o�x����ᬋ�ђĴ�s��T��hNR鈃�a����A.t�^l���u)x���`+`�p�K]��ĭ�:��k�ʤ+�E�T�m������;�?�����nۛ����wFfO\O�h�t���jul�,�-�>R�Pb��<xd�o��'@�IF�Gz�T�7܇���]Z�������c_�I��H�,o
����d�c�U0�u��h�H% �b�X�7�zݒ[��?ᑕ�=<}��mDn���b�r\��q��1�������gUO����h�^�'�E��cW5D/�%�[�2�}����T��6y�s�P>��"��Xxci�,�����&b;
�-���n�p�@��h&�=�����nL^^�c�;�M��<�%�? ��U�\������˲){�w�S�g�5G)x\��lT>'��.�G�#����Z�����/���������ƪ����$�;&MU$}�������wT����uHe��CL]����T��0���=*��q���74d����rR�AT4�q��&o��a��c݋�Q� �|�^��}>���$���g/�j8�eXA�{r�[�!��,����z����l�����8ߵ��v�&�#G�L��P���ʽe��-N$W�{�����X���1���M�r1g���o���	����]Sf�sC�N��l�q򆒺e�jm�m�x$�B.~v�+gܬ�ؕ�vLd���)$����ǟ$�����⁫ŝ�Vw����>��\�!K�E$������vx]̮Ʈ'��p�|k��U�.r�tsH$��L)���+�0b;�bKTa�S�O�u�\�׏��#�N(/ӅQ��
��l�2gT���\�]!��u35�s���� �.HȪ]�z�͂A�5���e�	w�H���Fm���s�bb7܁��b�&�gҩ����&x�Ot�3`!��'�D!� A�Tg��L2[���н�s�J��L����IB[�JL��;�i�3\3w;�u�]w��b�}��c�$0u�|�n)H�/��n���U��Gp#���p��	�R&/��uI�����֕�	�A�z}X��[ �-�o/�\�"�"�]8h!�h�Fɏ�����]��+fdxa����$�f׵�UYxP��ԟ4w��j���"w�m��N���Kw��O� �R������֢1��h0 Yp�jn,���~L?꩑4�u����;W����:���X#%wH�#w����"�T�6�}���#("n���w�m�5����g��q��H1����=}I��e�<�p�"��zK���Ǘ�h��P�9��Ä���yp���a�]���RpyԔ�:ҁ�Pp���6�ZL��A�x ��T}I9E=Arp$�K��y%�74/������q��4��`*
/ .��@�4��a��k�i�wK�O����`�[�XF�P�q�����a*D�a]m����B�_��5��l��e�A��Y�K�ޭ~gG��p�p6��Fq�u6GE�'P!\J
$�N|E�rΚ��{�癩�?��m�C�4���ݯ����3�e��n����;I�lӞr}4��eQ�k����z���y��nB݃&�k�>���:��Ϫ�&�t��&�e���c�}�M}��.�I �Ё��y>�~�#b�FZ�wL�@gP�l�_^�s��b ��4����NAj�A|?5��������Jj���G�i��&��� ᷓjD��2ި�!��J�5�]ef�^�*!�V���&EiPn(���2�'�+g�÷<v����B|,b����r���<.���'�`N�H�[vc����3������ֳ!�7�ӹ 3/��|���sD�v�׻;5n�눊�<���n�{5�{���S��MWB�<B�h-^;���F��l��2�
FfԔh�%9�J�z ul��g��X�Qt���?jm���=-�S���[�G�?�_^~�ږ����F�"��������©��(!�����W�1��l���Җ�����		�dhyh`ʙ}�]�/���;-٠<�2j���(����AM�)��SP�w8o[6�迎hb<L3� �W��A���s��C�L�Y1�j0Ãr�bDO���y-ru>j��s�:`�#�aIƍ�{�����eH�.HEP{�[�X�(>F�.xC�a+P�ŵ	�#w���f U�;�p<o&��֬f�f�^@Jt-�!Ԛ�i@3la�&xY�>�@�id`�؉�TUC�p�e����&B�������n�E��é���Ȓ����0��#cI���5���0��RD}�Jg�����#�����W�-7�0���vSJͩ �����#E�������d��P�oR>t�ǃ�&��KU]��������~�e�"GEV;��F`=��'kQy#��F��"���]=�;IA�5�D=�Y���AA��q�� Q|�c��3�$%�;�/ݏy�A8�k����q���p�C��R��q���(�xH�8��;����*�bz�m�YF.U3P.�E��=�r���ɹKP����\u�rŶ���L4��?��X��Г��}~�a���1]y	��G��U ����D��U;9�1����@��5C���5����+/�F#�#/�̜#��>Wcj�f�ⷃއ~�k�s�m��4T��\���]['��#�״7�C�P�:�N2�ץ���YdZ��V�_�qe�VC8�jw�\���!؄>�(:�"U���[�?�j�<*�Wm��������K���x!��+	�'`g�[�J����z7?`5g7�uOk.��/S܄i䶝2>y��A�hv뻢�J���ID-��Z��o���c�u��RkNyx&�8-n�k���h�Q��^�H��c�,��z2}�M�L\���=�	1�Vb�<���S�?�_��$�C�:��dV�6��a��#v��cn)��=˾���[��E���S��1��e�iFp�7�1$�^҇e;"si��F���3���̠��}������+p,�T�s^aɏ�����?���^40�Չ�)@���23:��T����t�����z�b��w�^��0�9K�~�Dp��_"m�\EN��UUH�`X7.U�{wa�-1g�${[Y��<�����R��rX����`0�����9,<���ͼ�N���(��W��b�j|t�!�������"�t�O�?�ඥ��3u����[��`E$2{���4 Ԟ� Jɖ8��˃���'k�w�]�&�g��|�2֖��I��L"�K�����7� �H9^��߄?BEFU���/c_��g��q���A���ǣT���pC\�?�Hg���^9˨St}���QI� �ʫ�&˻ �z��b�#����lw%�����PM�3��]�u���I� ���Ϛ������0�ٛ/�Cy}�u�# j�{YmWb���2��~�G�R�|O�jZ�zo�I6�R������Q$~Gu���00�W���	8�.o�+B��%e�\���%�;a�V�Jo�1�*-��a��N��L��_����QQ:��C�w"��'�ٕQ�Ĥ���@�nmp�;[�s^��}~3Vxxݘʅa�h-i�J�b���K̶�*'�(�sdBQn�W,��C`&���Y�zN(�P����\��a�o���T�zyk��[5�,o3�B��Q�lU d�X��e����dg5z'ו�j=�<�r��N��H��̐>4�;��)�+��yU�L�Y�� ��M[Y�1���+.F%O5�P:�h��k�J�D �Y��K�$f���'D������~��l���@�3��*\ån��z�`dJ)�|V����O�L�~:����Y�M"t�WKא���� �P(����Z��n�u��OSLB)$���|���P#�KBڷ�q�*�;E|�{�h�%e��s4�W]ϱ�x#rA�UNv��02_N�V����M:ҡ������?��g�j�:�r�%����
9m:�թm�f Z�v��W�o�fͬe���I{W�Y�@�R�h�����y�+�!��A��\B���Di�y�T�m��G�E�Ϊ϶�b� ڗV�S��cT�Ez@��������./����*��
�*��C�G��n����KW)ޏ8�*G�?խ�4������h�g�R'�qpO$�+��\���f����agWm�504xM�|�x�zZK?ǒo�Y�tj�\��,&���s��&��.���>,��Q�=c��a�9�L>�L���&7P(�:[xHo���I�5y���ئ#����z����7J�VR��7�?iP���1l=s-&�.��o�������:��{W-�?���9���Mz��P]�㸙�p��6�(g����� �mؐ��S{�,��@�q����զ,�Q�j���*HW)<o���ȡR����2����%����{Fnx_��^ }��;���@M�rp7�0O{,���{+6+�B0�|Ϊ�7O�U�7z�Yv���K�d5e��w����5�H�l����ѹod���ih�Eh�ǝ��Y\�3�>�V��a��[�7Y�l~�}��ʤ�qV=��-������7'�F4����@�NWv�K�픋YG���ӌ��NW�|���t1a���eEV/0ha����@c��X˪G������<�.`������}��X˝�v��ї)�W飰��@hJ��3J�b��щ�kR�+�b��Q�0��;_Nt�B��k�l2�wc�Pb����P�YQ�6W��\a�Ly��z;��mg�#1b)��)�e��1fl���&��Q�����Y7�s��Ǹ�$r�IF�p�P�j.��&��7�!b�i���cA�D�e���a�d�r�f��iK#D�}�-a N�WJA�-1�v��a�B*l�	L���4wb�)
0�jR�A�����G HĖ��"�"�V� ��@��0ђ�P!�� �>����<�82��+�Z!�3�x�O)*�s�Fu�G�D�䝸r��w%���);���n#��r�{�i�yt�Gb�[�h) �L�������ru����|7Ʌ�!����^	��`�n��������õ��Րq���Rw�[ͷ/bι��iZrt01���4�o����j�k변A�-u����:����gT�r��W͎�����g�U���^���>�X|�N��U+����y��qi�3���1�!]�#�Ą��Ge-�������':(�$��E��i��RC��C�w�Q,	R��2�'?��ƍ�$��I�*�v��"���WJU0�{�Ҕ���6|��F/�3nUGjK{�ZI�~�k��N�?�����|���M<z#�8�oG�y��D���1c_m��-Y"mD�%��o2��iz iLkDrձ�PY#�ĭH���!T�����k���v�6�	��z(�Df2�;s�r�b��q8�W���t�Gv�g�M��b�0 7!���J�����-Tr� ��ʭ{��>�p���o����&�sJ9�MH�w<DHW ��)9_�*�N��2pit����Ӱ����JjA���y���09وՒL�%���MǢ厀�I�z��Xt�	r��=��n4=ٶ�HG("�\Pf��:p s�V��,*j��2��Q��2[����0㈄c�$��<��W�������ݡ�YJ�a����d²4s���A�7碌���o�^��\�v<�ɖ�,�ziL�vpqF�eLd�G���c;jS��P���TX�Xo�X\��Hչp�+�7���B��J׃'$��.K���S^3<�S$��[r'2��	�J�����f��j���7��>��ӃI�����n�ہw^x�� ��lrc*vnW�Ê��	�8�
#�A���Ƕ��k���U�1;x�_�\?�}x�i@�!;������Su�(A�H����T��i#�q��V��TY�6�K�����}SU>�����uH�(��l�������E����`���H���N?I���X�F�S_5��:.ĕ'#�R��n�3�{��=��K�3��7CW,^��ǘi�m1��iŀ�k��z��Ô��q�qM�#�(��L!��nl����I�?{6��t�{F/|7��
%��j����%�@�:4��g�P/���~���Zٞ�v�=̙��<͐��'��ό|����U��>.�RV0-k�3kc� �͠�P��`)/�����jY�[Gy����6?���� �K/��._%�&l�k���4���a�F:%}��f���%��A��zk)D�"����na�R��cd��P����)*�RY}j�C|"ָ��ڑ�}�(��('1�$!�.�'X�K���^��8��E���e��.'C��-�)[�]�Ju�yw��v��[ՠN*�((젃7�/�/���E΋��,�Y�S�j4��6z�؍���,x���i ��C����� �Kp�3<�A�T?a�_�S��u0�o�����Y��mcŊ��-u���M�bO��R��,]'1`��D�����Uw4�d9�f0� ���k` �. �-#�S*7���`3���UI�~Ǟ���;�IA&�������kA�u/����H;s��M�"��u�_�:\������	�'�`�4F8w��4K��D>�@4�������8Hp��ry�C�~��u�3�D�?_x�8��j�9�a�G)^�P.E����؈]����#���N�rK���������9:�γ�aZ҄�m)"��u�����k�8p/�P��j��h�fE4 �0�8�Z���ӥ����K�e3e�M��3s��N�OkyO���<�[r0"���	iv��7b5��u$��Y�9ck���xᙥ~eӃM�E���_ذ[��Ƃ���T^��z��C����˵�|�T�B�]�2(g��i$&�A��{�[��G�-�z����?���`�[X��bc�����BfPh�����2�_G�%�ջke���WMs?B+���q��藍�*���u!�7.��)��6U_�x]yPK��1�����8��]o�D���i�n�ݵN�yT���ٺ���N'��na:a�;�R�|	;��l��E�&'8�8������k�yؒ� �����h�����ּ�����b��|��v��5Ҿ_����Gm����Z�0a�c�WZaneq%/��͔Eş�g�FrۍecHR����^��j�=/���nNu�E�O\f�Nzљ��ձ�����dA�	C�Z�O��r�u���
����[S�Z��0Xkw�n�ĕvt+��g�����߶�1��qJ
�F�!�<�I�O<նx���9��V�VR��7�]i�Y<!w�G�=ˤl=�_D���mwW@Nj�YE�>��/ `DG����aCWID�{x��$k�=畈pǟ�@R�)�t�u㓣���3Ѻ4Gп� �4RRƁ@ o����1�������q	�p�l�x�ӯ�L�x5�����ҧ�� ��m�hǼ�c4��1p5�R 稾I���~�x�A�Ez��}!�C���T� :o�"Nh4#@�ї��$�(
��@<���"�UI��U��b��R����l\=l���C1'R8��3��l4s�;r/�<�J�
W���.�is`R�)\il���!�L�ݎu1�H�ڀ䗻�P��6V%Z�����s�\�d����K�d��9hQPf�\X-��D1�@)�w���'��o�N�X\���zS�mH\4\���zX�Z�+$|��Ə7 �-l��):���H��}?R�&���]n�Y���A���?�ɭqU���*Ѥ��O�*�	�����}����p>����������@�b:\KĨ%_"�ANㅩT�k�]E�x:����ew!m����	Wd�ۼ��j���J���'�B��ƎŒ1�J��VA�;�Jƃr`�Ցr��2�5����1��ABG����y��n?�,m�L�[��0�i׌�6�zS�Ś�x��sV�N�	)l}�}�U��}�N^̣�DTI^�V�稀���V-R�&D!���4���F�J`�v���;����1a���C@�$aR_X�C!HfK\�U�~g���\1�rgZ�ϻ�y.��$�.�^��������,�T�����憦����ӿ������'��m�&�dMY�<+J��1�5�2M�㋖leo�+����g���Գҕ΄q7�zu?D(1��k���r���'f�al#t�}�;c�GA1]X�R9�uT��oj��NP%���m��[XA9+l���F�f�s'�w$�k�|�v3ͫ�g�	���� ������e�bq��B>`�l�������b&<�o�yٚ�����xd��6�ëC��Һ�m�3 ����ͩJ �����O�[���w'���Et��-{��	�~lv��4�9���}o*@�����,��h+ڇ�ƞ�s����>�샗��M�|�DTd����4��%��&�V��C�#^����:s���;!��ާ�d����CP#$gS��#�*g[���鉶�o (@Z��
V�z1�xa�2`�����/�n���\�'n��o�;���[���z�y) ���4�>��D D���#�z��]WS9���U2����!��e��}p���ӄ��?ũ�R�5���-��߇S�Iw{�O����x�,�ݰ�rX@��<�(�v<"T�3��*����2qQi���(�e؄M�~����S�#�ˢ���g��"j�:��)Vr�lVL,�s�-���}�^
� FC��G�5��١qF�z/.V�O���������׃�g�|���]MX:CU��}�5���O��c���.<Qw�-�B+�pJeSTw+��)f�.�ZU0[*T��Ot�Jn���$}���:Fr=\9�'	�H���s}�6��� ��ѳ5���q3�L�zL��F$����F6C�.�����skq� �q������{��K���aQ�k'$"�~��ϐx�K&j7��p�L'Yga���۽���c���ʰ�$V���,g�5ٽ��4�������}�J$��4~2��Y����0B��ߞX#5�a!���v�s���BO����c^�����sa#���G)t�&�m���Fң̪e� s��+��g��G)N��Ni1�gh���?e�G��'�
��sDzv�n��7w~
O9��,�p᎑�([$��,�갫��%�S�&s�#���Ǽ��ƙ������Ω��NZ]�[��r��$�<�qf-�qU�G��Hư9�bU�a�Y��>̴��J���^@t���D�K ��!z��/����O�'�ۇ�އ����Q;h���.�wR9{�$.�����cU�x�y9��L�9ō�aZ�T�w�����A�Q���a$�k�/���e�P�K�ć�"q�oUYE�
b���4o�Q6�T�x%hw��J� ZY�-d�(��]�L�wz�0zR��LX�0K������[Y�e�i��W&���#� nG�*�s����0�}�"��n��$ֵ�����{-�[!P�C�^6�r.ǖ��`]�aʦ[�tl���f��Kn��@	�-
@��5�\��	XU�'\�t��ct�>�$�Z�b�T0�0�a���^j�~�e��lTW���BH*�U���;3.��E�������L�|�[�u����4>��U_o}�,���w�/(�;�o����z/Q�sq[����v3v|�E;v������@z2����\d7^2�L皧� }TU�#�����p�b!����a���u��~�g�3k�?�&���Q1 ��s�!AE?:��'r���Q�6��. F��l/mę��\ʵ:����ս��Se:~�2a��4�rc|.�H�yg��Bګrfޑ��6c�h5�P�j4p��k��5\>�h����z��<Q��-�^	_b!vR�H��}MІj�wo˒��^`�h"����׾�w�7���X�(x�x���vB�qEU����}���ݣ�N�O��[7�w�ש}"��V"m	|����i7pJ��Z>�?Յo6�����8���,��>�h{���q�k����K="�����]�bi��N�VC78���1���͵tϪ��0���2�Iۏ�b�;�|hh>��NٵA��8PGw�ya��[�{�	�_9��	n`��LQ�'�A����C	ر��ᶐzK�V\c������j>�Q���� V��|�_역^w����<�LW ��QǾwZ�=��@����%:���%JQ�-~����2aq-#Q������i��^�3���O[D^���0A�R�:�/���q�G��R�N�������5��ף�3[06+�{�kb/ET�B	��>S�-��'��$��[&���K��u?<���p�>�V�7��C����Ik��rh/��W���q����z��_�4�C4�lj�F��0V�:����S@����Ck�i��.���3�:&��lڔ
�gN�S�L��Q�	��'��A�ڡ�o�k���p<s!>{��(�q�V��:[#D�l��k�e����!w�����	y�hB��k٢�yX/�r�_ܥ���L?v�"�0�)"/"�#Ԥ�o똲C��Y�_'u�2U�"G�y�X0.OJ�;�V�ӻ1w�c�(�٢��\O�W.�u���̸R/&��V9ld<�����o'���7��oC��X�Aa���<q�~�뱦S��6�8u��w&l���%�̄Sm�K��œ۫M��~q@�߈(x�|��� ��T�}�*�/p�*Cv�L=n�w0��nP�Y���t6Ҹ5���@�a,r�1u|�LrC1%���W����ˋ@�.���*o�BI��gw��x�HN�V-M�zN�]jj�Yc��Sa9[���X������e�fI�Q�����=��=��ؤK�67GW�@s�G�b��D�hy�%��r�tt�	ή�L�{�ε�+�Ҳg���if�EnQh���y5�w���3 �/.J$8|z`s�"lJ}���>n���-um�ɶ�5 +.+"����ی��	����O|F�rnWBg[�E�>[nqd����* ����ע\����-��gi���t ��}�-�-��O\Mc��ӳm������a�2bK���4�#�CV|.U�N �V�S0�Za;����RzM��Gy�Uw��-Xs��K�m�������x�"�b�+V<G��[�ՠlq�{�$n���bR�\'MQ��J�;?Vda���୮wslZb8��4�X��r�ybS=�@��C��0gJV�{Q�LDD���w�P��J��j^Z�\�"G���>�6����{}8���̽��Ӷ�T���Ŗ��ֱfK܄!I��Wg�C2�jm-q��^AJ������]��^�Lh*#�f2�M�`78��h���v�}��B��LX��5��}<���2c�T���RQ� ��y�R�r� o�:��7�\�a�n4RV0��#�����qtX��\������������(�?:ju^{`'�Ր�>A������0V��֮���s�c�"a@l�H��D�L�&9b_�����ȷ�K��!g�qg�R/�Y�6ԡ4^u}���tG	^��Rf�P������[�"7bg�Y4��{U�(E�h0���<k�+S1Z��n��Yǿ�j}C�o��!\#Le�6���:��~oԢc4W��G1�?%�w������0,��f�Cv�܎s; �?�}���-�hSH+
;te�0�� �^M2�M_h�����?8���{�9�CJ�Ju�>�v����T��?���g�=";1 ��O0�%F���Z!JtyG�+ޠ\�"i�b+��P��կ�&�r���ƻ��S6�q�ء�L(�����"�3�з'�BGY�|�j���~��W�>�6S�&�mC�u�������ufO��HrQK`���M��"�C��U`�g$�̍"r�ȂM/�{i �_\CT�n��A6
�y����%��?�es�Xc��%~p��e+�_lO�}���w����j��D+�И0��WM9T�Q����� �3�$�ʌB����P��ʓ/���g�=bj榵<��BvF���w[�(�C���_��*�;��S"�(�wN�3�b��r+X�a�������p��M��ڐZ����Q�E �c6� tI�G9~��,�D(�%��I*��~�qI��G�d�J]�i�����*���B��暧\�j�3��6Up���D�<�sj�Bq��;��}y>�h�Ԇ7K���tC�KI��Ȓ��@��`Qe�/�@=�a�y�c	i�D\�H�>x��'�ȅ�3P7ф�נ�A	��}�i��yT���Ɏ,��\���k�?u����+Qe儅��%� ��ײ3��8���և���O�{ˀ#1x�Χt� `rb�e,R���zZ1��[����&�������s�:�<�;WBq�����)akA;O*I�e�пM����v��	�wxe��6�VB�Jǀ�Lٷ}��ΫU�Z���e-��	7� �u��ǋ���׌��D3M� K!*>#�-�"|0����C�s��(_)�5�k�e�W�n�ƏlAn�o#C�fV�#�ȚFQ�B�җc:�������]��L�]c���;?�,ԇ �����/QA6�G�h�z�Q{�3���D�2�7 )X�s�)�Z���J&�nP2Q��>��Ӧ����!�*������%��m&��K[(G�W<�]�*���W~�s�aB_f��N;a����B$���J�-�	�C��-ۭ�&؟��G�N�����iC5���7�x�N�~���M7d�+�/4�Y���Y����A��ԓK䙭�3���L����ORg������U���������l2-@����ֱ�+�Qԃ���5d��&-�ps�ɱ<��@�bp����ҍky�@�P�2۫�͏T����5��.��GȠ%�#�I���+�{�����[x�e�f1���7$���GtٿCr�����0�r��)��Z�n�c�4e��I򇼴V�{�H�#=�J�?��5i�;�ga�~vf�fEh�HoWsF�Q��#�N��Ϯ,��<;���Sfs�.����Ոl����r�"�#x��u�^�2�Q��0�PA��㗇���@����B F'��s{�=�͊�,Q�����'����L����h�rc-R�&�~y��cՉ��E>d��T��������˔�}�I�
����Ck� �P�΄&�3w-6t��h���h�r�d6��nZ\ 08�Z�)�_�y�Z�y��	 .|�Wz�!�#�v .t��'�6fT?�-ם�Y�0;�JH!��1=���N�^�|=Iy��T?���k��H�O��9]!��R�l�&�J���+K�"����j�r_s���Gb9�j�t��LƁbڮ�Dq1_�(�aNA�`����\�u8��yT�ӶY�Ĳ!m�}�Ĩ�� o�M�����ls}������rw����70N{O�-�F�/|n�l���5",�ZrI�v�}u�z��N�#�5�$�����?QCH�H�I\ �y2U�#��\��jP2�����&���(.TU�%N�}�UϿ�Yri��U�����kE��/j���h�O�w��o�T��0)���@)jW`���DXp��`sCb-��K�����2��su�'�᧜���!bz�V�2�n�_X��h��m\��1x�+�C@�`�sJf��ў����1��/�7dAs����vwqu��;��b���כ��YWH�T>�]��:2����Oݼ춯��o�N��ڇnt��f���6�`�pbm@��0� c�$KK�%m%�	��Oߞ�
J�B���U�@W5WF�<uX~qۦQ^�t��q�A�]/�1{��Ʒ�����+x�q�8eTu�F�:�'@�����ѡB�	�/l�T��˶���	��n��?/,�l��=1$̶ݑ�yL ����L��WW�b}�2%�����)R��5J�ɲ�`]϶"�
YF�XX7Y��s��&;�85,�m_P�X�z�������>����IX�ꐟ��-d�<,~7W#��� qE��@�dze�d���08!p�Q����Լ�-׮�f����o���:[Ԗ���*���#1WsgG�Zy=�<�o#����+��(�l`sB,ٍ��5��wMIAA��9;���<�O�kd�f��G��JoX�>�N5��^W�j@�y.ƱiKj�2@|�����T�]��k��B>t���бyz�|����ť��2��ȵ' ���7�7ɨ/�t�S�E	��U�U�*��?�Ǵ���UۆOˬ�A���Kα�L0l�B'�G����o��i���R~��fI���/�E5�Vꡥ��M�f4uq�C���}�c�5�|���T�\J�OTYm|=�ң�=��ݴ��罸؟���5�6�R|�GJLQ���i�U���~#���T��m�r���w-EkZ�ըv�D�}A���J|�#� K�Xzǖ�����h�{�K۾b"l���W_���#K͎�<�i*�EA�m�y���<�e�F�m�K{���՘��Ŝ����7�o��Z����ت�.N�� E���^$�F��,�-V/��B��!#�G����	W�w'�>T¼�����1)y�Q�1�6�$�k��|(��	-���d4)��8��!��M���<3x�,A+�����N� �ʈ{�����z8������g�e:'�$���Zm�X�����Ɔƃ���o�˱�}8�� �q��>�����z �0��f��p�8kh�)لk�Wi��tv�w�C퐈wK(��4����k�|�ֺ�/�%*���;{
�M�}���>�H��JA�4�i��� ,\̮o�Z
&1Br=�/����:N�x����$�O<A�#�y��c�j��4lN��� �.O8n������5��������G�@�2����Ng7D��{&��T��§+�`}�T��A���l*��E����<?��r�yo�7�k�cM�1!
�Ri{4ҥ�q�_�"T���H�kwEg��Νvr�wi'�˽�a#�xℼ��ֹ�ƘO�RWNF�9��f���j3}��O�0n�l��jg���c�
��ǯ��ѥ���ˎ���6��~��LplQ)�n���|UmXӚ g@H(��<�Ov�s�����J���0梌�3���:�Հ��0�����n���l�� ԉ}��C_�,��.��ɝb;Wd$WĿ��Za���g��$k$��o_����<;._�T�Cs��lC��B�>S�aAe5����({ᖅb)��>���t1/��"ɸ�e����=Q�~�D�c�=�؇i�т��і�ː�2>�����x���F��5;e\��NѬs���C�DE��<e�Pc�_X��+3jһ�.Qo��]������6��ɕIc�q���V��}��u��k�Wl�k6g*�S"��߯��UM]R�yם.ݬ,%��h,����]ˍ��B���G�8D�޸D�^�^V��O��y��	���_�:+��|]y�N�.d�<(��C-��'+���9�	4���v4��<<��}JHN�U��'�v����O�hs� j�>¹�n��x�pu92L��	9i��j�!;�8Y����:^�"��>�d�'����Xs�b?����7�c�V����ٺ����4�%�\p��{��Ҟ��1�&�i>K��5����
���1���Q�8X�y�ͅ�5c>�s*�1`2�=�{��w�<̜��H���ŧ������ٝ�	�J7�Ig��9h�W�H�[c���H[�{��K�VUB�)T�G�g606���ͩ��{OQ5TRT%�[�p��BZ��5~!��VZ�~�R�8��%K����Quh���eF���,oȾ�Or����ݐZw�Ppi>���<˴��%��do��]JlZ$Ռ�iғD��k�wF�ey���X��48ʡ=�n9Ԁ�ܻ�v���Za���!�遴�c���q�I�������4%$N��w{&�>LT}� >X�-A�x#��J@kT�+�E��v	b����jY����6����f�_��j���a(�D�uR�RZ|{1oJ��֪�	?�A���]��k�.�sP���*�ل�|�@kM�{�K� �8������;-i+��� ���a���'��k��W�x��Abb�3N���>Kv�&�x�%
��P�
�7����[�(�ȓr�䛼]ȄX�v	 *Y�٥f��5�Z*�I��8e��\�I��B0�`�k��	�m�$2�o뒍��#	6��Xaw����&����q�ҝ5PB""cT@�;j��}����n�l�����T���\�{��L`�W}���8pksY?0XF�b�Oc�q�D7)JQf}�	�:��l�����ax�qr=r�E��<�Σ��45�I�vӣ�/L���&~���l�9�I�o��<���&��1��p��kU�V�(Pq�e�Z�e�c�l��ϛ�Vnۖw}I��O7�
���I�4Rk�e���m�d$��P)�5�>��R6j�_����A1�Ջ�J����Jܩ)���G�D΍R�b�}�Y�>���D��],��ș�Kߵ�Y_���}�w�+4pWݷx�1��ɱ�]#�e�&�D/��`������$j4�
JJ�E1�Ͽ\��*p�~<FT��â�Pa��_���9�e��Sf@Ysr��az��p�:�K}�4�Z��Z�w�V�����Hz��pf=���N��� �q�����kO�^g����wHZC-pR�9K�ޮPA�Mf�.ì�g���3����Ou�&W�jj��B�Z����S�x{���v��w�X�˼?�D��@8�G��,�e��_��s�Z�
m��'�Y(����]���J�s�R�	-�6u_�%�4�}�D����o�B@�*�� ���m=s.��",���$�C����V�$C��h8�Ի;e�ɪ��o̭���(Mƃ����Q��O�����V�|�I��m�:S��1�^�M%�N^�7��b������A��D�W�-W&fF��&�ʌ�T�>1�MV���忕e"J��!?��NF|�0|��9��/'�����8���A�q���Ⱥ�2�L����܃d٩�hr~��Y��G	�/bdi�w�y��o"���Ц���!����s���3�,���] �PĬ�u��U؄0��2��H�a�,�����s2ЭY�c1h�83 2
ʋpO��up�)�>)�I�P���ܓ[O�A��|��Xm*�O�!z���6[;�d�/��]l������v�?<��&�:���h��)��۟�E��IS'��Mw^�*\�(~Ng�c�+H5r� �P˷	��s��76�CN.o���,6�_��'Ǎ��)��E�]%9������D�ZE�{jݜ�޺k�&L(F8�Z�gX�wi��n|�mJ�����uy���E����e�9�s��_�!���"B�y�P��@͡�1m�X��-�V�@W�*�e��?�/�������]��
�����]s���,a��,G�
��D�%M1�R�Q"� !]�=��ȃ&X��9�JZ�e���c"����UJ�z.v-�@�v��7����"A�?�߈�TE�8��oH��EC��6iF��q�D��������M0k�s#��w�+���6h��"���P�Bu�c�'�؉ÈU�ӬSH5M�D�p�w�[�O�y-�4���y�Aކ���P -K +��c��β���B���#��w��@����?�׊aȁ�]^�JQJ"���q�]�$�/m�#S���B��'�a��2u�v8ZtiZ�E����((�Zy��ퟲ1�L:oa�Qx�X��u�=ES��zC�Gr��j��=c�퇀@J�}��o�RY�i y@o�I���ѱv�����?��M-���]g��jR��9�� �ʌ�m���9�F�!�����=�I�$i�q�/��:{�kݾ{V-�cI��ukHS�o���t�uT��<�$������Ё��ǁ��j9��

��"#��,ȼ%{�s}�t�6l��d|���o�-�^�Kd_֦��A�T�3��������#\�fz~�≹�ӝ|�A��]�`�_[9\}1��`P����O80d���;ȭpC�)���%�TcZ��X-��m82��4{n�u*�0����H�~��jt��A��P�ɡZ�ݍП��J�/�D�	�I�;��ndH�

���9��b쫋���_���d��+J����k��%�-�-H���5���s��n&ѥ�+�B���Vj|�|�Aq/rN_�}���)4X�AПH��X{W��).����*�h��aN��!��)�Xs�{��I.p:_�9�D�Rw?�-���|�d�v����Q�+�`�S'�&r�Sh�}��'1����߉B�u9�չ#_���/��W��}j��FV%���7�4�Uu�Ls4��N�W�A	(�Y���+��y����:{(D�s㦏`軝u� �
K�9�?��A��a��xA@
�W>g�A����_��M�)پҥ�+�(XƉg�����uN���F����лN��B�#4�0�Pᥣ��Q�w4��Lx�T=ˣ�v�!iuF�c��|j��j��^)�߿wwb1D��sԴ)�,��\���Z����\���\W�߶�����������>3�p[A���R����K�-`�9����|��n*-�{W���{?Y��$W��� ���<�F�Cb@����?cm�^}C2Ӹ/u�V9��_4q�٬�:h�X���N���nR�K�j;�Bq�d���e�-��;��{B]�vNo�)���S�H �kB"=�c�|�G-ew4�:��x����)��=�x��0�����OmtN.����Kx������.8����f)�TI�>��~Ys�F��Ja�m���W�=L��p�S�H��@"D�xM�f�nT"�d�{���V�� !�ɓ��-u�*��$/5\�'W�^е*m�jo�� �]�;�E�G�J(NG��� )�ft�}DTv�1v��N��a ���|�U��8׮�ke�T��~�|Q�I2.��T﹔��T<>.D�fL�O&O�����$ �.s�B<��X��+�I?\��a��u�����|]3�ǽ8��H��|�YD1W#�G�r3r��L'z~:#^��Av�gي���(�ȇ�p��t���X�ͣ�Le�w���ms��m���(���r�i��IJ�/�'��<�|M��.����?��2�NKv0{��	��R���j�@�Q�a�^D�TOhx�/�L2���Bh��,8Κ��d��p����W�2g�I�����zۉZ�}���S�+:��=����� ��|P{8����"�1���\����U�u&(�rN��ya���p8����%�r��0nRe$E�0���.6�ͻ�.ю�iiо�W�|/���R�8=�P3~pԜ��j^u���)8%�G��|$�E.ϔ
h�k��5�P���y[�Ș�4�5��7�|~G��hB{K��i^�{�sAk�k�T�D�]����F��E2��Tb�c6��vK�1JB���ȑ*ĪW:o�A�,�z������B����@i��]��Q|��*�r��}{�H��U xc<��i/�l����	"�ɩ�rQ`'����{��b.�_+hN�[tz^��y����U��/�6�a�@x*5:���:����a�ّ�K�ۛ�J��s?)G�l/�������������ҺS`'�����rR�M��!�ٶ�����Y*�b �{�v)U���
�s��&�ۈ܄7���'���N#݉�7Q=��T����҇���9�q8#��R�<(ώݹm�pVT�!A�.#(�2L�YԷ��NY!uO ��A��e �y��t("lk��'�Gφ0"�DN��>;���+8r�5ˣS��6�<����`72q�)�������~�b4�kU�%�'���엧��>�j�b^#a�I�=�����g���s@eO�Y���bdt�3��p�m����vq2��q=K��]�sܘh��r?���?�����aE��*�m�v����D�̼4m3�>EŘ�@޹ȓI��H��� ���l(W�j[�d2Ӓyo+�8��ח��0���o�G�U ���H%�:��t�A�o�C|}��Z�ϱ��f`^W����$貮�Z�}��b$D��A�+惚�
L� 丽!2�jzlq3M��	A�M���PO/S�'�[��YJ0�#É���q7	#/�9�[�'�;F'�-b�N����W��3��i}Td֩�wE_\W�0E4��-���%�u������<�5��İ�8]�h��U�V]�Vq���i�� ���Rj?�j���
�P�.��Ɯe�T��-Ŀ�Êw�W;��d��~�,��v�Jr�_s/}b̳�����sAc/��b�2ٗ�R����<O.�4nc5s���p�g��;�����'w�7�lD���0`Ej�?�5��m��f�^|���t/�Ѐg`]���g�������L�A�M�C�F�^������+�]��P�W��6�H^~�Б(�#�C�'s=���)� W���z�{�'\{Z�.G=N�M�`"�Z��J�����,O\/T�!
^�<��)����c�����v�:"\E״�͍�(��*���A%)��eS#X�#Zͬu�qOrG��\�}��Oh�4d�FKBA�Z��Ŵ�D��,��2�w���륯�d�Aꯠ��$�M�{�ШH��u��\�� ��.U�V9�Fx�U_d6F?3�L����u.��n�<|Ab{��g�lR���@��a�2� V�^��_�9Z>�I��"�!F��j~�>�{��>p����?#��S�Rmv��;"ZS�XcėF� q�?ӡ�R�!���0���^����eTN~��������W�)u��ydS{���ʖ9X���Lg��
�f<��21ۡH}zmg!�z§;ۓF��F.��H����� ���꥝xb���P"��G�V����CbV�?���A��Fg���H"n�+Z��pq���{��e&��J�˳k�3��a�=�N5��n�+�5����aT2�;gd�!�i+[Ғ��8m7I�3�cシ6������I���4�{�����u	���F�QUS(�������_��p���/�[���_�\e4��]���1,%�T�+���3v�-I�Ǭ���E1:>._���u���%L�u<�q�g��oTp�5\��l�чEj��8A_�x@������{��_O��=���MI����'�?�*R��?����#6#c�x�.R�&�j�0� s���&���P~SU)�{AZ#�F��(�EC�&1�Q��^=`�#J5�w����o�F���{	I����jV ��r�%O�e�0��'P���z(ćͅ�F*]���lMʚ�i�!d������$Ԁ�����7�38��^*m		���z�ّ�s���_�]��0�����b�TkpT %����{1w��/���Ą�͔����tS.�Lա���t��Uq,)�N�q$����q�(yqŞd��e��g@��/C��5
����qo,�|��g�9E�ݧ(嗤ڧ���:���~�c �d
.4)g��r�@��L8S|�9�0<�S��߸M����ԑ��Bud4�&$����ȟ^F8gWW��qV��gG��!� 斡<|�����!D�b��'����hi+j�ٞ'��a�Tu��l.�Fʍz�pm`��K�c��F*;�ύڧ!z���8�+�j
�^?<�
�!.?����}d\h�M	���	Au����X���x�0�waP�$�?%���i�¶me�(��6~��B��ܙ��$x@�t��S�X��F*�����]�\�́��(2��χ�˵������4�;@�fQa�a��]�ǚ4Y�W	Pt�fd�����hG���4Pꑜ��!��}�%��U��d[�aڬ"2	=T|�~�/J�2��ACF�lW��_+׿���n��{�k�ȶ�d'�i�MH˦̒�3=�(����Ҫ��Ә�/���u���+��+�]��!C��Ǒ�y�=6��9���)~@����l��尌�/����wx���q���F���v���#X��d?��qU<b�Sm�)���P����̲��%���A�:��;ü@ �`q��{0�^���Gb���#����<�ّ�*(�epe�td\������
ț�ђ�U�I�� ��F���h+/�{ie�Z��?}!s�� ׉���H�?J���lz�e�Q]�����t\�*�4�]C�u�YmV��҃�F�܁�������
�!��\�i���������®�x%�Z.NwQjkB��M^�#�+�O��Z��hH��#^P5'���{.���B$Am��$A�B�SmȐ7>��8�{���E�>&@!g1�Is���]�]f놰�U��B�����}�Jhȭ<�%��S�5�z\�Gp7�)� O�IK3�5�L����۽V� \���������2fH��b����t/vc�+�!�?�:7�,�{�y��2>����U����P4In���c�,
J�U }%3�D{c���hz&S��@���_&7r�C�Ӻse�L��[��Z8�!���6謾���"~A�Y��q8��3Y�c:%*~W;��o����N��BLX��W������֛�����^�	�3�]�؍g��H�B]�~����Sv�s2d�H}_��������'���>�����@��:�Z���e�I#WM�27!Y�<���q�-�'bm�S�2�rmv�c5�C������D�>��4zY����r�q=.��:ߌa�m���~��#ؖ���Nw�J0�f�V.�(�a�� ���{��`��Q]�yBڨ�Vz�4�� ��e�(��nO����t�m豗� ��d81�𲙓��N�Wp��Y(.��[P3����wB�T��g�n���QHT�չ����[���/�{�����{�qz,P\����M
�\@�;���X�K�M]���V^)���x��j��}�/�,/ R	l�~)���eȤ
����'E�]���;r�!�(��.����њ�#��o�Pp���Ɛ�FV
\�U6\�U�}�����L��攫��J�|��?�� ��R�F9�zG'R�m�$	k[<�v��� �R;�T���r��)��zd�N������h-̌�j߰Xbz2�����!��M�����a����Z
�@eM7u�,��c��ׂ��6=��M��Ҥ8��@�F�����uO-����~l�:庾�Я(b����NF�|Ã���2���MV6&R��֎��*�!���3�_����M���X�Q��"�Hac�u
2 �W��}����9]/��&" W��Y~��B+0�󅝹u�G�]��$>�;�m�m���:�U]�~6b�]pٷ�b'Jt=�Ž�n�AZla�ѣ!"��_�a`/��*.ٿ��8$��2'��>���+{Rjzh���3��p��=�*�k�D��H�^-=f��09IJ�*�2�.��	ۓ����"@��2�`5��|�z#Fϩ;͑v�Ll�y��U8��U����Af�%A�k�5�x�� ���?��"�����q��5M�?�^v2�z'1A��Q�)(&J,���K�F&��2�}>�2�A�zx�^���^0�46t��&��:n��֐��bU,��I1J���ԓ����Z�#��]�
��K��E�Wf����v:����m{���1�u��*:�G�S!��pF��Le��i��7o���<�w�)��T�����o�wI�'y�LJ?��*��@T�01�Ug����L�ם� �H"�8�Z��Y�U!���09ɮ�����M���X��
�:���^[�c�.3Z/���5�*Iމ0�zn��N� ��a<�Hxm���&�6+�}r���D-y:Ӝ�]�z��M� �2��|;�����d;eM%�01&�)��ꊪ��;:)M@~3���Ȗ�!j̷�q�1��mg�հ+h�5�T��iq ׿�n��W��4���i�b������ĉ=��C�Z:BL��H�]4����k��" ��
�E�l_�0�H���Q��H&�8�R����cX"� �0Ѱ^ף�w����(�f�TI�$X ��ӕ92Ӑ��N�2�&� ���?Ռ�1���8�Y�_ͶQ��E�8�W��m4Z��ȍMy��~-��'.��6mi��>�z
��٥
w<�����U�!�<��p~(7�	�����?,L�^�p��:�`R���)��*�{לh�.�Yi,_]�}nK ��M=x��I��vo��wY�Ӂ]B �Y��2�B�!��b�:�/b��)��CI����n�{�$E=�NH���S�����X�W}d%�M��b�0u���������ċI�"~5�a�������H/\�u��S�^Kv;߯qz�yf���;U�r�=�ȰP��
᠈Z��0�<C����0� F>���4|/L��r}���v� ������wǞ����('��Z5��x<�Mz�H�zv`J����xR�K7d�sE�c	�#.�\�E��c���ವ"pD:ނ��E'|�o3��\���\�(�%a���`��k�<�	U��o[�}�	��
,{���[���́���Z!��/i'��w	��t�g����뵨�c�"P�����އ�z�v��qN�D8�4A�CH���w�=���]x��Qx�L-G��S��9�X��s��4aΚ�0��9x��C��m?l<P~�8D���gѓ��3!���I��~[�8U�}��KZ�m��+���c��w|4q#k�����މݢG��e;颬�&����s�T���ao� S�	�:2��&��*�T;����:_(�O�M�m��b�׷+s���M뉄�r>���@D�i2�v�J�����K��n���:{��H��Χ�d{yK��c�2_ ~�)�����;��X�:8Q�
'�k�����_+wD��t�d_$���<!���8R����ܺ�����T�A4?{�h˱���}/���Ǆ�Z#��4�M�X�(J�5^(t�s@��k���sS��r��O��f��%�~�!�Z��m`
Sg)?x�?������/M��gB~r��ѻ.A����z4�q���{�!��.lM邋�
_�`����Kzށ�qif�9!z��Q�w| ���Gv~~"�+	���k5,F` .V�#v�vjg�ߔ$Ϲ�������4��SO_�4lބн烃��/ZMX�B�Cx����S!�i�N����&�e��7�)�Z�]���.�"Q�|'A.�lUdR���F�J(��7����Y�Ro!��n�b�}���Z �H �f����,-*�[A�f����q���R�F�i�Rh7�s(���$շ�?X	�+��"�v����ikk�|�7AC@i��;y�-�?J�$b*=�x�*~��gÏ��F�5N�B�B��i�S�R��mo�z4�#n��.�귝Ƒ����|X�DD���~��&�MB��N3��Ve[6�42	�;V�����e�M��
�9�ȡ�bF3�n�� *Q0���+��L�^%D��R�j:	o|��ME�����mOy@�2���Ew���s�}�3%3�_z�c���P�	b�P�OT����N�E�>J�g����0�SX ��[���1E0�(	i޾��,�Q�˅0[
w�%�@�*����k�f19k/fo�XT m����m.�}M9�r �����7 ;�~Kl	��Y�]��m��e>�f������%ɛu_�RUY�P�.J�'Iz3�资i�b�\"*���^�璗m�g�!I��_Q�U3���yBwT,*MC�q�gSjl.��D���a���{ط�?A�D�yTNMņ:h/y}<4�V�<����l�]�9�H��B&噊�T�A�Z-,srؒ��d�����l���@ʈIpo�*����z���
 �A�D���
�*n��߻n2�<~�8⾅b���(�<�K�~7@B��IW�$�u���IĨ @`i�vz�����B6��R&$j��7�t=1�l�ĭ�G�uW!�_^�&�?s1�&��2�@y������rV/��"dɿ��-!�@��K�lHr�9����KR^�԰`L{��o��J��o��<��O�~�L66�a�qu�\ڗ��G���`9���8m_W�.;���������tɗ〛�����t�L��0��_��չ3c�K��vYZ}K�F׀j���r�X��_�ߦl����" �����J19��R_����)���?< �����z��m����PH�)��ޗ��	�Ϣ��f�~P<�D�C6�~t}���/�9�>�b 0'��������Ux����o�z?�e];��|n;��{̀H1�~�}?	AC�� �l�?x8�
�w�4d4S�r+�������:���&�	��5�R�V0&]�0ʥ��ШH�-��:+ܨ�3�rܪ`�5�c�l�Z�5����ܮ~TD[��F0;��^<�f:�����΅���42�[��s5"R�)�؇~G�˺%�5̀�����12��G�u
:��W������`	K��e�#R_қ����.'��Bte��O{�*}��&5{�.gɃ��mr�s��Kk��	n �}����-I�!G�8���63���^�s����C\zoߓ�iv����n��5���2�N�K�ۑ��x`�d�͹!Mh$�����^e���vP�蜐2� �������tIH���
vm�*ϔ7�/h��3r�S�/�00J3��ӿ�������C��,[\�G4�����ۿ��VK�N�%wԠ#�⠯�ו7	����#4��uy�Y'<j��J��l�,��u|zI]K!�1�3]F�h΄n�����V{/ƒ��q�d.�[%Hљ��#̨��:���|/%��_c[���t�lg� � V����Z�%d8D��j�5T�ݢ��w���Y\����u̸�t���"=v�9�\��^~�ƠY������D�j�R����d�C�~s�PM�sq�=��S��[�J�_�{5�+ުx�9�(����T�����i�/�E��X�"��c����5�e�#��1fW����Xް�|�Q.��0S�=(�h�ǹ�� �`Wpv�w"K�=�Ĉԫ0)���	E�3ݦ*�p����F���*��D/��лC�i�u�$�9Ob�����p�bN̶m�[��P[���?�|?�~�:kp������~�k�?�U�<<M􈋪�5{�]1~�	do��׵�`x����5���v���U��h��w0��m����u�p��b	��5�f|愅H���5=�x�v���*<!�]G⟘�8������T|�؅���� 
[�2
�2ok ����]Y8|�����q��z�rjʖ�d�U���6Ņ�h�B˹i�%�x��[0!���^���Utl%,~%މ��k��<�k�d��-�\3"*�����挚:�[�)]Pe%=�p�3�n�H~W��S�|�U r#1����݂�g��c�9��x\E��IlM���.��K��ѳh:~��X�܇GV2���T�ʭ �(�j7�m�^Ɛ�B�kKw]������aݍ[�A[��9��]Q4��˜f^Fx����gS=�]w�l��"��d���wm��VS��jF��$v:�OrZ6:�Vg0��Uߋo7*\�����,k�����16�RM/��K�$դ�w )#�����Lx����Bd�`Д���p���:�<���4*��$����F6�-�#��]���P}�i��F��54è�T�<�����:R4�����uy�1K䂾pQ���S�_��u��R�E�Am��N���{(ڈ?�8d�VK8Ң	��{�u�s��eߟ8�I�?���i2���UdD�\����j�
�D�?u�辣����6�v�Y`m3�����=y���E��-�M�'*h9�zm�߷�L'?<6f}i_hm`�G���Q�]O����B���8�#��#k���y
�/6p(���%q.��Ip!���ġ$�Τl'�+�E�-ws�ޘ2�d�ق]�i}��ъĈ��Q�;�`��Ǽ�໮�����=�i�:j�N\�i����ٜ4�p���0��m�$6�+�F�Ŋ5�������I"��� ���Y3K<�續�`]��TM��ٞ����&�Z:��9b5b��PeCvo��KgJd8�`A�P��;-���q+�	]��Z����ɯ���ݸȿ��XĘ��AW�e�����,��vn"!]���f�،�~�l$`���*���Bk�o�?a��9q�l|^I>��./&a'���zTY�.wH����p��@v�)dR�?����ω^q&g��L�CK��(�,>�+�������$!H�{��MP@�so\}f��/��6���S�]v X�hQڗ�ʡ���)oS=�P�P�5���f
X3,���㴉(�Z��{��w!ml����,��?^L��_��En�9"I�rX�HV� �AO2o��)g����ȴE�M���Z�Uk^�z�|���<x=��gm�?x�f�B��C�Ƈ�B���a^��~�oާ�E��!����'l0(�/�f�=��5�s=�������\��L0�rNZ�oa�x(��alV�Lq6cޏ]�����&� 2B�l��ߜ�l��H�=Y��p9?\���7�(šљ-�����s�2K���2��t%SU�V0��a8r���aL�bk�o*��j`ˋg��-/�K�#�&]����.
<h�@W�PUd�w���o�,��o�˓��n�?���1�ۃ�^B��i{%�b�m�9@�����E؋^�ˌ�Kj���~XO���>[v��������\L2�>���Z��d�$�@U �vb
=27Ԧ#RO��u0 m�^"_0��of�3�?�rG�UJ�bs��RXT]P���W�Ac���9_�.N���x���/҅�Or���ƴ�?���}٠�,��#F�NY��'�4�`s��L2}b�y��|����^��mx���D�rn�Ėn�O�##u���B��qëc��8�B�����7��L��)�0΁#E���̝��(ᮏ$}�,TF��{E��5���?CY��}4���+�ԓJ:e���#CbD~���11���
�R$a<�b^�g0�b ��|�B���\Ejg1	�J�P�5��GR:M뺫]�}!ׯv�(n�ͨ���R��Grv���r}9.td?歈�\6Ն�UC!K����$�7�*�5�}�kOR��0Q�U�b�h5A{��hj���	�~c����%D�a�@Z?8�����F��^��ms�.���^������\�%ޚ�1������E�!C��{-aA����:�\��Ik�Vn���Vy*X���瓗��]w��m�?'}��O�Lr��:ө:^w]�z�lЯ	<ܖ��>*����z5/�/w���פY�]�b?GA�Q��Q7qf[��D9/#���t��A��KI��mv3їQh�=�Y�(�Vf*ö6>��z�"�p-��Vw2~C�����)N�6�52>��*���}�d�^ߞo�E�aj���ߪ$���\-�K��ܘ'��;��m�����z���[ـ��p,�V!��������}�I����տ;�]#�����e��2��et��ȩLEκ[PeҜ�K&�h4S��d�a�Ѱ�l����o�B�{$����ਇ���(4��FLs?��m�V��U���u�^ر�#c�PO`4�� �9����ưM���Y3���L	��k$��V�A'�n��]�,�d���/S����%�Ί�D�*<%���,�S�_Z�[��ʡylk���k����I�,��FB�)�N�i�Pu���Xv�lv�mr�L��IS�Uu��0(Fu��h�[1�h�Ee�����kH��nn�{��aP���S���W����
.HH��~�KOd2��A?ߔ��bl�O|�D5�mB6�} ��dn&��m��@� ���=U���b�Sf��h��N㔢�I�����R9�9w���ZQ婟n[`��.���7�Z�"� 3��_�2��w@*�x���&��(27�d���M{~D43���#�=���L6Q�nC�+,:�h�%����N�Ƒ+]�$p/۹���~C����� �n���-��U�ߍ�.3FXp�D��AzL
iV?̝5V#�����d�,�9w�Y�����O�Vdl+�oyX���/����3��n�I�b3�n��~v��G�+Q�^'����2Si�>�ُk!e'�txu���w:p��MaX/8p�&�:N�f���-tZ(�f@q�z1L�3��lpEm���_��T��+�f_^
�	B��s��37˰��WLQ��xvJ v��d��!�j@�R���O��88a��t�+�Z}4~B9�*B��p��=�<�^�����x�P��1z�$�����Ku�~���T���0�_C����%2����1]fB��;R�.S<Eɞw]���E���Zdr����+���	3�NC_\��P�Ю7m�x	^�0�����)���ı�5�������t����R�V��*1���[��C�vC ���Qp�.,w�*�u��֒���/���嵆�g�ˣe%��LQ��w7�c�Y۟�]�Ej$�N[@��H���޲������D�/������̇e��c��~u��x,]\u}�<)}b۽���Z�A�F?��-����.#?ع���zH�b(eav8�z;XO��~��������z�"�DL��έ�I�-�j�lnة����B�7���[	-��e��m#+�M�%����9��6�ڍ���R���m�ɋ{�t��9�dT�R����lgMP�����dǊ��"����w�k���cDF�q��Y'ۄ�;�Tn��ʅ�����*\Bs�˿O��2��H�R6�>�������;�)��=�vC�=X�݆a��*�t�� P����9[5rI��X=I��S�:GOUl}�6��IE��0��Y���k�Ոz�?|��y�pW�y')�*��j��7��G��a�����?��ͯ��?b�C����LG��Â�PRO�2��NTFJ��Z�"^��p�4Ѫ�?�:�%;xf䠜�	�(�E3�Hk�;C��!�T2u4���V(jAi-~�LX��r��_�����pngz�w��b�9��ѹ���8�)pgt�m��&�I��?���ݦJ��G�J�BIfy/�)�H��|�'�(Ftk)� %���T!E���\~B�
���u:A<��M��!����K�v7�?]�����P;B&��uAUt�Q?���l�牉�v|Q>K�g|y�襚�I
�_��{�&�t
V��_��LD��`�5C�� $�6MIm��� w�vȠ/���r'�%�Xqίj�+o�fi���#���r��!�c�vMW�Y.�}�x^5�5t�Ѿx�F�N#2�NU�+�Z�"R'g��(�����]>z�p���\	�
G��?C������ذmC�D�vuG����[B�5�o��$-���n�Ǧ�G�+��޾�=�c��=���ol�?�iaw��iF�a�6��0�ƙ��7jEH��	*�}'ej�A�r3G?��p
0��:B���]���R*�zu8���1���lS�fV@�FAS�Ċ�D��is\����Vl~�y�C�=#���ZP�2fF��3 ź�Y���!���4B����1��f�ʰ�b�w��0��Z\���+�@�Q1��c�0z/*�쏴�����
�����y��B�8����i!�{�^��zgم�������WUp�ѺU*<�ԑe���]w�9�Dh-~�Ƿy�{�N�]۞
U��%�:���Ae��ψо,t��'��ߜcI� �P,+���r&�'�ϱ�I��	����AJ*�![�3��T9��H�΃���S���dG�C����CK{y��W�&��8i]��Π�������T�� -����߇�77fj!`����D�j��ml؎�],�ꄢ^Y{����a�wW\b����|�;����SRv�.j���G����T!�˯@�<�B��:v/K��G��Z���k�ĠB$:N��jF�l�꼘��@w�`&�Tϫ����b��_
����sF�Ϝ'!<�BQ\@���� ��ޱ�9�c-�5����4�?~�U/NRX(�S�m	Ql��֍��^"��ˤ�ts	�QOR�E
��dN�i~�nFS�a�]
��Q��&7B:�e��ξ��v~�|F�z"P7��0>q
��A���*<o"� �J�+�)���X/EN;�ա��E��8X�������,hҢ)�(dg�&�+:�3�eV�b��H	�n�}���A�8��b3�t#���?`�|�DxcI��>��U�~2��BC	Ze[_�O��Ӏ��էBzu����f���_g�����YM$��x·������{.黭J�,�2��"�lȖ��/��n��D���=�ar�]��@�����
����>����}g�v8��&��uϺ���S��1��#�����e0m��C�U�2��~�g+���rM"hk
@��S��c!���%ױwpH����,ۄ�i�\ҘV���֪t[�@[�������ǀ�8�g��´{�����+�]ߴ��,�h��ߝݎ��Z�k<�0�ê��ψ=*�1��U��Z��c������5��;�1�U"��_���R�a|VMނY��מ��+&���B�*;Kp;�a
�?�Q��7R�+�:���UP)�9��VwD�{˫BO�U�"b���ߙ�����8����?�rb~��D Qd��!}�RCmga|ş]D���8�r�JԻ�+#@�ꦊ1I�e]��cŊx�y���M+K�<��"��7�Ǟ�J<����6����T�=���wBr$B	V��+T0�|�C����'�	-�(/4����
�H��_�zt�=!{�7�Hj@]��!W�ĺ��pdpsT�"������-HA���mK��ԫtP��^��ۤɘ%"�o�1{	Ft��5��uq����{F(x��e_��(�2r��ЖLsE�@�r��*1��}nhG
��t���k�u���Uj�0��D�o��W_�&ac�|Z�tz�i��3I�� ~+�}��-��Io
��?�R���_��ywcj6z��r��%��u0!���.qz��d�*k�_Ŵ�DGN�E���̪V���R���vrc���@{�~'�\r��J"m.:���%oh}��+���jz'��q�i�[5���Σ�F4$Qa�R !�[z�,y���D�O�A�n��E)��� p�Z����YN��d�]�Q`�y�)\��� WӃ$����v�a\ �1�X�(7���s�-���	%o2x}�1f���`�?�ж�O����R5ڼ��R���l�����߀Ou��l��|��b��gUy�^׉RN��޺�`�����������o���qL}Ve/s��:i@�L)Ū�A�xD���]"X�<��i6�1�c�j(�AS&�sq�43��~PB
�������,<>aŇ�ac��"e�{죜����U��c�6bW�������T��L����C5\���K4��0t2�xT�����1TE��R��fI�2����3f�&S:��F-=�F�2�ʙM���Ȱ����cJ�2�.�ػ����d�@�`ZG<�}*g�N츸Df�}�H��j[�����Ɉ�>A�z�/�8�k�.r�O�O��ww�#B��(�	�����t5i��}�~�b�uq���u��I���v�lu��� �W��˪N��l���"��� $�F>�:�N(I�ru�e���3�`l��d):5��Ȑ�5@|�߬�q��9Lԍ@���E#�.eEoA�M����n�b��c�$��)�7zD-& V�u[e���jet,��D��?g	k���E$���E��7��^?ҽ�XW� ����P�kQL9�1ͧ�����s3�-$�� �){J�"e���J~����t�Dj���l�����Z��=7��d>�����K����Z����U�;�[?2|\����.ͬ�*�җۍ��)�J>�|��ah �'Ņ�ب�Qn�thw�]��6�5���2狒/�D�n��f�ʚD+D�q�	��*�4,N=-Ff4��r�DO/��a��Dj�7?��_7 ��R�j��sG$��	���9�C����+C�gԺ){�Ҙ�l���O>��[H�����A�8Q�Kj8ڍ!��H���?�7�bp@��15<���MK5#9�D/k���Rl�Tc�Z��Sْ��MLf ����E��~Ɣ�3AS�9~=���\�7��5R=ڂ�:��ewz�rR|�h�����Qġ��~����b���M��D�������F��v+�ISʀ����o�פ��B��k��z����83\m"�*�Ƴ{3[��J嬚����A�]�{ر��c�¸-��EUǞ����;rG�P�Ëڞwޣ�x�7�ќ��^8G�͆�1SG��M��dWu��#�	�Ѩ��QB�ۿ�Yz�^zx���ɟ�� ��0o�)�^�hŊ���V���V��Ow���9h��o��I����� �>��x����R�DZ���r:��g��%�9�.�tp>�2�:�V�!�^�ְ�Ɣ¶	j���>X	�U�<DF�~ �������<u�%8E~mL\L�?o�*������iID�n��k�Q˺Y��V�X����؃ě�������#��}K�!7z��9�ֆ���ԡKK�((/%�`$��C`t+�6.�q���v�lQ��Ѻ�R!H�]$�9�
m��	�=��a���Bn�<�p�d#���p�:U۩���Nv}mxS�ܕϛl�ۧ���d�c$l���n�^�T��{-��ˈ?��cK:Ш.K:��W��Mjk�N�ص��ȭ I�����M�&g!��c�&B3A���>�d��ܠ�eh6�a�RVF�o��x��$�U)w�Y���9�� ���D~u'N��Ur�Tj�%�g��{�l+�h; y�̕�u����J���3ǻ'g�}?��|��Ί��6�G1�!�1�/ɷ�{�q��Ō�i�oO��7��a�G��V��S�A���=W\'�������#0�"��o��Q��	裬�;���15���Ev���Z+M�s�m��YJ��<"�ޱZt���?>cz(O���-�"�N���Hy5F�3��0%k��(в�����!���B*=�u��J�����>O��l�)�A�✇vSD��]=��j�Sb8���<���i���·N���Uj��h��+�B��lYc�ߡ��e��F	����a�8�,!pZ�Njy|T����gӬ9�.��x��K�緅�	CdkxH�9��d������H��/�#���S}�1���?-X����
ķz=�'�i4A��EQ���^��
2l=�sh�])�e�j����Qf�6��jȚ3��1A�{�Fz��c7�w�E�����"ig��x�C��_l�
߷�O>�7
����}u�̇��ub�:yl�^���ʲ���Cvh��+�6�^Y�4)eq%}��kd���( �E���S*�+MKˑ�P�f���{W[͞�>O���y����tՎ�?�Q�w��QQ��gos?�s=x������7�tJ�ͥ��X���W8��t}p��)�=��8��$Y����s`oY����E�+i��i*)���f+찀L*hB����ٝ>1T@�Ռ���$����\�	g�յ����RסA���/Po�����U24����{���}�d���	�~��+�6~�3�Ly�#ذ���b�sr9��.�β2�T7�����!K�cfʁx��|��s�-<�rT[�MC��4��k�$Oa�	���=q��q�e?�P��f�|� xr��fƅ	�P�V~x8�v��ԇ�M���V�@	�e������P��k���jm��	�iN 2�;���9��� Z)�3a]���	����7-�±�=�?FI�&l�(��O^v5��I�=�5R'X�_��\�٨�P;�U��>�	�<���?��#Ol3�M�5;ܖ	G�A;U��*��C�#��-����ܤݮ>izl��5���$���2�B��8=47@��tȐƐ����6�N����pk�o��.������|�M+z�e2���}$v,���:�-�/G��<9�H��B��bڸ���!i��P��iDb�JГ��ɰ}*�\K�'^�D.�0�i��C�?!_���>��I�K#謅�dK'�M�1�R����+�76vWw�/HgR��H�!��i�*�.*�[�2F?T@yT��/�''H⼞����E�pmg�,��$���2$k1C�o�|�Q�v�D���V\�p6�l���7�@��##�rpGi�i����v?Iy7�b܅c�ΔY�C*�r�W*��3�cy9�4okgE��~hV�?�<�N�؃]"������>SN>ݠ�s�K$$t�����N�z-���6��H@� u�u3��H�����3FI�	�?8~�
�b��Ej4���o��G�0q��E�7Q!�hdNl�;j�y	�ST�}[�>i�V��;P���]$^��͒�F�H��b��V�CUD*>[I��������vUX{k��]��]�c�]� J������[��H��HZ����
�o�?����˩aw81$��@Z�����$���n�ibʟ'�-��D�­�c�����;���S5��{�����O~N��n`߱P�5�]�ͦO^'��T{���,9�8�������
�5$Ժa�=Q�&e��]�'��,�K��}% Hf���.��?�V�+����NT����n�
��q�^����D��k�+'����O�y�1Ko����i���d_ �B���,�/��;�4��@�hA#�{�{�̶�S�&�g`'�<(��Y��� �I|��*�����p� ?�[XM@��� @�c�'b��� .�߃J�yzǨ�xA�^`T�:��jc��/A�>Lli�P+:�ԡ��!�VR�}�h�c��~Avr��l 1s���o���gS����oWpҒ+��Z�T6�e���d�5�"s58�q/3��\e^F��S�'�Ѷ;�A;�jH�<��T�v$D7�&�� �/KkD2U�P�l-@���g����y+�ݷ����b��D<�:dB�Ƹj;���ǉ"��^b�1�9ZS�ld^Po֙����G�A�菁��S����J~�=�I;�=�q�9+�����>t�l�yL9�J���0Rj�����v�9�O^�X`������{��?	�Em6�B���)�l��z@	�s�G_��̙_�M,�2"�0u^Se����.����a��\e��۩���?t��.��1z#p� a�Wk���0hؓ�Pf����+;p��`Xc�2���N��� LD*��� �,�����;������<�²�"
����/�ʲ��g��v����ouD(8�ѯ*��O�T�������Bt&1�Bi�40q�Qg����l�x�*u-��IS��au���g�g��k����m�BbB$�n,���r�j~���]��f"Ab��e��S���=.@�bG�m�B�ly�N\��ÑHc(\T�k��Ve:pdF���Ð���˜a����g�%MNV�����{��{c�,��,f��Vr+U��6�5��]�I��Z���*f�xMO��1���Ғ�ӟ�ե�[��
\ў����?�/���;YWb�]�ʟP� �i0ЛY�Z�����1Ч#�L�Ͼ����-�C�%��1���B4�e;�8Ϣ�h*����\�x �q��m��yL��LV؃T�.[�c�ZLz�ү%줯٩�48�.f��)��C�H����Z;h���)�z�����C�:%����f5�UWC�3"GPY����0�/)6����M=[+��P�,��u�CR������n��S�.0����b$�]q{�S�$�(A��S���[~��A5���{'��E�i����:o:P?~�x�kZ	�v=YII�2:�>�5J�=YM���]HI"^�^������j��H:錡�HM�P�Ѝ���:�	��SY�a1����H���C&��ԟ�gk�?�gCΙ8/�ڪ�]�֛i_����&�5�A�g��>f1������7�6�䤐4���oOWnBΒm�~�:�	I�yn��u6P��Ԧ@�o�_�a#g�� �8;��>�BQnJ�
�h�):q.��[�[i���g!�x�����$��~����H����z�������_nh�O�zg�}�U��ط���q��=z�漈�[����E���Y��8*!�E�'��4;�G�'s��|~��	t�׮���Ԋ��0��}bҰ!����z�]�e�t�0�o�W�ޥ��A��:��kv�	L|g��ț����5J+��:{��	r�i.*҈�w���*O�wM$0�����\s�Z��n+�P]�� ��o|w������ܞ�A������E#'z�%7Ry�]��[i�X�Ke��d�vwK����<�N�EH�m��dP����`c��\"�.��`#�ZHU�
�d�b�_�K�L���œ�����'>>z��O	�YM�?
0��iU9R�'rD��q�e����'��ϲ$�JTT��1ZC�:m� u�����ϔn���;UN��9_xQs��j��L`�1���}9��2fCn��B0�
k,�B�@�;�B(��S�E٘���u��~��ڴ �1;Dy��;�.�)̉�����@�iJ+��ɞ7Aꅎ����Bה��2�&��A�ktz�v�R�����,RhX��z9���/�����J�Ц��ł^v��X��BָW�M(;�|D�ЇM�m�8�H�G��C垦̭i�	��_S���0k���F'Z��3f�YI��į�jC^ms��XH}��u�Y�8��{��Н=9"����+	�FOꬦ���$ז�qxN&��s	�*��F��Ҩ��!V���^
�Dp��Lp��u cC����kU ˜?!Oላ&��*;k{�@��e���|Z"Q�E�]��٭H���71ھ���b�����rҪ�@��h��}��7�Z�+!K��\��N��5A�rD6�������N�[��� ��eX�����{'khL����W�	���>SS
�o���
9I�:s|�{��)��]:�	,f�H1
(�TM����������,�L��7�M���˱k�
����
�f"�!e(]��@bT�Li7�ii '�p`-�Z*��JT �Y���=�%�#A��U�e�ż�"���~%j�����0U�	_FD����B�=�a���N�>s��o��Q��ˋ	|�U�C5��~�a1��H���w�������#���Z���Ԝ,C����ѧ
M��F�&���I<�[_6�W\-GX��w�+_M����Y����Mj�e��-V;��64<��Ľ�`��E�4��O0}9�Ųw�?9{���<:Qx.U�{���bk�qy�Fu^D�ԧg�%�GAR
4X7s�&�±^����B�?p��B�g��A-Q�7/�o�]���²��>>�dˢ�V}�O������Wv�a��/[
@R��,�9{h��pYr����π��{�zè��,����9-��Bs���,���� ��J�N�Xخ�͟���p���ފ�6�vyDդ³���w��a<ʃ�y��c��ؿ�.@����-�H�Ai7妝=�,n/՞q~a����"�W�,�)�8xm�n���: ��1_��k����ƺ�8�&�W�P�B������Pi\��"C�p���?*�O7��-�g귘���R��0���X:�$��o��9�x�۟�6��A
&çâ?���b�")�MTS�g����3� �n����A��� w�q�6��,��v�Nr��nx���D�x<�1Ԩ�Rه��rFs\�U��Ac��ہ�,9'>�<:�+{d/PO'�?���jc5b��m&Z@���
�ԴgK��f@ZV���c= u� y��b��0t��E�`��e����n�����:G���\I6Y�F���T��d�sM-��Dpʯ:�� �dF�$��fM?\�"Rq�=6��r��8؄��:�X�:���@����L,��J�Q<v,?�����'�H�g4�%DO�̳&��c懣8�74A���%���Cυ����X�&�a"T/B�ڟ��-*@�7H��J�k��L���tP�4��֦,�w|N���>p�]w?`n�'"u���`Sw�\y�
�θx)����P6�,����?T�|Ej*}VZt�}���ʰ0t\���6��M{<r�^�$t�WI9�u���\+�����.M�?F��H�*D��m������ʃ��p#^L���Ӈ�����ߖ�~�`�i=
�l]�bܸd��;%+|'�# d���ٌ��7��<M%涷���iaT��~*�}+���G&�#:��2����bs(&��h�ɞ0C��E�R�f�D@�S�/(h�$ �PH@30#�!]��LZ�;��>�"+��oL��h�|��(�&�p��Ÿ`Q>0i9���E�Yt���=�-�܁�2�9�K�f�!�'}�y��+���ϸ����|Ko�d����?���#�S�i�opR}�D�P��`��FFR����P^��i�]z8Q�RV�gԭ#�W��U!�Gߜ�}l؆uȮ�3�A6=;e�v���B3����	@܋Rs��[�F_ɟ�kk���6+���RN �՚��r�&���2%U!���~��S�N���ո3�HZ�@�������(�)X�%�^bAT�-�mӊ5/,7��sZ���,��s�C�F7��������y�0<�����µ{H-�i�? ipL(���@0ٰ�J!kf�%LOT��$��N�� c���'!o���3h�ȹ����r�v[U�.��sq�l$\�\��q�e㲪n�pۚ�=�ոb�$zS�P@���@��+�3�g8�L�SO�§�F�ƺD�ˍ`����ۨ�G	��'�q7���goE����F)Y0�T�V���v,rU}d�d�K��]�tt�M�*:@���-YûkFb}�VXO+��g� ���9��""�+6���}��P|/I�w0Z�d��{r�!
�<s���K�:R����'�f��d�T�~F�m (���&�q(���Y�"�S�~����g1�������x�ӎ������,A��oy9W�5I�c2��{Ŵ:�Ze���p��bV	�~!r"��rR�����A�ʏ����{�	���ր��\U.��D�@�	\Xo��mn��3�O��c���#~ǹ��p!y
�~8���{6Uy��?�ƚbϵzc �o��O$�kQ��ӛW�XLB������5��t5XV'-{��@,>X����7Î�-��+�vecY?'�1*s�����%���	@�B��;��-���`�9_�A���}� 6�����?\x؄50�S9�\B�T�?����
��l\_�`-�P⿫Q�)��R�"ڢ;B%����\ P�ԏqTl�]99^y���d��N���0�î�Cr�e��_��`����X��.�*����� d*�2�IH2t3�Y�d�׼'�0c!KT�s�/�߃��ú�u��F���P�>}?j���+(��K�����{��T�x��doW�qFB!ЩI3L!ƕ�ʒX�������δ����e)Tm�8��-!Cΰ�{�5���=��h O_?X��#c���}����n"�O2��>�]�'>I�\�  ��U|�q��<�R�n:9A���6z�^�8�- �$�W_�O��/A���VϠ�A�+� `[:�ᴁ����\�aJ��4 ⭐=V*�@38��/�͗T��f��a��R�G�)x/;�8���h	�4y��mD�@'�����Lhܯ����ˁt[W� ����»&9_�4ү�;�k�.^H-��%��n���������ȧ�-!Z�+8�����ʵ��ݸ��ay���1�3H��V�.�s�ѷ[�ų[7���D;�p4�@աg�qX&�1�D6����cS]�7���Y��\FE��`�A�q	�__G��\p�Gl_�F� h[����c�'�J�s��SGNlks�Y�Tk�D���*ɮ�էR�цYxy�@!��e�g��Y�?�U��|��1�LR�d�e-I��M��f����y�T���g�7�S<A��L��~T���uJP�%a|70�>-�[d��7�'͏�6R��i�FNa��<��Þ�p�{u�M(�,��n�ܫ�~�i�A�����J���t��g�`rp���g��J.��-�0���5H��$� ��u:��p;FM��{I�y<ܜ�td�JiB��C�`>�RE:Xd�?��3�kΖ��J�U�I�|ke*2��!�T+y����S�8F��g��d����i��s@~(��(ᩙEĵXd��w� e0(C͟��Һ������-�fc~T̒:#5��L\L��q�J�p3m�Z��G#�˂�ytRPW4Uǚ�'z�fgsc����́J�AN�/P�k���9���!�L�#I�s�z�������j/BS;�������==���0�/�� �/�-㼄K��g���d�&�mJ$�O��M$��v������;zϨ�ExY�]�3-*�	�{�_"��}-Y���R���c�\]��>���\�5 ;�c�2�Z��t*�I��#�|An���yM[����B�s�q�;�O*�"h���ϴ�{�i?���&���Z�&L�{7&�*LR�o~������C�1!t�ݮ�-��%�_��9��p�a:u�7c^$X�3��;�-�)����O]�Л�&x�D���� 4滇�3���K?2�k2�����Y'/9!�/�=NE~cC~G�$|&��X�08���/�f	+��pu�&�b����kA�5{N)�U������$�5]�����q�	`vn6�O��(��LZu�C\'V�u(}���Y��o*�L�һ�)R��m7��gm�~J������c'2%�^��������/�Z3��92j�)鈉��%�� �;a�`�S�+2~k��a�}�<�K2�ș�Q�͔~��Z��F_�`���>l�HV^5����5�:���S�\�,~���@{y����H����}T�e.a����� ^=1 �k%�gmC�������aD��/�{,�;ߐ$�m�j7FmX-O!4� P���{����#"�+qE��A߇���M	/���`�G6��hezի�^�Pd��z�#��hW��Y��hŵ�c�i>4���4#^�Ą�q�=@�zE��c:���=����Y��w�����B�K�c�,ʞ'��X����ߵ~\'�s'6����:���E|��p.��(�` Ϊ�t!�QX]������p�I�h|�֞��y B���O�1�9��_�{����� �˚S�kߺ2����Zd��pR��q�,�ܤ��B_����O�UEg��6+As�%��]� �s�l|������O|)-h�>3���?�0v�ֵj�v��r��V �؎�9l���8$�7�N4�� u�z6�����P*!3=�V������*C�_�m�⿲>b�Ր#�c���9���.�>���zp¦뎲���x�{�\Gܐ'<2����FT����n��I�����*�����:���7~L��4=23j��@Jf �"N�Rf��L�a���-#�f�~���`Y̜�>�\���<�R�QJ�f�b�ۺ��g�-����D E�`�2��������\N:M�J��8(r?�=x�M�i-I������V!�얒5�6��O-qyC�_�Sw:�M\�x�N��0������6�aB�7E���G�#�8�	��$���Zo��PoG�YJ̘.�fG0��`˦m����H�ޅ�c�'������S�Y�3f��\���XJ�:�w A폄��{(x*rf����g���H�-�OC���b�ظ�����
G!�gI�	�@Hd���1���N���{�c�6�A��Vs*�S��h�}��M?�Po�Y�� ��Ɲle=�[�uHb�b����o���:�NH�ł	7rX^����B���CܰVV�D\o��-u��p���ԭH��?#h&�j�@k�dj�Pǀ�� ü��^�#�0����g:Kr�#^?��=�����l��mB�X�m$�qZ�-�ٞ1mU�%W��E�c��ρ�+[ʖQ����feڑ~����a��#�O��
�T��aѧK� m����@����Ξ;���;]X��щ�cT�r؈9�QEb���9Q��_�7e����;�-zEFρH��Td�V��0]HE�ϡ�� u�^.��7Y�#� /V�*L����6t��=���7v!����#�r!�ffB{,�q����?I��>*I�Ob�=u�q�R}WM�K󜶗i;v���/?��ﳟ��;�}�ͩ��V�$񹧶��z�#˽�a:�P����h�����rL�BIW�@eצ\���A޳��f�X��S�\m�����n��̡1�TV?!��Bs�0��/d�7��`��s�t�,�&9-���6��X ާ���eˊ!��:��?a�n�Q8J���BXS��ɍCFE� R ��f�
��pe�:��&�S���I"O��t�yx���; �S��R:2��0�k<CF	:���VON��7�� �I�rOs>��e	 ��ˢ]Pz(
!�	�2�b���&�4�Gܓ�Wka*L	��^Wm�.?�mW`:�Rb�ڢ��D��^gQ�H���
�z9��<�I{�J����n��+����{/����{���33B���X�m`pIv�^�%�ނH��_��zՐ/���*�%����TJ�=F�K��nG+�ӭU�w�?ܐ��ާ��F������A`�@H��Fc��;ݗ���7��%q*�+~�l�<������q��ѐ���i�Gxa���{H%�e��%v��=e �n�ܤ�[�5�
�W̑�[��=���f�c嚉�2�J</�L
݋W����:� �p?�����f����f��K ���gn�X���Z�?��V�H5��(R�<6�a��F�������tQ{���k�_.���N�*No��`ߑ)�!������>|_��{�5�[��^f��kO��[x�RA���.!��e ��V��:��۹��͉ծ���+}}��nٷ�p>\qr�! ��k.HZ}�#4T���g�n&����JE}��Խ:�dB��Y���]w�� {	��,�[�ζa�X���a�Ww��K�Zkn�_�j�N7��U��.{��K��`��,�}�~XfJ5=.��Mۆ��Br���mX�3}�(x=�O��6�J��$B��ɿ|=�.'w���� 4���%ެn�@�D�P'A�Ȃ}�r���pe'��"Y�9��-]tUի���		<�'�7�3{��I��d}r������.[�� �px3�p�����,���R�����T��P�y���Ql��?�I�:LE����۷E�[�
:��{��U�3�HE�O̾G�<�Aq����ƔB��Yu���I�b1`�;��Г�m��j|�L�$X��8����Kk��e���a-e;1�Џ/°ÿ���2$�Uބ�����P�.0�����n�V���_3Ȏ��&�[��ĥ�n9Q�'9|dPck��8�-�5�:��,?2�u+�R������5�L�?U�W��P(eÁ�W�G�bXK�gŔU����?%?�4���|���'���`�B��_����}�m<�6��o��f}�;8���L.��Ma=D9h�	؛��B��<E���	=4�@�c?�uy���T��)¶|rQ�ܨ0D��`6_�#��ag�<<{�#"nܙѨzn]"�HXc��g�R^�i���JQ �"��h�Kb�>]Ez�H3lBv�D�t3����gY[��OX�l�����j�vx������'�Y���:�I��R}��j�F��>F�d�u�GX���1��c�� �3���*�2��$��h�O�������,�'��1���S��֥Eg�ϊ�,����s�oarqh�#bU_����Z�XM+��ZB$?e���RX���~Lנՠd����� P�l#gpj7u� )�/6-h�a�m4�Ԑ�ǒ��_L:`pťT��|��w7+��9*ieC�;��c�}~/���+���DZ��g�Yc�D��X�����{�,L�-�i�т*�>��\��̪��f���.��ջQxC^�Bm��w��Ƣ��w'"c;F1@O�@�f�����9�$������@�n�C�^*�oj(��B���؇<�Q5X���eb<<*=y����vG��{�$�^K���D�Od����;T*�O��J���m��<C�u�Š1ԥ"���;���s+�����RlK�nخ�g���)��z]9��w�$ܣ�A�������7f�z�V��J༡Z�h�'�r��p C��Ŝa�� �Tm���(�|�dl'�@r7��Rz�o�U�ڗ4˼�*�-c��K�M����,�ߍ�v"�8�؄�]����!N�X��Y���E��^������.�x)�ZmZ��}*�6`L6�L�#�x��E����r������T,�0�9��z�X#|���@��So�ϓ�O='k,"�/�S������d�٧@�X�4Uf�8�E�m���<��5Pi����)�r��x��@,���t^�:��i>
�[ȗr�^kŮ�1�����1�9?�>�,�}��jo�\�x�l!9�����@�!�%���fw~��}�}1����n��u��4> �8��Y�6�Aߤ7;�����;�o�>,~L�Ν�Ϝp��Z����xtƛ&MLu佩JJ������1n�	Q�jh1�<
�g��� ��*���������y���9D��	<mt�;y�?��.��Y��v�^�%6h=��^ q32ˏ&w����+�{�k0��-:��!�=߈^�\z?�G��F��hAltd�0Nt�>�@$ޮ/)��v"X�O�$?��tCM��w����Lo�W���h��uY#h��ǝlB(�
Y�N��	+c:�XY��T��6����e�6ժ��6T9#x/�.䋰�f��t#�2ۼ�0�͓����Z�5��/�z�T(	" �"H�3V��e�q���d�%���������Ѭ�}> &=������{$�r���<�2���y�`̦1~�h��e�M�Eb<Z+?���g[���y׉�\��\�x��@�Q�>�
����<_O�`�-����YC�����>��p���eF���xO{F��1G�.��;'�Łe���.��׹|%����"�����Y�����
t�|��4��̡`;ה-t���Q�٨H=*'ߔ�p�S��UAJ{Ȓ�&?��1~�@�4���x�u��a�E�L������Lmj��"\׸�
H�`Wѫ ���tng��v�u+�&�x�U�_����Ιq�KG�|Mn�L�Gt�e���nO^���v/���W�O�!���� �Q����W��N��վB�����IQ'v�Mѫ� �o��}=��Mg{[Io8��˴��o���u_<o�Teo8��-����oV�j��7F�/�'_3gkw#����>laYc�ɩ���l���̼(�����*�nR�#�anm������C�g�"�h�OA�F'�;/���P'6o�-d�eݥX�5��
^�d��L�[iP��ZoZA��Ŏ[��$U^ҋ��9�=�w�Bo����iS��V�V��Pm�S��*���e_z����?��'ꮛ����/1!f2�x��i$�s��4I$�4���<�R.��h�=�n6�/,��%���%� ���0Mו˙~��������ٚ~���� �+��h�ɋ:�呕<���4�bA@��I��j���a������ԁ~#N�^��[z����o�%��R�ئ�T��=c0�-)i�!����[��!&	�%T#G}�����(����(i坻Yb�>��R%�����i�5�)� �]�`�LWkY�t"��4��2m�*J���N�!��TI�������Ѡ���ԦF9ϸ���K&Iӣ�gyٚ���m��PyK���9�)Xh'>RDJT.*����!L!J��[0��<O%R����2;M�N0�Jvv�嵟[��k(�����S�g�\O���y�d�L�׿2���o��B�E��J�N
w�[ �x ;5�����A78�8�s�w�	&/���*2��?2��P��`�u��F���ڣ�I���u2�J��'��v^"�d���1�E�B�6ݯ���Dȹ�y���ںp���� �N�~ޙXN#�#(�N�S�y�u�vy��D�2Q���j�Xt�|I�S�D,X$ze����d�a�T_ޮR�7 !�HWt󓁢�A#��x�;�F�9���dƞ�F
�_x=5wщ�I�� J�t�*�_� �Z6�L ����t�/?�3d�rk�������^>g���{�
Ź����c�[0?���=��T�Z:���i�0�{\=���,�,�o?�`e�����l:]�=��I'�����q\��u�U�aұ+y}6�X�����*��+�m}����>�-
��Cl�-'M��nXp8_��̰r����`��вډ@��Z��Z���F�z����C ���l�fK%���Ҷ<[��|܉�.�0G��l`�4:p�$�H��YFc矱�\�ӌP�e�
v�h=�e������3觤o�|��u�I�w� ~��	��䰼�Y��Ǧx��� �i�K������N*Ά*��������u��7��w�e	�@� �s�y��bg��↭E5��ဣ�ߓ�̃r��*�S���_tQ�'����)��e��u��P
�p� ����(�y����6B
�^���}9���x�2rO��l�i7d���ܹ�a�Q=ēw~�jL�h? �r1�/U����&�+�q3�T���4�Te�ou���ŏ���˨:�+֤�� P�"���ꗜQН(1��Im�jv���Hb��ӄl^X]���V��O("ۤ��;���ې+�E�iLz�,�������}�-	6��3��؏k:���H��o�|o7�<�ҳ�A�������ߧ�Lĳ�)�4�;���9�S�={,�C��-������}�AJ�d�0eݥ�&��z�	֛Ξ��z��2D#1(r�Mb���US�ͥ66�Bz��M����<��ցJ���}��^�;�c������.f��dZ������I?�sMET�v�HTH�<�z�^�����v�e�W���87y;���n�;d�h �q�A��)fzXz�MyA��/�_��$���W�U�ҝ���Uʇ��&��Td@��2����'�R)`
*J�?s+������V9��-�Ggz�y;ྚr;rɷš^�u���HN7m�m�/ �7�Tc7��R~â�ߴ�w�# �޲&�	�3R�{(!��$��"X \�����}�1 ���PO�+�S+a!&~��->d8���^�8��eXN1[u�ͧ��vt�~/b�r5�$&A9	����J���Q�R�j�Ft����9�r�ND]o0"S�]f�K�<�[ryc��7c�{3�(�Jp�̺@2��/ʊ6F��HB�@y���K��d�}=�ӓ�Y�'����F~��&�O�ֺFu�j�~�U��x>k�⌀yS ��~�C���C~;�n�V��̣�Ռ �?��G�,�Ubt|xZ���vR,`b��(F6��-�f�FlЦ����Jc](�>����<UA )��~��Ny7�)q'�<�6Ԏ>��6�S��
ޑO/�;~�w�
bĮ_,�j��*��A-��;,���ז�r-���w�%da+�Y�k]�߷�)���J((qWi�߇K���5�s\wh�����u`�IO�?�����S=6k���NG-����}:\����زwH�?��Y{ہ/T��K��Ep����Ǧ�P��5�t�j%
�e����(I��V���R9��xk�<��������/��7.����eA�=E�Z�K��a-���#�e�`�������!L���N����d0�����D�D@L�[C��{�XZdEW��EU?�lNh|�O��DSy��F�@|̳��T<�<7!N�!� `�d�]�Dt��'"F}��hhW�}7��r���]���9�8Žc�!�j��TZD��(DH�X!�o80_�o�}&fG5�� ��5��g2����ey��C�����%Lt���rx,O��	N��{�@"�]�ǐ��!��u3NR�=�����]��~'���.|�t��R�t�����E�2�`l�C���V�eS؊S�N��0bO�a��� ��][��X_?ԋ�u�,.#�{o�r�O6��I�	�����MZ�m+��
<ɋ-�1�k(np��x1�T�j����[oD�B�8�c��N�!#�������Ѡ�ph�1��m\C��t�9z���o��#��Oo�p�	�j��'���օ�#��-�#�]�2�� ����7p�}�N1V��1��D@�Њ�Eto辦i��"bؿ�5``��Y�d���Z�$1nQ���27�t��0�ؚJd��,]�j����
��;��F�̯��=�n���p�5��8n̻Õ��b�W�\�*��!��Q�$���l(�<!�0<�fY��y"{SI6N6_�����e+\��~j�����"T����Ej��s�`���"�;V��91$���Х؀5�&$I��e�aQ�8�E7�w�,L���rD.Q��Hdj�VӺ� ���d^��Ȯ{�!�V(�z��8�v�R�/��ْ[9zpSHZ<�c�ܥ�u�8`�d��v�q�G�*.!z��3_�<�s(Ǹ/� n�x�'qc"Z:r�Ѻ��t���68,n�f"�����q��U5$(W6����y #����|N�}���j�7X��d ��� V,4��Q�z���?�>�g7�ز�� )o��}K�����ơ)�*�81!݄���F_���v��ذ�e%[�h��\�y��GHĲ{`�{S0����*��zH����Wy��S�ML��2p����Ū�;���m(���/�	&
�\���eBd��Ҽ��/^y�e]!1�Z~l<�y�Ԫ�L%��L4�n��c(��P2�A+����2K�� |\�BHȐ��ٛ8v��
NGJ�wUV�OІW��3h]�[Ȅ��xκ}��3
r�_�6B�1%��Q4�+np��ت�H;�EX9m�[D��6��^���
H�'cOz��v��f��e��=�XC�v�r96~��{����[�|�QvF ��� tXѢ�����0~�A�I�*q`"�WeB�T��2�%�L�% ��/��_3-��V����Z�f˺�`;?C��=p�=���\�8,|��}����҂:7�#���Zek |C�;�Q�F�՚�X�H}�{�'��J+G�PJ%����H�����WE	s�4Q*��䔮������I1��1i�W��M�<฻��r�)c�t��g&paSA�˳u���޴��C��ǫB��~ȩ�f)u'-Sk����y:_ý��tUHŚ��W���koβ!�E�z. �� ���]��9m<�ő�)�iě�ʖh,�09��pzQߊ�;M���t��S���?]f,�,Q���v��� ��dS7,�qs�{�;}����Fn�I���ߨ�J���UU�~A^�Q����+�Y!���0�� ����@hOK?e-*u�J�d��2C$H�,���T4w:'��׆jN�Z�հ*χJ�M��e=�m� �ݝ�}�����l-b�H`�����h����!U��g�B��W ���z=��P��5��ϲ�^*�O�<��2���>#��q��b�XCK�ݍW�Ͱ�<Wf{Ђ��+�O�9y�)u���5~�����n����c��T�]�8����0�ulѢ��`��ؖ�==�K�4���9R<0N�Z��e�.��� �2/a�+�]~��7*�+̶r���dgmރ>�н����ڗ���p_h��ρ����)I��:u��9����ACйpo@���m�ou���n�i㺌*-�ge'�@�K>���9,�"�Z� �������1���e}�*J&�e²���L��l�fG(~���D=0�u�'������4���d��h!�ے���+���C�ha�0esxì�o��κ'�,����mڧ��iZ����m������0`�@�ٔ�ׅ�E��;b���LO&\^h{�9����]a�
taѾ�Mz�͛~��?�u�O�J��R�J:Sj��~�B�)MJi�H��.L�n|liS�%%�T��4>�#ژM��^Z�P^��A�2'MS:P)��+�B�o=�5V{���rׄw��*-U�=~�Ա�@7OǷ�>��bB��6����4gt����J QR��IJM{�]�e��9	��I ���܀��$��4S(!���a����p��8�̶�P��+(���i�&7,w���<��Ԛ�I
��FC�i��_OWR�1�ˌU٠�O��݆~��(��kr}gc�=U��̙��R�<�N\�0J-�K��9�u[��Zٮ�-s���&�_��ikd���Ϊð�;���f�Nm��?�;e��?�5��t�YG.?|	�d.��L�R�a/��ڦ��,QN��9�PZ�Ml�;��~��,�tO�>]+\L�A2Y�,%G���8i����V���4a�[[T2� �s��fԲBr�J�J�Dʞ;��ɬ���p�Y�-%%��e�];�EP�S��% �7�a�gqO�0�%E[v�?�f����-&l\��kמ�@9q��y���%?M�;mn��P(���k��t����9�0[�i�Ia�x$2�1��Y>�jB�a�vn������m�V,�p�?4�A!guXllR�L���S\��Ѥ�7�&�d���n�<�]�
qW��i%ٞ3�&ԘL6�_0�f�"<'���.��S�v!��sv]GRͳjz��j�[$�#T�G4�*�y~��F]�Ѓ���G�9�[��e��|��OF��Pbq@FW��<*��ӿ`�/ԭ\r3��k3Ĉ�&��GY4�J�����D�ʒV���?��ˋRb��ɪkdV)	�+�!.z;�^���<�1ai�B�}�;\mR�O�b$�J�p���|�nU�*J��},�ս,�vq^�!D�JC�\��͑�:���l�u��w�-�%��7b~̒ó�!��a��,���t�פ�S�̆�#1�.��jDd��¢��>+��mQ6n����V���dx߅DδOe6h�[�Ā�~q�"�Jύİ]�Ҭr{M�
��9-B+���(<nR�t^��]�Q�Q�3������̔7!A�Y�κ��W�n;� �q��{���q�.�1�hxܰ�������X��z����CW�)h�X̚��I�Y8�]�;�YP��j�#��,7c�΀���Y�K�^2�Ck9Ɗg�*^��Y�*D�� orO��4΅wbGg�p V`�ol��Bs�Dz���X��P\&��A��A;��WoOܲ#Ź���i���ƢfZT5ɓ���l����O7�wa9}���K����ƋP%�6��O��*Ufţ����UJs��g:u�mG�"E�s���V��m�6����~�
R#����]�۱P��se(yfk)�Zx��)�-�N�Ʌ|�A��Ǭd)��6����ΨP��L��מ��M>a�ӥsb���M��OL9��moP��Lu���������"Cx�!Y%q���m�eE�-�*�~�ar^s��_#~��m]Ay������I��ט�2k���0�k�����gQH��|�����Έ���-��W�K|o,���H�����N ��&Bj��Q�y�'!i���i��H����K.�I�uI�sEB�#����o0]P�u����o�zh��ú9��
�M"ʰ�����2�I�&��-�fss��IL����`:ɨ_\���>a�y�2w�������	v
	���>x�G\V�����#���;�nX	�[(��i��گٓ����53�K]�U�=8	~:��%=�c�}��� ��y�l^��s��dI,�wT��R�02,��T��TS�sl*) e�h�O�I��81	VW��)+0>P��$�k��O#:��=)e�杉�*�|���M���7}���/�t�"j�������|��ɻn�-mv��"����jI�
_�c�c�!>��Pc��ItW����.��ΆE,?����`7����ƀ`K�5؛-�"�5��HYW5бܳ?��(�dZ��� ���OE�UĤ��p3�"�0���81�T"�����Z�5�ze�aG�[8�]��5qS	�+�wW��t���h�dwX�2�S�s{��\l���yqbPDo��a���n��8���Qyxq6�KK�o�:����+'>kޅ���}�_������e�rK������eda��x����#~4ߺJX�HʸP��)��Ā�0�HQhA� ���CN}�f�����:4Ӏ>��m�5�)���X��U��e���#ۓe�8e��BTq�;�Z!��~o��	P���5i`���`��Ei�*��T�D�F*95F^�
_(�;��8�f�DW��l�tg^ܙ�s2d����5�_�ue����D��!��gf��o��dT�d��N���U���a�=��Un�`vۤ�A4֯͛?w�*�4�#
w��b�Ldf��8H�uS�PԱ��9���ئKg�薴MQF����vK^i�� ��	%��i��$F*�D*����� �?N�ǋ���C9��.�Z�	TxMQ�S�uL���cF�
�R�щXn����?�����#�F)Y��	0�r9���V�����.=���=N�@��	�)��~IV���(#"6�A�!k��j��q;H�hp[���dm���HM�;01�p��t��|�+T����(k��n����?��>jD�B1ٝ���gwC�&���F�(��m䘀E��vRa�Ϟ�C%z�5D�Jʛ�
�@�]~�Y`s~R�*�]���	�{+@���N��?h��9!��h0�vC��F��r���Y6M��6.�G~Q�/�d#�O��I�C���K]�R)����="��Y�>�V���W��G.�"1��]IF�j�Vn�� ��a��OgUS�O��>��+d��#dB�K�M���P�`�m�7�t���s��"�j�r�y'Oc3�)��N��m��������'�^ɣ���߷
��0��%^��|헊��H�L2�4I�J��-���2���li��<Q+�Ԇ�b	����
yR�',U��ģ�w5Aj���z}#l�c\J��NZ	��j��^0�.��d�1]L�IZ��z*bygt��� ���z�ٜ����|Ջ?s��vG&4�>=�Q��?��9���O��v[E��#��X� ܦ���{A到h�"� �w��4^@X
��b"���P����G��|�U����Et��ar�V��ƴ�ۉ�Q ?�h��xٓ/K��c�x5^�_�i
�mw�̀��B��	r}���!�����Mݻڪ�����$���t�
�?О�y:�ۛ'}#Q����UW�s���]qc(�I^ӣ�=,��RH��18��%��N����1�ҷUx�"�1 u>I����o��6O�Č+�������E}�5t�?��,_os��5�����뱞7Q��,Tu2y��7��{2�ѡ�^/_T��1h�j���uι�{���EJ��������o�V.�T�L����S'��c�͋�)wi�!��#$�G��Żew�A�v���͒�@Z�r<~ �ډ��6~>�)�Ԣ�M#�,���B�H�g������*i�K��ha{��gT+گN���Mt��.�ť���ŖκS�K�(�n��#���lt�T��%.�7�Z�
��HC�	��-�<%SYs�qKs�:�'��,��4�y�����x�+���c�o
P�٦u0a<�'�A��l W��Q@7�p���Js���y%�7p���0ez�߷^���G7�\������� �-l�g��~ݫrk�`�d���PؾYɍբ�A.��*n����w`�>��N׽U���N;U40#ӥ��p���-O�4�r�n�p�	�$�"a.�{;��EU
����>Ɩ�:
�17��*�O�o}��s�=qJ��{S�a�M!2C�sn�-�86l����>z=WtF8A�g��@��8}�Tf]{)�<-�F�p��	�/2�ͪ��<��+�^A�%�+�H��8�'��[	z��W�q� �]�E�s�F�k���l�[��#.ֶ��[�g�M�8�-\�Й�C:C��C���T�;�@�f�w�&�+߭v&�B����Yy�� ���]D���;�.E���P�FR�C�P`��@���~?e�C�|��zR*d[_�6��\�?h��a����}	{c�ND,1,�
�r�ע�KT�z����o��R����roE����P<#V�_/h8�q����?�A�k�	_�wO"�^�e��??͂��#�%ܣ� �7�.�[�&jr�es�� �sv���f��?ۤ��-BD�uaQ����Ӕ��r^�I�3��է���FV����zX	'�0�+�|��:J����.�p��̍�����%��]���lk
������/�Һ��"0XUaN�Ӽ�-ML�����K�_�B#��n�����<`��"jqյ� M��U���i`i磊>d .�i�1��:��qbϵ���f���J+��W	��3eN7�ʰ��M�N�y���51o쬸���-��g����������:?�HH+`y�����r�ێI2��=?�5�nK�n[B,~Ԅ\��'�&�R$�5��Ȕw��P@(�K�Ҙ���� �ɤF�g8����ʝBk	�*�͝y�����J.Q/3�x�`�2�خ�u��6U��'�v#%3���(�~�|�3�$�qY��/���0c��O+�c�7-�(c�K�W�g�8@[�W�J>�CZ��~.��Q�E��
'��K(�G+uMf�-����o���#������bo���UF)M���
��<%T4̘��S\[�çR����I��6�$��Cs���&�b��'���fB	���X}0��˨jNF&i,_��Q���'�S:U
��u��9o���g5p.�{4M�ふı���,Ð��p#gkv���#�����IDzʅ]���ED�� &@��D���/t�a���I��z7��@��t��Nmᬍf�Pͺ��i�B^�C�>F�R?+�Ud����w�6"����U�+K~Γ:p$�T(-����s�k��:��[g�7Xz_�����f_�+�>k���)"�[�6A���ڀA\�A7��C��?X~��}�
t��,�r�2���X������s��/X���	�{ޢ���0�H4��>���"�cBI��P��~�^z>�l�a�tF�F?���?�2���'�t ��*M���[�wJ�����gh��]#Z�j�@�uf|m�Y���z�`�)��3�	�[�,�V5�b	!A9�v���z�'s>���r�2*��7�W� ��T�isvѩ@>^�>�W�χ�\�@Q�����4#�J0�#�NC�8�[���A8�������r!nc���N)���7I�P_gyʁ,͜6zyϑTR�j�{�}��� H��E�^��38�:��.��V��b��58җ1�sD�Oz�������9�Mq5p,���؛Tp�o!��O�:�����-}����؛/�7:�N�C��'�ɷ�&%o�*\eb�dh�馅�ʐ���-�� �kr#~	�(�l�HlҐ;�L`o�L��8�h�ύ�`_6��5o������%�-I��2�#�|~l��%�/����	����/���%���)��]���Q7v�i��w��io�蛁9�0�J�t��jDD�,eo9�}�Zɂ�Q�Ϻ��0�_���s�}k�Z�9��C-��!F�q���x��_�'�dЏ�)L�-��#����G�=��Z)�����Q�@���[=�v�e;��v!ق#�=��uhe ]�:>�Ccu���a48�!Z��ꦍ񻗁�@G�u���y��]c��]�l5�V��f'h1��T�����d��XgAef
8�ʃv ������;>�MB��t��k�1���ۦ!նwě���r{g����Oѹ�Z3��o�4��r��Q���-H���`S�����݌��{C�Θ0�Q�Ԏ)<
5�� W*��.t����>0\�n�Oe N�����3#���2S%`)bL��t�zb��3�n�aZ��k��.1���aÌՕyzM�,Y�o�+����]Fv�"�{�R�o ������4��o�un�'Ă�|�k['�t-负S�.]��+u��y;Z��e�&��g��w�|�ݦy�Jy�;?�uW�T��,���]��:w��0+FU~C�V��V�4\�%����*Qd,������	p�� b��}ݷf������F��be�8^��t��ZW�KXs���
�Ȗ@��K~������Q����-a���0�g>sM���O��~UG�(bqV/�޻�����Z�cb�7U�:Q4]���?���"(��f�Ei�
o)����(u����P�O�v�7_�O
��i���`-�z���aH�j���	�߹o�3s:P���K��j�(Rb�V���<?[�LO�9*� ������\�d�Ц�c��6����yG,�p's�{[d耳<�h�?�+L�x��UW��MM�:�����oP��ϰ���L/@p���͕.������f�I@��VA+�1D� �z�$ӫpZ �M��E�f}����И���-&��:L�\���7�ݿ?�-]f�����Mj{f�/y�>�f~�֌�a���_H����ͩ,���k�Xk�jP>b��d�T]��{����,�y�C�5�� eL^�z
z�F���2�@?�a�M���g����}��Դ�A[��kns>�׻D��(qo\R(�?f��b��	q�9n���G��kG5�<䴶��!�sHҏ�+-a��zN��HA��(v�$��_'��$P%e�	���d�p,%8�E�V���H^y�c|���8 ��/�i�p��ձ&�a���>K,nOy �3ܣ������W@�>#���@�C�/E���Tf��"<���b�@1W���cP�U�ȏ���ULn�#;3c��_��P%$��E ��=u<�=>͑�j�е�#>Q�!��]W���"�q��Id�좄�n���}��L��9o��d�I������CC���V���Ǘeicn]�*��\���p=n��=�H&S*��H��i�$=M59�=��q|n�Y��ʬѺ��� ��y{���%�����4���'qk�Q�S&�K�!���X�UA���,��D��L����~��S���O��Q�9pe@���Q.~�Ѥ��=׋�#���+��]E�	��W�[��ѨL��	��>��	�h�kqy�4�*��2�DI�giI��w~v%c+��T���љ|�w@��;�l&w�CM��UIKH�\��%��3 0�V��Z��D�990c����������m�����}l�6���H���;h����$E`��s4�Ƚ�Rd\��A�J�b���͝�_JwQ��������h���T�v.�BS�6�L^kv���(D��T��9��9��Rse�B.�P���{�M]��jz�9{�p8N2���tO��Z���KJ��i�Z������v�@���r�03 ��r�O[�Sk��o�޲2�}��.��H��L�v�2g�~!��?��"�Vȟ�"lb���u0�i���v���A��-����NQ��>\,/�+����X�*6C���� ��I�$L�eFOX����	 �Q f�Ϡ�X���2遧.���8~�������q�$�j�dwU��|��G����OMh�Zʭ�'�������s�[�6�W]��PK'ӔՔ_�12��3~C�⹲1D٦����'��V�T��� ��X>�S�N_S� X��j�����n��M������*8�K��i������P(�% ���ƺ�Gc����b3�1�ݵ'��'�G��a&���Q��$(K�Q,�umBU�v6/8-l66��O��5�ْf!�!4�����N�:�\W�E�P��p�+1J�_V�o�\����֜�x�y&Wv�����{����/W����֞d�6)3�� �Wd�h�pmק���j���y�����z�	:�;�o�ٳe���gԃ���[��7�E�QN�k�[]�5E��+�&��:�:�?�[k��V���݆ ��|Ϫ��nbCB�4O�w� L�P��P>�w�1�+o���Er]&p�x��}Lik�5/�a�W!�BL$����
&2+���)N��,���;0��n���t�˺T�[�^*�N��D�٣�?��5��~��Mf<E�w��(�6-Y2��!:fz�9J��dj/��DW/�x�F���C��!���)|���z�B�9�~T���F��8�;X�I����X��E�&���+Դ"^�N}��X�[���$;�M�j��u�-Įz~�h�c�f���#.�|s1q=t�]!��FNө�K�*QK���	�S�8�7���3����=J ɺ��RTxܕ?;O�@A�B��W���"t�`�w*�Bf���V�Ɵ����^����~6������N��d�6ڴ�,�M���i� �Q+6��x�;kfq*?�'5�y�� z�hr�e��'�'%����v�g"ݸ�.a	�,7���T�����焙� ��Z)O����|ZI���Q��C~�|r>6C�shK*#� ���	�I#���c�Z>;�&ۻs�����B��aXR�N<������� �z&k)�Gwoa���ɫ���3UN�
�t8�ֿ�@����1���}�?I;6�%���9��Q���a]4���9-���mB���}M��XL�e*mD���V��5I�����t�Ⱦ��)l�^٣Dc�î�.�g�%,m��c��q#:�+�\�HKuvMI^�m�<���9	�=���� @/�:Q�?	��N'�[���V:���i�vu���H��G�=�������=��XF2p0r�SR�
C�����l2Uን!E)����L��+��M�D��*��XT߱	-H�&�I�3��DP�9�g�؛�B![V=��k�~�3�4 >.�����}qR�ߒ���� �J���/�;��j+���_t4�	�j�	�Ex�V���r��y�0��]!�t��s)��tm�0�ɉd�]�f��+-?���!�۫mQժ��X.fV���ڜi�q�Aj�P��p0�I>�-S�WV���S2��b~���{_VY�	�	�T�I�wer�$�y��s�Dj:S;��)���z#�5�i����F���7Vh4�%A���S`��h%X���e3'Zt�=-�@�5IQ1����$ќ~���5It�׮[צ�ۥ�X& |��\3y��_����e�UE���^�*�<Y�б���%����x��o
f�"�9W[�J���QB".��ђ華c/�>�\�T��Q4_�F|��[J��1*`�V�Kl٧x�+������ZA��F�ڃ�*�&��3�VQ�����y�
kꠜ��"��Sh������ۉ�:NE]�D]�8�{MP9�;:A�!`�b���G�<{��~�f��PJA�J�OG�#��c���iWpjْ���iƏ,^0�[��]��ޱ1ohh���k�-�3P�'֋w]a�H�}W��oB��RK�@kV5�]��@�kY�v�HX榕L���!�T�5_Ԡ�(�����;r|f,���ʅm��06FR���e�d���˰0Is϶� Q�T��e��K3*��3�:]�oX�g��C2"��>����h�|I��l/K]L/���mF�E&�����Xy?���T��oQ�R�PG�j�K(%�.�L���g�;�4|2��*�0Z�A�Q�|#b����v���_aL�s���#&еT���I��4cy,y�z��r^�%߱�N%�Im���|���4p��!qۤ�fS�m������$��I�|h ��?�]
��|د�;�8�QO[�8�Z
5Zմ��I�#�`���v2��6�J��t7������`�d�Uur�c3��A`��2v����O*�J!�g�ge�a����Vf �n���p�YU����4�I���u�c,�:wU�DV� |��ـ��_��,~��򂒙�êa��l������ڙJ8��_���q��XI�Z'U��;����`�Cf^p�[9�a��j���^�*,d�`TK'��z�0Z��>��xX��oKWj˚6�IGF�q�8�%�u��'�qK�U�by���e<W�>+�Q��IJ�~|���}xW����K����*��#�O֡��c�,���T�1+��d��jFֲv���?�S�[�K9L��)Z�ɺG�`Q����p`(6@��WBTESq����Գ/�4"_�U�Llz���	J:���PT�_;��{m.2�=&(��
�^�;E|x9P�~<�Yy�jء�Ąj�x�Q�J����O�܆�AhG�!:8' ���*4���&� ��\>��A�f�80�p���N3�s�{����"��G+{�V�p��� x�%Z�+R�F�}��7v��ɛQ����}o`ϓܨL�Ѿ�w�6B3i]��/�H�dO�΁����l��B�`���>�%˲C�Aإ��^�W�	Y@���LT��?���Dd�,�Y���nzAS#&[4-�9&�3�2K�vNc:/�����(&��!8�n�B�D�p�@mR��Yr�Q^�ؐ��@��3z�L{��;hl\"�0W�u��;Oz.^�v�����
o��9��pU��k�xCp)�?��	Rv-,mC��X�t�x/�̕��H���؉S/K��F���LҶ�'�T�[|�sc�H��{W��5\3S��@.��\�1"�G
gꃒ�^c�aO!Mot����e�kL#*u�]rT�xz�?�h�E#gMĻLX�[����������jK���߽�� ��͐nD"q�^��0#g��|�H�Ҧ����ް�`V�gv$���Q�!R�!+��u���t�RǬ�ɏo�8!e�;k���9Oh2�^ь������T#ly� �=�4V�Fź�+ܠ/d:
^莌�ˊ�鸼ݞ �Y���>8/[{�k�7��KO�+VK�V�ӵ��_�n��K�:"��ܧ0M�!��u�'�s���W�ї[���V��+`b�%Ϟo.0&�e�4�e��yl��Lq�e��%�~�u�Έ���W��<�xl�H�WMril%����;�Fw'��Nml���)�Rm%ո�&c
�v�I�n+�K1�r������y��!S7��]�b����S%X+Íj����M���Q	�{�,n�hega/E�1U��|a���rCJ 9��Ћ��Qt�0uz�"g66j�ʒjH�؈ب��-�.���q/���Jq��''�>����G-���M��j��8yTTd��GQ5�w�E֮	u� ����U�M+�?4/P�;���,�
��Ae
��:ᡶ�~a��B{)t}�ԗ��q
��h�l)�I���:��!9��I�s�0���$J
�-B�С��f ��&��(������3�"ۓ�:�ۉ�D"(�'5!�9�S8-�`	��w����_7r��P�&%�6�2o9[nNV[��{�R.f����>���ƥ�\�ƹ���@���$;��=���U�����T�&]8F?�}a)q��Ļa�� �"�4:A6!l�:��R�}-�Mn1�ū%�ͻt�_x36j�0�5
���n勒���2)-}�ި�&��U�h��:�߿z�"XV���..�(���<��v �j��T�Mi�sٙg�~����U�q�ܕ�*�Lυ?؝��q�)�f�P1�b����(x�}K$��et��w��
^9�z12o�ň�&(�A�O�i�^�2��8�)e���	�6Zh�X��LS՗g�e�?O��[��-��Th)���<��ٗk'�����|S#���f3K$�4H�P��.ŉt0F~YƤnzʎ�$~~�KٯPۍi7J����z�Z�9y��:�r9���T��-o�b0jQ�8��JH뛄H/��^1O�&�4����A���H��ӳi�e>�8�z�wW�3,�K�4��*�����㊖q¶r�s�mR�`��]2��&Anm������C&ݰ>zD���#L׿�/I�p�n��{y|Y��+���R���*<�'۶ ���L�Եv�Dխ��Q���Xs;�h~���۔�7��!D"b��z����:"��/�pљ��4ޫ��v����3Aɍ�*��J)n`�4x��Uf��F/�z`v_ƨ��ƍ�_R��F�N��{�?�&;%�2p}Fr��y��|cQFu�d޴k7�W���l�؞ij��Ւ 4O*���~z��Sd~0�oB�3���P|2��R���4COa=0�ɟ�|�2�8WJډ�5nZ���"̯�G7=��C2{�x����{Q�?!E���i�0ː���б�j%]���9R���0-ż �\жP�:KM�1����䷓���O'���<�aG� ���R!�X��XK����R���e�bf���w
^�4W���������C9�fkƈHJ�Sl$ݲ[p��������=귷��K��`���3;Q�|�(t_�eDE0t�����������F��Et��V�1 
��`�^�����=H2Q��ae����������I1<*R�E�^.3�<�Dvwdr��!���,&Sՙ�)�ɰU���;ιa�2��G��l��{��v5�5�d������A���a8Z_�7!)���HH!{�Ҝ���*����Fm%��[��?�[,|]4-��@R�����N���_<�k��͎��7!� ��F\��~.�7z�6nC�{)C��H9��3��^����$�RY�v���@�ͬ^��:�f��;_Za_�M����o���Z;�0!2Zr�ȩ*R����%%xT`/s�]��q?S��/��o���э�J�-�g����*%�9��Z��(ii'��p�^K��F��<Q)aϕ<�����/#o�|'����<��l^i�B/�5�o@�	��v����D���T�m�
5�}�8��pO$_;� ".n9@y�8��ٷo�Js!�Z�;���[�$�i����(�O�U,�.eKB�`SH�C���"���"���j\��WX����jw�GL��n��q.��PhҦ[D��)�A�[�[�J���AV}��l��,r) Ϡ/�,s�\n���������!�ϳ�{Vy�}?���%��}��$AHq�gjZ剦�ތ<�T6,$$U+�	-�_-3y:]ؼa>'�1~K��7���S����$}V4k.n�\*@�O�S�e\�^?��\��3�Fr�ľ�������C�{].Ϥ�)����!٩m9'��͐ٲ�
��h��4N�,�n��?�?xS�m��@��N{�,���c@���t��S��N�*�*��\>���5���3F�u�������17�l�>����2
V�]A��A?�??I8�MO���0��8���0�v�"8
��W�]���d޳����(�"d�OuE�'�;BKݭ-^n��w���c�}X���X��d��B��y�K����"0�40!�Bf��b���&/{��L¦�yN��OH����8����I�6�&Og����'���Ve�fшX!^�]�0#�
P�*�!@�Hف����-�(h�_�AL$;dO�|wb}�T�,'t�)"oj H3D˵���H:�q��zۈ�9�;�ٚc"�����_-��h�%I@�}��OF�Fj�׿��� .k�\5�õ9Ůt..�G�b�z�X�.���8o?�t������#�_΀�ը �-#�aW�,����D��:���`AN����=�ܭf�?�r��²�ȅ��?�+|2g��29Y!�{	=����S��=;a���72��D�#���i8�W��i��g�� ���Ap��^e�l������::��
�����
��r�D��������´���#�H�ʾ	�[�Q�J"Ex͗��f7i���-�u �2 0Z��{iC�����(�m��A=��V�D:�FH]ѳ	$f��[p
�45�d�9E��������wR�ӟ�T��&Ø��K�����5vsO�����$�oEƨ���'��Rx��nts�i3o��*�I=�-���Æm!�S��ɛ2��d`�������U-GXv�!�WuY���Xe�21�ؓf��������j�-���զ�f�n�ixku�t6�~�q�;/���TO^��qI��KC8.�G@��$tXI��\�
��׫SmH����o�穜�!��-��[Z�1F/��˙�������t\�2�ꡂ�Ab�VJh����GS��4�ܣk����/�R/ToEe$SG�2��W�$��k����);���U}�����e�N�@u{~�3l����,Ց>���#��X'�ա[�Hz��]h�9\V���fGr�7�e[�����"��x���������]�5�q,,R������#B/�W\8�	�}9*@Z�-s��`�`�ד��q�����	
],��o[�Z�fWe�"+H�b3&��{�����ј �!�
u�pF��k	J��a�����g
�*CU���7�!����nDK��������F���	�~4�UxW����R��ڱ�J|�{J��Ìb��E��}�O��O�ZY2e���M��V�,Z���˷�Z����$o,%#;Oֳ�5,�2���^KfE�aL+i���ɵ}G���=��#��
�l@��)��;��SS�j��&�6u�o�p�<�߶�I�$V�z4�U�CP�1K���o�Ʋ�N`�v�U\pt����
��*a��8O� ��Onj�B��.(��
���RT�)�W� ��o����ػ���TW�c.k��(n=�0�� ����&Y��X�_�G�n��P!���]�^.�Q�'Q�duV����c��N'�B���a�3>�N�����0�@�幽a�0f{
M��R���dqL~OO�^��P�5G��#60�\�*|�zC�Gj�ϳ���Zh�Ka��';���՜BG/��<d��L���-�p���!�E�f��ڼ`�9�a\ueP7o��^��6���1r�?*����§�TCIZ_T�V�{�<���_���dB����T�nk)�����m� 7-zkMt�^P\s]:�ǣ�)L |.cW����>E�S�g��;��ck�{PsQ����D�N�N���*�⣋57u��R�,�Of����β�/�I�\?��h`�2	�d�`&�<����G�ث
��qBa�(��r<�� �+����h�e��L�
�ZlrL `-Ԡ`�E�#����'M-U4��v&�>f-�
��-��6ǢlSA-b���x�fT~�+�qj�S��,���6c�3�� ��&TQ���:v��_	�ꤏ�U�U7���� ��Ҝyz#	ǿZ$Y�a���ݰh&����?	�5��� �#�N��*bD|p%!U��O��\��P�Y�v0�f��}*�O���I.�Cf=^yT���t���)�f�[�v�G�Ⱦ���s>��n��K�C���HLXϵ�m0�P���h��\b�����a4��4�Y6����8�B�����o�Hݜ{gy�9�͆�K�io�H��u;������4LU�d������i������	�<b��`�N�6�!nC�xs�À��0���&s�/��5BR��H��1��}o�`ML��<���ۮV[*�8hu��c�'�m���'T/]��f�
���/�- �r����n�ҁ��/f�~HۭI�:��[^<2�D�^d�vH���-���RںK�CT�^�=��D��c���Q�.\
D�l[�r�^?b=a�AƠrB��V9@����D����J.�f��OA���j��=�,�dN=�YK���'I۵�0��@0��N+��Q��k#�臛YH�j&i\te�ߴ������W�a1d�z�����J��JVR�"��䜰��"m�Hg�_�h
��H�� os`��C\�oNy�5�V�Fح�ϩ�SK������z�]=s�����u�w|hԁM,�^~E޷t�ON�1>�R^��n��v���	L����g\�,*`B��r���rd�x��qS������q_i"����44�d���:y�3m���x��-��T+�"��)Q��^�ۄ��^������C�y��x3��V��ix9�$�O��>c� ��?����7c���e�;f	�Q4�6�N���Pr��ct��Fg�h���B3?����"4�V%s�:\�v��i]E˓#�3��L����Kh���0��!��~"tn��2n���j����:˳A�߱1 (Y��25ًz�J�9��1�1���A�����S����Bt��#9m�Z���*��?�\sΕ���O<����3��pc��8W�[��U�P,`<���1k��XL��Ԫ��`�X	]-KC�֜�g��.Hu��VGc����&0�Y%�Dk;*�4�B���'����8ʊtʏ���;�^����.�*�_(����k&���q�n��߱�O#֥I@�s �d�)ۦB�����#*�Z���pAm����P�&0ǌ�&">8=�vy�K�R$׭,�MO����Ct܂Vj#=��	҅BΖ)C,�[���T�qY	Ʈ� xWM����a̟��aB3��_c%a߯V���dk���b�'%,��0�[���Z]<'ke�|���5QE�+��&r�k�VQX�/�wXd/����=ˏ��k?/i��{�؆'+�,����<$~��x𖫿�� E�zDs2ʋ!�k
z,2�-�M� %�F�N����<*��ݱ���v�F�:'&6�6Э��k����1��;c�#ϏS�ʑ4�<� ^�!Y��,,Nm�>>.~;~����d�!���/�=��&2|�YČ�唄p�ݰe+��|`�L�*������� e�̆��/���]�dsؐV;�+�Y���2\WШ{���6���������h���P��P�˩������ǚ���nx'"7�'�vZ���:�����{�b����/h�><`�胣I��e��f`���w��#@^�i�Hx��B�	�X�3��cl<�x��B���i�"���^���[J?�9$QI:�ҪK�4G����36�(Rv�l��px�:;��:�Z�����=&�|���Ω��d��s������o�����-��L�w��B	#�����ЪċJ��p�����ĩ�4�������7��G<���6J�7�2J��+�����0���g���(zߡ؆Uz(/�҉���x)kOm����*Ԡml"R�!��"K�Q6��ZU{�+O��,�<˄��$���;���s{Y
�tq�j��� �BC&�Ņoi�%/�ܮ,�>�Om)gή>#�t��nD$��>%�h4�0�زO;�˥�^�=nק}?b8 ����:8c~g����S�'��:��0���<K0f��Ľ�}�~��2u3S����;>�����޵I�\��7���vUf�+kZ^�5��������ݫU��T��wN�e.��~K�/�p�Itv��Š�����Ӝ���jS`
�z�{.:�V�Q��U#"�܏IP�j�����g�k�ϻ���� �H:WN�;�Hb�U��A�N��mDK�����^X9����dW�zl/��<�X�[�>�NN�bXr�V���l6��Mt9���h�Vz�ݨ�J���>1����b�{�H��$�'�9���!�+���Y-0K�P��g3�����1�Y�Ru��lٓ��w������򺺶������������i�>-b���ӥ�G�")�N�U���"����^_׉(�?7��9M��2̐�+6o
�+�Jo`DH T�%^b� CVT��iJ�9�s��W	�v�3Ȫځ���S���PQ�,-�w9�����������7��<v��Q����;�K�{�����U��?��Y��ǝ��ح��	��l��U��J@����a���+`pF3.��"�C��B�|Hbm�0�f���q��!*)ph�*뻡�qysD/Xb������w��
/�
�1و��+wٜ�XO�=i�7TjT�V�I�o��|�F��K4|"XjDKb�� :���fc>'�dx ]׷;p�p ���&�'��o�i��� M{����!:���k 5�k�DB�z�l�"-q�e�aO�B0�Kg/��et8��U;�&��X��T��&�rSv�^H�X���������ڟ�f�Ԑ�v��*�偹LR��^H�c��k��M���#UZ��ί�9F���1��$!xuy��3�����(O��J�`�_q園���0:U��*��]{z� iW��/�D��<8U'.��;��:�l���m�v�kqn#�iRp�+A\N��n+竇<��Ra�՝l�)L*�?�-�W�ڶ�C-���]h%�֢�)�����m��3��k;u7�/1p���;��v/n`�!+q��K�n�������sԔ)�+��������U^��a^�����I%�=�ք�V{%k�Ɏ�U�[��ŋ^�Ku���)X�QA����c2��TK�U<f�o7Z1r��x�$���< S�`J����o�Ibc���Z,ʋ,�,M<{��Yj�$T��u1���v��3���g:�X�x���:L�	��5ʖ��I��n���*���7k�\^�g������6�xb��2`T�>�N��BݾRjTX�\�N������NѤh���(R
G}Q��T6qu>�h�����U���~�}�9Ĉ	��� %)�@��"L��Ө���"��|9O���/�Z��ޑj$#�nj=�/R���=�Tf�c�7[��ͦ�wi��ָ�ɸ�t#�a]���f�_�t�*�>|9H�I�<{������s/4!�4�^~5^����V�u�#K�7!�Tyٙ:!�3��gR�B��A*?�z�(�`þ`Vy�2��I�`�:�`
L?�A��=2�@�l��3��:�����Y�b�@�r� IƤ�J/��Ο*n������$O����+ :����)����S��	W~����~��)F ~���9d� hȌ����<H�6����\������<���ɲI�vl+�$�?r��-���G�L�kGM�������ԛXUFf����!7H��o�y U��Ep�������;�Eg�68��g�����_�����!����#���˧�5��r���kӂs�Mw6A�v$�9h!P<���RpB�޴F�6h��ٴO"u�Q%��V��b��y�Li�F~�,tDh��_���Gֽ��(:M����$ܹ1�S�%����:Ɠ꼣��
����:��5O�����I��&{���p���_�IqI������ "W���kl�O��qy��Y���E	7��x;g�59)��~�Z��DJz�iߋ��~�>a^���C��J�R�J��6YC�T�J�d�5d�9{h�H���95����J���F7�?�Pq��-��?H�"�Q'��;��ql�=�i)II){��5���M���� ��VDJ��8�y�t��� <Gd������@�}g繧
�6�$[�?;A��d�L��*�Z��p�~�X��x��_E�h���6���O2�.�Ѕ�A�U�%
~o���g��#��"�x��<�f
��d@|�2�5G�߼���PLۛ|��O<�3eP�ݬ]s+l?ޣŞ,��ώ�a�Nw���6z�{T��Rcm	�
oӚ�1G�lF��,M���Lz�J'����!f��4i�ajҍ}�U�<a��w����8U+m��_��+�����ߓ��2!��+�*ٹkso������ճ�	?����4,�զ�o��:H�ݚX��s^fI�^1˜�&�I��~�[��m9ᲀ�]Pȡ�C}�Bӭ�>1�"xGL���j��Y��D�6�.�';-�d��m��6�rP?��搻�è�b>��sTq�M�i?�k�Y����TPѰv�n�G��fs��_��=ʰXa]�Yu8�^1=z�2e?��#N,f[UML��ȗ���|��A��%'��v�~�NPhG�9���n�;���8z�d��]��]B�&�]�'�L���<���y4��E��4�M8�=��O<.'nCP���t�?��(����C����:@41[�&�"�=m�z�0 2���	�Iq��8��lp[;?�'.��jT��tR�}�vL
zlR���v�����A�Ǖp�,�h�'{���/��lz�&�!!!���3�rR��*��L���v}�Z��O���q�����i���xx�Q._��
:���س��O'�*p���
����g>D�x��m"|�p�&�i)�@#��g*8�:�=��Y�`;�(�;�X��D�к�\)�>�����QA��� �z��
�P�:<�ױ7B�/���jy�/�᳿�Z.�t�.�J�XS�$\M,m�f�Rĕ9 �?�j���FJ��zwՠ���uPU�����H� h��vEx+[��[B��g��>^��n:8�.)L��e�w�w�6��'��*���v[��ؗL
�!��^�g0�^S����e��������Ҩ�F��E"�޼"�:�#=������9��۵����L6�D+�����1.��q�X �q멚%���E
�X�L�<ّ,A��7��U2Kiޛ`J��zG�m�_��j�P�*;�H�r��#y��g�k�y�ƽ��%���nޘ�Lȵ�g�n�n<�e�s�ƈY���m1Ͳ�e����E�����t��p<�l��|$���b�k`�u�	��_�{�E\?�L������Gz=a\��Iw�]ȣQT�P�>Pj��� ��i�3T�p��0x��:V1>�H	�c/�� \�'�ˎ	?*�:9�"��}��8�9�)=)���摡�o%�(%g�Ng�'*��&� �0d��=X��!��Xx�o	�{��#�z�]fDk`�=�X��� �݋�
e�F��Ow��gX3M����xbg�v�pA��;�aτYup�U1��o`p%pEV���NW�z�``A�gd�0_��ԩ��C�{b�D�M���.㶵 O�Q8�O�ӓ܂f�i��J�v�ɒr��?tQ�@�R����6�sL��/�H� Ɩu���7�Ǫ8��Ah��;:e�q��`��{b�����]W��aB�����ƗG���Q<*����݉��5Z�Ꙑ1�'pS������!���
�[�V���)�D4>-2^_���yN�K��Ӆw��Tfm7r#Pki��i�T�|����^�������B��^�L6T�G�S� ��N�܍��5�,�涵l��'QL�:@��6�TՍ�eW.#x������O�������&a(p��闸�v�c��	T�AZ%��4|�����8l�Ze��Y�e�G+��U��@� j��A:^��������d�]�V���1l���Uz?�y=GA[�T�������~��t#����~�n��H3���+�-&�.��+��E�d�F�����+d���a	s/����}6�NEV�*\P�#R�z*���� ���6�x��S�*vĢfnؖ��f/����pD(M���h5e�7F�n��J�r�r��2R�)g���2hw�;��jR���a3_���vǗe4�p�k�L�T���w ���t=�̞�w�f���v
\�w�F�}�բԠV��������i����}I/�8y��Q���`�%�P��|����lp`����!���m}�/1.\�h"�ئM|�`Z�LGݵ���j�2B��%��ω� ̗����|��t�g[�
��A��3�wJ�:�S~7�Q6D+���gi��AB$f%;�o��>.�� `ɺ�P��k�3�k0*�!"�x����W7���{�,rӄ#�
���b钋�t�f��N�H0���Ue�,J��#H'��v��iѶ3����� 5�@HQ�4���콡����&hƾb#*���e�jgi*~�F���<�M�m�p��q,���u��L�7��8z��\#x�	���ڀH�<؎4���ml򸴨8�{;-��W.���(���5r[=h��������5.��9�/�hXD�٥ܘ�KҌ����zE{GTHy?��\�m5���E�A���6�y�_��i�c���������T8�*���� 7t�� f�Y<>xM��:'-d����ͥ�< �����S�`�A
�j�K����������V�B�?</�M�PN}8O?���;t�#�S�����w��URĸ>b���4�������{�:�0.�����:���+�U�v�F�����2�Ⱃ�a��%�r�lq������'UD�Ő���dm�U�@�0�!0+��&�#�v��*�`l�<��ϫ�B��2��+j�ܗ�Ҿ�y�Wu�
�j��zo���Si�Xt��dP0T���5��x;|q��"(�#C��9|J�1멁��vH�?�q���I��H����N��&6���l�i��7;T�x>��0/�����DH�H��R<��'��3T���<�-�����B�D���$��~�^`{��@IwT³�!����J)R^1�K�y�FI*�]��w%��Yp�d	�f�(��$�O>�aE6�b��=��Q��
�����ה{r�w_�:�Mۍ2�X_��� ɨ	6������U�|6�3��,���j�{yE��ҷ�L�Գh�a	-�.�s�a�����ֈbn,|fem��,hV�+�h�"S�5���x~�l-���xS% �[u��Q�8p���Lp�" v	��}f�����y�[�洰��kE?�}�ҏi�oas�2���Mj�/�C�:��Gj�r4���f�����2�fy��0/�r���F�;���#o(E�P��a�}g
����B�7������\�Ol	:��{(_�B;J 6��S�=Gce2T ��h�a��O�fS\���f�K�wD9��u�1�M�ZD�5�TRW5��nJ��0�ha�8є�D��0:�I:���(i�S��K�@�y�x�v�}������]��`�(���o�@��B��6�A��~Ռp3�#�#^�:�����4��p<U�^���A;�/�=���aD4��t��<�J:�8fn�%�a��US�#�!K�s��x��&���`�o������3f��v�CV2p��bT�yW�I��`8����������N�i��)�~W�x����n�� ��ى��{��e$1��Y
�祐��t#%Z2�Z[+?@���/S��Ueژ'	�~�@>��<����j��  -�����?�w����)1u���P�ǣAb�W�@#�qX�f���J�1�$����g(]^#	o��'�F%���e�n�Qɴ�h��)��Wc��F��sw{N�o�R�W��������[�-��ӿF��qM���L�!T�0~�a$����S�:"��m�	NL��,y��8�J	b�*�l�H��nc�5�F��6��]㙨rD��^�v�K �� ��ͧ�t��Έ�O�U��f�E%D"s-X�soGh���ґ�=��3.�7��3�	YțB��!��xP���t-��b�A}���6Y�Ҝ��T�q��p�h�(���B�2*u,
��=����ӑ'�4��я��$�Q׶k�c���L�m�َ6���.)3�*�B�5�>1b}��7�.c6����~ꢯ�)k��nG XV�Nj��\�4ѯ�É�?v�-|ԫ���dyc�n� �T�eXlB*}@�ɗ{��R�����F��P���w���'},�m�x�{*%'����r�����Q�d�d�`��f���$pRD'F���׭{Q���	o��$z,�Ǽ��'"�prp���l�.5N�R�=��J�H�q:��E:AEL�l
�@�h�d�kj~��ߠD�*U�WU�`D2��LO�G�{������R9����qQ�.qB:ns�q�����$�����Q�w��>���:�ȣ�g���)4 x��pMX��I��)��\%���S�KJ��ۓ��ݜ1��z!m$�n����W-1g)�R���2l�X���J�k�\�3��홝L�P����%i���S�H� �yд�R"0�����p���.d��V�iss	��G
f�O����b���h������媗_�%H����W��K�7ΟF'rT��(�"i�9��%�ʵ��:�>�P���τ���N��r!��*F�׎�����i������u��-j�peǨ�.s�����i�<[�� ?0;x�7�7M�#�Bd�2-wun
��PH�q�{�,I+��]��d�c���Wٍ�D��E��D8�bΎ���f@ڏ8�C�0�ɤ����[:�d��>9��oY���G����)ǔ iMㇱk��ŏ�xk�B�t�$!�~f1���b�B����-C�xm"MN���g�a���}���<R���H|��(Q�n����z���%�K��޾4+�,w�A	6w-6����ҕ��K����B���H�/���g����|��@�s��Py����*!OC4w̌cs���O�Ä��ۣ�#a���&�J�O��N������N)0]R�֥���W����D!M��8�Ӊ�{h ��g���lldͧ�ga�.y	�����\n�ӭ�I?Z!��Z`S���2��u��=,� 7��6�zP�Ll*p�����(_��Idy
7p�sk&ޓ����qݨ��w'W!�8�	-tcLf��jty�;-��b6�&l*����$�޻`jTw�o��s������҆v��^��*�������+����&Y�dF�?���(��1��*�\��	i^@�S��8�p�����OD��Q�A�#Nj���:ĉ��4�,���uH�NΨ(���:r�/�4� (�Y����&����Rh�	X��n�.,���a��qn��˫��]���ݲԶ��;ZR�����0X+|(�@y��+���.m� @Y_�-�ɑ���΂�{��9���W�Z�e�d�i7�܊���[�Xj�G�0�̫m�N��w[֞+�̴I!l@R�SO_[�{h�ϴ/�N�Ė$Ms�jJ^7�>���)�ӷD��`l>�q<��7��qT���S�%;��	����!o��q�D�eJ�~^|�Lܱ%m�=Ǵ5]��E��jM����9�_�'���@��Sv>�.,��[�A���t�81vq$gu����+�.�����:��:^Ҥ�Qn���r�߹�/z)���|�V� ����q��t�cZ԰`v��Gn�a�;2?��"@9۶S�<��+~~CZ��� ���)]��{���VUٞ�7�$�Dj�;��Iڟ	QX�}���.��X&~\�#Nz�i��@Lˍ읈q*���`�����`"'�9:�3Pa}�!1�C�D���uot���;�^-R���TC�ɣ� �ݡ+[(��=��3	($9��t!O QQ��Ʋ�fy2�(�~(nc7fL����e�t�o�i��?G�8�M�A�2ߐR�n*�F®�[<��3r wHM&6�Ĥ���(��,L/�C�����u��?ľR �h�@�v�1#4>D�7�
w�ۂ���P�+y�^�ŏ1ae�/�%"���`]�'�D���ٙV��<g6/8v�
W�N��yf�8JG����91j{��$k�����F�l*����-������Z�|�+D��y�(3`��wc�N�ƨgb*f��uX2pZ�S�u�	��\57��_;����O��B�O~����	�E���iܼ7���:Ή�%ESំ<VJ�����k�#�E��b�CČ���Q����$hp����UF�_.�7?ȵT$��HZgT�␓�@#
D[��l��O�̡���.��1X^h�%ZʇB��NVl�D!�2����}��W��u�]T�`nۜ.����G��PA�oM�=;���9!�d�$���Y��(�3��.�A��� 쑙"��o���_	M�a�F92���%��@����/�F��ؠ�n:_�D�#�ޮ�ѕ���a��1��G�����?�K�����������8� �Q^~~����F�f�s�c3����%`���2#nqoQ8��#��]_�$��s������f&�lb�bn ���W-�Ҥ���|?��<�k \r_qe�ޫ�D ��	�	����@"�_֥�_d�	~�������K
t �>1@!����6*�0�_oHٱ�ᴼ��ӗ*�����=��hL�rZ��ZKĊ�:H,�����B��s>S}�:�c+k\�)q��Z�AQz���������"����^�fϘQ�����92;_���>�+GB��"V���%QM�8�=�0�e�f��	!�WK�� �m֫;n�`5�s:��zfC�6/�M;��N�ꋁ6�_#�eIg���SR��Mn���N�������E�)?^�>�ݤfl�p���ɖ����m�0�~%�p�*��3%�Z���M~�9��B��1#wV���{J�>�B�3�P��Au|Ա{�(�T
'�Om��X�_��9�I�HqD�\R�еN/�x�M����FY� ��=D�,%ׯ�Z:/.v���/��<��c����y�\��n^�ㆆg�Q���[�@�����&�E��u�OpG��7�S�me�U�m~���>�A����{S-�ܙ��j=p�U��&ŋ�`|�)�t�4"r�t?Ò�!�s{���Ð[�`O�M�*�t=|dֽ��q`�z��`7���u�q�bW���MJ����oJ�e:���J��M�Vő�~�L�$�"y�h�{W�j
���U��G��H0l����s_��e�>�I���Ju�����Y%��: ^T�-9s�PE:մ!����~�jyg(��s�H�����ͤ����v��� ��sH���'����X!��z���=�01>v��Gj|Gڦ����O���10&Y�%ےf&��@i��,���4���HE��cr��q��B�d��f��	��[U�7�
{�Q�]O�`T�"@�P�ht��Ҍa�������;���Tk�/��~4�l�^?_t��͠X
(7@gnO|�r��R�3�J���c ��0U����[v��(�Dk�a��t�n>���Z-��[b4w~����_�H�Z�f�O��VD�G��tb�ș,���Krn$����gV)�*����>�W�a �CWڪEI`q�;���Yj����kL��s�?�t@���3߃��B*�l[ϼ�'N�l9�;���o�Z���:�_XO@�@+�T@Q`KC���Ai8A=�EHʅ�J�	�eh��#��"��:yxio���p������	\�CL��nA��`��TUsW�L�������F����]D��4	%��_�e^��k�����ͭ�.,"�,�2mH�y��SaMk6W��X��1�[�|�y��ޫ����ePOo<�
]�����i��L �i8���4�.�3!;����9z�Ϳ��縶�b�p~1�l��3���' ߜ?�s,:r�8� ��f�<F�>6��ͷ�'����ϖ�й��F���o���i�op'��� B�@8�="�FQ�������ƹ'(�c;SJ1`�3��׺U<��������0]�[������3�k,9k9 ��G�;Qyc K�Ť(�s WU�dŬ͡��c)"3��{�EA#���=D���|m���C��z�'���ۼ��;��V�EaMY;�H��ear
0Р�JI9�M���԰���?� �� �
����	�W܉r�����#��h�qP�Dd4x�F�R�!���~�-�E��_.[�-V=ztlV�̐�w}xZ	�E+Ϫ�Jf`ISm���ds�T��>��{�1G4}/o�Fz,}i���Az�}-/��BF�r�4�-�6*ǦZ-�pf�I���9=�g1	Ԕq�"7����x�$�)�*����O^��şT,��dz������̘��[�`Jj�p�f�@	x|D�g��fǊ��
�6�doʊx3�A{�6��W��f�e��XE���/����a����CS���|
N_D=hX�+�	mT�	�<L�*1��$�J1�\eE���gi"0-�!�T��խ�|i9҅M	�	Ԥ�L�|)P	ET\�#���`j%�@h|{E�2��6����=U4a##����c�c6o���#�-=�9�rR�H�-��v��[� ��q�YuH�11s;���b�"[��Ŀ��Z`��WL�L��* o2޹��$Vx;��*�b��ko�Ԭ�c� :� N?am<6s����z�J�Q;Kԃ�6FFsZV�J���{r�W���I���!����c�ǹT�n<�as1�����qv�򕰎���[U�r ��}�}��iH���A{�X���E��pl'da��s��j2�xv���{9q ��ٛu�c���d1�Zq5��.ǘMJA�b	�vx(�g�9�$+�l�@z]/���Y��4;�7�%���ږr+����4�إZ��aƥ#%Ew]L���C� �n�/2��.����y��^�-{V$J��sk8�
�}oX�UgBH�R^ȱG��}�7z�����c���]Ӗ�8 �8`PkP$Ų�8�ۘr렐� �Ǹ �{�q���X�Q	ϣcj��-2�8i�=b"�m�uFCq̣��NS��J��e� ��fJQ�]6B+��r�E�A���k/�v}̆NAj���m�-�V��K��R1��x���#ш	������iz^�ɵ�P��j���V܊�w��k����/�,�a]��*��4_���ԇI����֜y�Bq��/wt�6F:�in�j�Β�X�O��I m��"&"?�(�gKP������
�l�Y��aὡ�'�D��ю>O�E!�%3�Jd;��Wg�
��;%H�붨ޛ,�T�D�g'I�� x����Di�c���X�P�*��V1:�9���%l�Mh�?���ӕ�`��ް��Q�󔢣�qRz��v��Q����Q����Eʁ�z��0��"����G���I&Fʓ:���tÌ��,6�M�Ld	��sk��Y���{��m�Y�B9��Ŭ�?e��΀*+#�Ё#} mj��[�r?��hGޏ�?ĵRH��&��ik��
��+Z;��d%&Pu$OZ��7n&��+a����� ��B��()%V�9�xb�tИ�z�$�r�{����j��}��4m��ܴ�j��:.2�&����&������9ړ%����E��RB�hhHͷ,����u�L9/^��$�W���@������Ͷ�S�yC�q�is���H��\VF���&�(I��X�S�M�#%�ѐ(\�-^��G�1W�⚤�)��4L���Fށ�("_�˯q���ޗ*2V�{�35DK��G,�%���iv��l��b;�S/]����>I F�2����!���R-VM#��A�-���z�o�dݿ�l=����Լc-s��~���wo߭$*$�*
]�
T��ՓL(��lA���3xL�'�����`���>��D��-�L}���ǡfC�����.}8�t����fE�@5��xĶ���ޟ�K��L��7;�vK���P[�r~| Yn�5���4�Z=�-����k|;p������c�J�*��u1���q�	Y�d .IQy�iIH�iL1g�R��k�z���*�s�2B67$A�B�qdc��Y�`߼�O�/KF�.�l�������2R��ƥ6�._2���O�شZ�Z���5z�Z���x�����! �A������l}jsNw0�'�����ʙ#�����7�%�Yvz֦=xG��[z]>�B�I��)N��upV�7��=�<���y�)ַlN�����)�(R{���_�]1�K{� �݀K[�D]Ȑ���Ќo�q��'c6ߛ�����D,�&�a��D�X5z�Ѵ/�&���E���W�w�]���GM+�^:��'Y�㥔����$0�N�\r]���S%�G��e��N2���y����g��b��J<����v�����ɋ�`�d�A��n`f-D9w0�=ܶH�G��+�۾��1~��3G/�]EgDF�$��˛�q�yH��0m�r�����ÏW���|���f���	r��gc�c��Ŀ�UK�E������?:�����w��� ����?�р�
�5B4<np�J�а����hF{#�
�L�bfo�)4c�. �j�Ŏ+ĝ-Y�B��K,|�]�HZ��-]ၼ��"���!OW������� J:ޛdO��`B�Р)&���dva��������8��\4
=��zE	Ϙ!L�~��+��Y��6��Ѻ�.�����86gm��=_�:�����0�􀪡w!��e�Z�p/C�D�P��\���6��q�<���2�(�0>)���_�\���\ɤ=8d��*Q�ٖ>�U�	��ޚ�� �s���J�B� E%F��$��A!��mm�r���ޒ�Zf�xI���;t\�Jl[X��U�,5�\�6������[���S�'�P��(?�x���#lAa�ඍ��a|.=�Y��B�cd�pO�"�$7t]���U��Z���bJ͊x[_���E/v�Zσu����1�k[�[��T���E/z���]�LHc�]�:<�N���<�p�&�<r%k�����<J	�ζbVu�x牀ԤX�r@�2.]���~O��E[��;��	:$/�wMI�n@����b��1�<֭w�J;e�v��<E��p5��rw,��a���xl�W�8�J?6���H�c4�L�:q�4���d�(J�G�G�4�s,���(�7�\n�2ͭa���C����c�tFs����2)Jm��/�e����ya� BI�LJnn�3��øKR��"ܮ�[�_'��>�5I^b��X��U:�p~� ��R�!����Ƅ�A�fE`�={O}-�uR����i������l9G����+$�T�d �������kw�G���\/��|�rI��su��l1`^���a_?�kK��#�/B\��e�!r}�kSΜ�'�_���k�*�7���}���� ��g�?1Q.���ѱ�T�8-��أ���O&�P&f��������?�_�Lb.�Gci�t~��q����Č?���=B{�| �wX����I��
[��(�O��[B0ق���ȽE���S=B��
�W�
��P���4)�eq'��vv7���_�d��l�刚�#o��n��~��F���kS6�"j�V���<�����j�ב�R��Mj��x2���Ho�7�J@�q{}ڋ�0�~���/�p�'#��6�@� �8�`!����Sk{���Q��ފ�{�&�1'�b��z�Z��LQ��/޿b}7�x�1�0,�=�5=�BH�J~C%�J3a��E��.�3����c�q����o����Q��AՅ�g���E�s9�
��=�8��U%Z��~��)���4*�i���-5����ƣ�R���Y￪
����m����U�PL�ע������I��'�o�Z�d\�����! Н�<?.�2z�9�i�LtH�R=Ƃ{��T*�Ȁ�$�U�U���ػl��ǝ\�q���ſV��v7p�]6|�9�����M�s	S����r��)d��A�@pu]�,����ic�2���! �9р�:i4�^�P�Mh��\�X�=���oH�����y� �~��q��k�c��X��W�gVd>�<ó��t�w�yd���y��Ag�¨��Po[;��5�&=�]��rٟ�}���[�l�/mؤS�5<�4�!�S�}�i�C�z��������pk٩-�'W�A�v6�T(�WU���%bE:Y�L�P������#Z'�K�WU"7AߔM����XD����Q.���\�dZ�iL�syO_��{�B�^y8ӽի���r'��Ͳ$�rĵ\�%������a[d��NK�9�H=(#uT��1.�S�H�nV]���N�춞��d����<��ͥ��r}&rl~t��l�a��BB`�ޔפO,��xV��M�������q�V��`(���s^`��r�����b�ԧ�Ǒo���� ���?� uK+S���l�D�%�����.S��*��jFRc���s�PS�/�YV����u�˯���A���9��Cj����?��]�_�rE����0n��G��u� MX�r��Z�:#=��Vh��	qt� �������m��H�.�DI�0Fc،�!YQoq(���3'�ڔ/�ݧ��2SA��4u+�71�c�����Ԛ�^̝F�;����r�H�˨�rdG���̙z#��v���,�h*X�|�O�2K�Pn�x�qP%.�z��ڕ��[����Gǚ�Py���m��	����z7A�ce�	=;��C�q���x�Oj)���U\N�3�D��J���mGYZ��^�I ���H>u_"b
Sc?3Y8'������|j�o����SU���ϽB�zH��!�*B�6�`]���51�oX�4=ަ��?9�R�|�S�V4K�$��5SRǧ�P�]���V��6�I��*a�"�ǉZPچ6�>���n��^�^�p��*��^�C���uL�@��`��g�*!�.�P��@���bʳD�I�X���Q �����b-�yڬN�3k�����9i��`�V1c��`ؗ^�D�M)�/=x���OYo���I��h����8��QD5�9����l��ϗ�4��������.�q��*o��3���_\�~�z���X�2���Q���#-�P�#Ǩ��0����~\$&�s������?�f@%.���ގ�t��y���N&��7fu�R�Eh������~�G�GM�(F����x����X�Y����-,/��@Fr�}��K1�\-� �-	��|����D�5�Q�bCe�]����\��Yz���KH]���h�YO�A��n˹#�)�Bl1�pG��@5�3���ź�^�+�URj�+������o~�Ə�˭�"&�u~K�m��9 {-��==A$���"!l1�TY������y:"8�\{�S�r�][__q��I��|�p��:��=�,�Le���i�X��'G� �!�|�<����oD!_�'��s	�wN�Qp=m��Ӿ%�}{,���<��µ�э���uT4�?u�EzDK���R��\�9�'zڴ��5�Q��EKX"�p N�eR����8=2D������Uk�;u�S@1MEKm�o�J�����_Zr&~����L�V�H�<Ӡ��H�CX9'>|]����%�f�'�AF���q���2�{�HE/���P�$h��	��y_3c9I��"�c��y��B�a���i��4�����?!uȟ�����Y-���d�oxGr(-���i�ygA�Ȯ[u�Q��%��{�q���ūr�b��,�Y��J�a9^��ds��6��V�=|SGr�KKQ x*)�Z�,��=�|�QZ�x���m�~�q<�ғ3��`b�H��e����R���KR:<�,Í ��?H)אڐ�3{��$es�CD�FoLmw<�����T;˗�����G�%�]i���3�����$�q��.h��bg'�Ey��jA�����߃��n{ �3�T@ŲǤP��9�m��ň8�Ew���O�&$}Pс�Z�i�G�gx��`��&�Q���v��q����*��u �Bt(��=X6:�1��
�I�.����T���K�TqԴ���"+ͽ�{H�
N�������Eo=..���(�'櫫x��Jm�Bb�����E敲��a�� @i�I
���O�eT��
ԫ�ɽ��E�ǥ$����N�l��Ǩ<%z��*��1�z��_��=6��f`\�ʙ������Ѵ��&���5MŦ�^.4ɕc���`
���Ұ��+y��N��4v��(-���ɻ>��<���TσS����Ѫ0BP/z+e	 �җ�0 ����]��~��.<�ێ�S�(Fvq���pZ���m��&����	S�i� ��Ln�+��[��7�A���+�B��>a��j'd���:�㴸����EAh��5J_ֹa�Z�n#��-7!tJ�FiߙT���y2�ߟ@�#�j�	׉�.'p��*��9�P�(��2��'3ak�;�5���J�$���8�����7�!�J�6�e_��s�9��'��Q�����d.�!3�y��?2�����o�w��:^W�/�UG��rj!�-�F^�J�68�F��_Z��ǟӌ<7�}^� ��Y�wΥ��L�hBU�
�wjs:��
F���{�����WV7D5�rE)fb|=�ʂ&���tc(h�n'�A+}�2u�t���:^V�'���}y�����X����=KF*՝����g���^�k��+��PM��K�?�)24F�e]\6�Y�Qo�,P@��*�$ \�;�F���5�~�XV�b�c �� V���a)�#��y�7���o�?�����Q���&�1���E��y�"-�}�0ü"�NQi�Q	5n8�P����Β"'���&x�G~��p���z+sڂ{��tc>`��aр3�3��x���%��b7~_�Bݝ_{�Լ�>?�ߜb��88����3��k��45�Ŭf�{��x8�6s�%������_dO/ZO3������2S�"꣰N���qȩ9���s�����n��ג�{K|�F&�T�:L����8�q?���z��o�M�X��7s���Y1�F���y�Jbr9��i���EL)�s��;�4��g�iW�_2��,N/��"w~��.g��=���'��F�gYD��r�n�U��}ߨ�^̺e6Ry}��Pn�/�����.�����|���h�}�/�os}0�£V����[�eaF�e�z�FLJ6斸a�s�R��dZ3y���,H�����3tt)�`c��L��D�|�򄋓}{�[�R�e�{~����l��%!kT<:�e��r���>,�-�]���V���?G�f}3��3AQ��Dq�+{��>H�cݐD�#dO��,�$`��|�s���c�u�c���V��ã~WP�t9���r�?�/q���ιڡ���h��Y��J�����S��s8aR�?n� �n'MV��t5I�����ɹ�1�p�V�ň�u�W1u�W��
����k�s�"���h�,O,�1����N�X�����O��
	4��q���˚�Js��xW3���[k��q٠�Ϳa�	�;���a�5��ͮ��w`���Y�4�N�bfG���"@b�A7��\ɯ�Q9��D�We��l��j��@��|L;x����[c-:[��m]r��a��L�E0^�iq��Gⵓ:wT�Ly�O�3��MvN� �h���<�ȸ�i@� ��;�*]�"�HRj�D�q"{�Q9�g�g��ieCU�F�t�({��$�vw��0s)agS�弲:�u��%4���i:�����ɀ4?o���P����t9��'�㯴\��mx1$�Q�i`�P���ee9��U٬	,�aʹ+�¿կʧ��M�)ȸj̓ %�J�0>+v=�å�=䄾GV%�Q{�6d���Ob�(����8V�����d��1Ƌ��[�l�u<1,��5a��mؙ� R�C�,v�yE�CC�I��'R7�X�a���V�K�lWu�Q��5X�:�tҨ2�}f���Ÿf���7���
C�2nz���Vm�	��l-�a{���aB����y7R�K��)�Ǻ�,�?U+T��5��c��Y=\hn���AO�i��\�C�H����-qC�a
�����s*�ej�W+���h0̼�	!m1?�8����p�W�/��ݿ\�1�8L���7w�zF�66:�^������ ��1'�J���pa�b��g��d��T0�,+�򦱨�v�ݴ�;A~ϯ��}9u~#�(]��-6��>�9o����Iӹ����[���� ���]g�=�^�����ϳ�r^*y�b�0 �G+���|T��D��	�m�T)�Z�A�O{���$P��fkՕ��N����ͥ�+��f5cm���FB�@x�鬫�;ґ@�V����4G.�?VҐ���)Ov�}=��^R��WF��}=�������^��w�嵀�b*���p�2�1p�o��.+�#C�0�V�'K�e�3���	K�����ļ�X�&2��� (�v[���;��#e�tS(X�P����ݩ�A�à:'�Ã�IQĠ�R�0]�����Q��
4���r�h�пՔ�q0���<�f�����2إ�%U<@+�P�пg�sPJ��cg7��M��|�)\v�;���t.��C�]y/����<�I���_�)YIJ�Ա�u����{�-����_ޠ������:�-��v{�o�1J��='�?����W^��KWa��:;}�{��[8&W0ǋ�_�t:�o/,0$:�6TKv+�1N���I���ך|����l��&!m��b(��Ɨ*{R �3�1�Zώ^�c�x���#�,�n�{5MB�}:�0/�Ik�*�DuM�)�4��)6"���
��4�ё�t��%L�l�&��G����%�Ӧ����r�{�&�3�ړ����b�\����?T�]�Õ� ՗ eYϏ�'�!�@�8��i��ضs{n�,Я�*���흋u*�W|�r�;�4js�iB�AM��{i��Jlcl�:��d��֓PD��8�O�Q�o�n���+�K�������+�r�H�����pk��1��Xᬾna�� D���>�i�ܢ��"<�b���@�]uW])��ĸ�j�#��薌@υ l|{����9M�����i��OY�%S�UW�%��uL�>�&[������p��n�[,2��i d���杻��'���0�*�Pt�h��dS������u�c>(w���B�r�%���nj�[79�@�a=�"���tZ&���K&9p�f�>�{^Z��������g��$TmJ�mw�����'��֫'�6��;)W��Jq2�dj����1�%d'<�����CjgJUʨ(�kR�|l,94F ��r(�ͩ~�Zi�q��!T̠(���>+���m���Ԁhk�ZzX6�w��Ҫ�7�=�|�,� ��Rf�j�],sr��logdbݸM�Z�	�?
[�O��K���ci��D�"� ���('�J�Ւ\gJM|�<�`�ʔ��[q�9�)0r�o(z�����tmTȿ���ڟb`�S+|�ˢ��n���
r��cv��G����K�f���R_f1�$�b!� Fe�mV����0��d�߹Wk?�e7��lR�?+���⊂��aM\�r}9�����rV)��?����@o�m���2�v�z���=E�B8�86�T+����[Ty
��.�Q<����$Ѝ0Yk)���y%��e�@��U9J_АM��W�?����$��L�Z��z�-�f�ZDL�h�z�$e�w����K��X0\l[��D���Ӄ܏/���
������~YF�ˉ%R0F��kV1�^���> 0�����i��

_@�ZP��<%s]yƌ�T�))�t��QmyOa!殡�v�0-�}ъ�a�R�F���/i	���Z8N�[K��>b!��M�x���&�!�0B8�Lc� z8���j�.i,�A��F+@��h�1���+p!�z49R[��Ce���1�p��J.)8|���#�E�MW�� g��9(nJ�Y^��{�����sr*aӎ�U��T�`��ƭ��)O)�SM�l��=W��;C�0s&�\�c�2��ef�&�6����)~��(?S���*)��s�N�t˛��X�P���N�n�l�VR����	İ�u�؟�ggN��6Z��[R 2�#q���2-����q6�����̓d6aw�R�� �Z�|ݡ���{F$�t�����F���Q���??�@$�L0@�r8Y��`wo�T��mH��b��	ɲ�m���C�Uʮ�VR(g�,G6���b���A��)�V�'I�b�b�E��9޼2�d[cbلd�?�Y�C�W�T]��}6���X �Ba�;�b�LE������7k����3�vh9�\7�V��mȕœ��g�Zd�P��;�0O�d��h����>�`��O�|:�B�_2��0��f9�s���F��%�%���?~��f����@�>(�y�^�`3pm���VHWRTh���2ֹz�5c����RcV<�U�j���F4�Yj��l���CL�����n��-��ŀ����y{�[Zl`..�Y}��x��9M[Bc���s<����|�z��!h���è��Ι��������yh��V�]�Z�!���A�4���G�~e~�%x��yd����XE��Ӱ3���m��gt�d6SB��'i�3'*��FT��5E��;r't��1��s�?��Ex�y3�!}�0y�x��tj��t0j�c��b�ϻ����1s�K�A�ـ��������"A_I�H5KŃA���`#�]�]�VxeƊ�NP\Gg1� Ş�$^���/��t�5,�����ŚAA�+H�I�?�@rbt��_���:e��8zܼ������2{�:�� ���s{=�߱q%%�C�����c�����^ ������44{�����Z�d��S:4�@[k�y@A��K��j@��޹�n�QCfp
�r�Mޚ(���L�"�p�,���Y+��.D�
���g��u�l/
�vT�xz�ؼ�!�p�&_��"Ur��!��K����p[����1����ʾ8�p���!^�Z�� NO�Ք��ML���,���`�Zp��U܌�nx՟��by����JU�|�7�JP����˦tE.�\�9!J;�V��Ǝ3�<o@�c�H�WA0�J_����ɖ�w�ɂL�8�i|�p+
��'@"�l�E�e�a@C�] hl}��cW��M�o�{o�c�Q��y�?���)M&M�M4=w����~���üf�<�F3�X�rUv�����mp&7�\�S��y3��u(�6fi�l��R��U��B��u�����Y��^wjwn3M䘮��3\��-�/�"�ml�\mޅzg��Y��LM�p�}�\PJ�Z"tl50}ƫ >�^r"g�{~u��$�7?�ä$����z5�)����8|������;o��Ie�y�?�����H���gE�64d?T.	~�5yO¾I�
,gE�Moq�\�[gC-O����ړF�{�N�f�f��4*�q�K�`W�];��/ZÓ��0���0�6p�����JgԿ�g�
?��|�q�{��i��A���	:�"`8�kOzw�M����@"��ʹw۠H
o���2��B\L�"~�}lX��V��qvxpQ"��!yX �f�Kx�]��!�%-Q��QO$rΌ�Ӎ���vo���)>� ����0�|?1��{n8I�4� ��nB����$�p��*5=�AG���Ss'�sD�v@.j�Q��o��=ޖ�����ؠ�iJ��!>�کr�-���-U}�����覀�e`��u�f�o�d���S���|�ȡ�i��#5�)�o��� =��y�e$w��Ցǽ�NL:$��!V?�"Ԅ϶�1y�v�,Y��[�)���i��&H�����TP���NL��x�JL^�I5/�<4C.8��?�Z�V%�Ώ�h�f*Y.C���k�٧r�7�8~���Q�^U�#N�eH[�wAV#T0�b�3��7'  >�:�7�{�L��NkJ'�/��`.]�L��T�8"�t��X���8�#DWY�mN�~2��*�1�L�Z�</
�IX��i᳀�d�����햻�1!�$򵩊����1��J�e?>#Az�+	&{�ϻ�Ʋ�t�}��F<Ǫ�6�Z�8ׯ ����x��D�&�xb��ￛ�k��Al��V�:�(�RT~NB�+��<�b�H$�xe��Ȥ7�*$�9<�Ͷ�� �񝗇C28-��"�y�+��^y�
���Ц���&��K =���+b��I]�W��mY,�"_�NlY~d�M��D���N*������ctM�a�=*_�9r�a��(:B����L�DT�@���,����tܠ�+�pܯ��E�SL���?s���0�D����塃-eiw�"Z߾�;�����z-�-���W���\���^�疁ʨ?�Y)��f����A������xg2�I��������|v��;}�Gf3D�ԉvJ�C@�YN�4�<��1;�z}B�l���.2�֡ڶ��'(���\
ӌ/��P%j����ҁ�0���8��A��Su��to���_���M`DL'
�W��P�i��Y=z���xs��:���֌'X��Z�Z:iS�?y{�eU�Xu=��#s˳g�y�{��0Չ�K1m�ùrLo&���'�6����RPb��0�(��e�S��F>��٠3��َN2��w����f���+�g��͎�;T	Z0龹20	+��
p%�/�{sj��	��a�o�����Gn�S��?�AV_�y<ݒ�������)�{gc3��u�.V���&��vc��x.U��`M�l���l/=Y����?P�)�]浕�&Q's�=�yT¤�_d�ߑ������1`h�#�=�Z��
��H�CR�U�O-M�3ء`
�ak�nZ�Ȳ�m���("uC�O�h���.�������w�S�~��!��H�k�{d��C6��:����0w���&&����x|�d��(u*�'"���]�D�&�<y�g�%�CJ8H��v�ҭ�����Uq��8��7���W�>|�-�n`j2���xUf�	~T�1���c�7DkD��7����� �Q��
>I�R��)]M˒�k�����>��_4%{Bb��wt��+�6IV��\B����r1"p��֧��O{X�*f{��Յ5��]n@vaϗ;0[:�6�e�F���l��Q��IK	{2pШxj�ppX3x���{����qi��̽JtK������r��}w��k��9��
C[���<8��!)�x�f~JR�����e��w��ML Q�>�Չv���� l�<%S�aѺzPݶFJ��)1yS}f���E0R��YCmcr�L��Q�<�6~�䈻���i��o*yY/B�0���-�[��uF�:��F�}ˎ��iY��:����I�=2G����!�f	+���@b��e�����n�yɃ8�$�הk_��A�F��PyN��yo燠^���-��p�(o�����&������3-%}�c>/�U���?��Z�{�>��4��� ������˪�d��pY��ZA�Qʅ��A?q5%e�^���y�@mz�_Ne6� �&��jS��:���OW���^�~%��%�,�#��i$�\b���M� ��������l�@���q���"=#5�=$|r�0fɐ�\�,�UX�:����_��ӻ�^m"z��Jx\õ�(������h��t.��e�t�=��իu#?ޝ.�ܐe!1�f��r�ѓ���%ٴ�Gc�@�/m2(�bb<��k/1��<���{}n|�K4�g�s�粀��J��~|؞I��bE������-ҕfc�����wU�i%�y*BC��|~S&��|�5|����U��������>}8���m����&�+z��껷g���La�ՠ�'���f{L -����"v�H�&�l�+@Y����1��y>S�	�b�ٳ�Ћ�|��n͵�j��ï)J-f%��ۼ�[&m�6,IBG�G��.>@��KR5�dI���D-]s��(�.di>��r�9q�a����P�t�~���5�ǧG����TU��f~�|@ ��b�=Fg�;��5{��3�@���^W��n^,V���A�V+�1��e.�,u�eʺ甋C�2ި�c5���-�P���d{\И:
�(\�B�g3t�]�Q�rQ��I��8c���G��:4IŚ�_�	a�P���KI 1�^A��_�#jʲ�i���+S�n��@E@7�Ɓ��7Kg���j>�D4�٫my�ND�mwMc��#7�bW�V��C�G�>����������9�R��8�K}��V?����23u������V�6�v؟R@��a��쇆�y�$��Z~Y�{;� ��f��x� �'��^9"5��m��6n�rjCq��0e��l�@�a�5�+�1P$f�������eK��m��EQ�T.��'�:\�~9jb� ����Ɠ?$�<z������<O�'?\�.��y�3�����c�R��?���%1�l7A��)1�i7`������?ѳ>6��X>�L��0���0��z�J(h�-
��v������ߨ��V�o1�B�x>��
�mk�)����rp��nċ�|��(*>QXV)Qܠy��4����,��p��t��5�>�"ic���$s\�axʟCMh���Q�ϚN0X��K��a��%� �%��k^��_kT�E����f
��_���\zwS�m��[�Ͷ~��N���hw!��1��y�i���{5��RZ��Q��Є9�O�Ih�����t�]E9��%�N����?hlu��<ᤞ0�%)�c�M��'�)�������ʁ ��/E���<)��ثe;d9��=7(���?�(�MR��b�/e:�{���y�m
��!AR=@_���+o�Vރ�X���#�"�*�S��	���OX�6Z��f�#FW��?.h�rҎ��M�ȯz��C ���,x�D6����6����4��P-4���b�*�C^�
�kjl\�DD�%�����aO�z%�A�?��M&���	��t_o�Ŧ����F����r���Ė[�Ӭ e�n�c���fڲ��X_��X.ba�r��e}fbH�r�Spq�	o����D�J|Z�Y
�Vh�l#\?y�)�( �o��u�4�V�C��m1j�2[K)4։�Bn�F�{/�������Q���}�Ǉ}d=���K��!�T]U�8U�&�c^�G:�$a�f�`��U��wb).��+���t��ʮ��hD<tv��*g���Y7���<l�	��L���b�]�;�K�/ճ���z �e5�-��`Pt�����Y���1�/�Ǵ�aR_�-��D�S��|>��iͅJa�m�|I�/O`��U:ظ��)a焤���8`0��$�`�[3����KZ���!�%Ϩ+�9-�� ]�Kʔx�/4�������ur6�{��2~Ne���ʭoT!�6!J�A�`pjl"Ͷܫ�-`�cO<K��_�y�Ee�e���fIV�9�N��z_�DᲐ?�E����qK�I�Ձ�W�T7F� 1�l�?{���^M_���a�Z7�ho�:�|&cT0��)�1\��_B�p4yQ-�6����q� ��'�c�H�V��H�"���
}�O����+�#8t�������vI���#n�z	��40HR17, `cce�ؔ< %�K�Y�Y�kW\�N"�<�"�sUyJ�D�P���PK�QFk����vo!�e8�g��U'�'�m��?�p5Do�K�诹��zT��mJ��φ�!7�-�4k�[Ì�+�EU��z��	�b�HRpI	�I|�j�ےtx�V�4�i�#"���O9���ٓS�wG�'������@�O����Dzi�l{�q���dzkf �T����W�#$U��ǈlC�.T�,�|��3$���@  ���9$��ƥ�Yڣ)ǥ]�O�phY|g`
|���>Um%=��'�h�P���7ë�	~�MGu�Php�)֐F�Q��6�t�Ű��ɝ�h����G2�a�e��SI�PX��hx���9w\j�O�"������Z�Q�|���$y� ���ZY8�ӕ�:� ��Mz�J  X��`J��y����:P,"}Y~�G�>-�c"妲n�'��*̃f���s+̛�4�psOC���$�@��|�GFRn�E��O���^�;!�
�ʺ�"j6�T7N
��;�vzXp�7ͺ�W�����9	�f�/uɰ�!D�/��р�4�G�a9#]��ڭ�Ž,�T��|��=0�o�W��M�KL��qLWv���N�����d�|,�楨:���y�:��V�,�d���S���]�6��˘��^��9(v�7�In���Ip07\ӵ��ܜ}=K���u�C}B\���0Z�p�q���;��q��աZ���6�Z�-��R�y�Z����vڢ�>-��h����U<2/�)"��<�����uK�cG��?6}f�
?�[y����!M�U7����  ��4��t���Y�P��QQ)F��	���K�����e��AI.��ś����wOd��wCk��ӊ���TG���#�6�`\)�#]Ə��M ���)�p�J� ��+Ե��9�2�Dr(2.ӑRX�m�!���#YZ�����f��V�V���%d��<�\���Wu���gNR՜z�{/x���� �����5ð�)�d�ubs2��p���={_��������W�M�s:9e9"vҐ�|�7 �o9�hU���^j�f�S�zj��T��aO �!��v��GZ�?-DfT�Oha�(m�蕧\mcVĪ�� m��3 h֍X����V�Zҕ��x�X��c����|�ˢ����&g��I]���@?��Uj/6�s�L3�@w�=[�`�
aӂ
d�����ю3+�`��ܥ�C�{f�.��죡��?���!z��/B3�mw�iZw�a��u�Wg]�0&	Z���p�E6J#�	���-SSΊ,|)bΆ:*y=~��(�@jr��!�XBj�+U��'�XY����
�`�!�\�\O��T�\:���iQ;�O�n�^-O�H�0��\7�����&p�G~�j���G!B�)��5 !�^s=���*bi��ِp���w�g���>(p��l ��ega/}x�Y�W���Ql��R.ig��N���\�����
A�a����q���;{N�P�cV4�mK����k�����-��R~��Ė�i�����t�c�M�JnX�A|a{9:.��+�0�#��C��S�i+)��#ٌKnO�?/�ˮ�l09r�I�(ԙ����6J���'�2TE(4�'��(� �~�ޥ��kX��F
_�v���kf#�'5��et{D��	L�+8����Е�z 4�k��q�`e'lˈ����^PLS��K�Z�AM'_,{�,����8�5熛AZ��$��h��_k���o���1�)�g�$0���v���A����L3���}v�_}��7��4l�rϭ� ��;Va�Ruѓ){Vĺ<�ب�I�b��}����^� B:7�/k"���g��"���G��*͏@���$[Č`/���#��3:�IS���}�K�v0p��M�ݮ/!��?�03{s"?'�����q,[��Ë�,\>V�^����R��:��jJ�~�8��Ԫo�*/��Z�F�4�Ѣ�q  X��ü���ڱ@��Y�wY�&!�X�q���ؘ���UT ��R��Sh��Dծ~��V�C�hC���↯��bB�p(��u��T.��i�)+,W�UC�b �~�5k?o6�~B���Icl�J�y��@w�o�Q�W�Vk����}-3*������G�7�nHp��Hry��nIg?� ��ё~��jݳ$4�}7#�܍�a�=?���%�.[j"�6g:��a�b(��n�(���!^)�~\��X��?M���_\N�0��"�����s¸��Eq�n�c=�Z���>O��G��K\�Z�E�Dm�ц��$�M�>0���~���8ی�"�IG���&��I�k����I�����:��zr
�p�������x��|-\�hb�Hу	EV_W+ _�b��,A7�6/r���&�H���x��`į2��[�ɚ�-�l�0�i}���V:*B�Q���%�@V(�ċ��r5�r��k���A�H�Qk�}���}eD�ͣ�G�� �
�v�	�7Ꜧ=\)��ø�7���Y;ưn�DՕX��[���� ��I4|�P���v,�?�r�؄�z���(�π�C�Jc���f_p,K�^����4j"Þ�ټ�"��(�Ц�����LZ;�i���h�ugartuPmrAQ<���2�Ky!T��g� 8��Әh}﫞F�1=�����%$7��,�"=�`b
�Om�;�/�ֶ�P�����)�	_F�l��v|t#��
��^&npnB�xX<V� �.0w���7r5OG�D@�e���D�"��;��qw��g5O�J�P3�)o����7���E�����+ؿsH�C+J���,��?���5K�k���U��6�2|��f�G�ddJ)�������UI�J�z�{���:��6^1��D�']�x����I � ��LK��O�ǧ�p��zb(��yɖ�r$:S���0|�Q*�[����|��袢 3ɸ�����d !�!n���g���8DR8�ˌ>Pz��(�tIqu���|E1�4��l�	>����0	��PQ���+8��1}�	r���ۍ@>�3��;�{#����z�!Q}*�b;$��Oi��;i����ɣc�K<�9�Z��;(����1�0L����z6^��1�$���]���%���g��x�M�����^��5ٓ�·5�c��s�lI���0l�oK��H��v�?�,Bg��G�a��!P����%K��:��b�_�w�9�/��,�$�%�}B:Vĵ���z�-/��c��S�M��,-j��?��9:^
6=W�����F �.#��r�Ԝ�M����oG�!�D��lvQ?�͔�������mr9�^����L��5^��4����t1lR.��^QL.��FGHR��B\_�/B����Y��)�B�����CY��C�v,�^?�s�p_Zt�{�M[A�@'x07��M��Q�x�]k�d��6��rD>}ie���z������=�."o�N��S�0}�w���4�y�2#�D[�L1|Fwŕ]kac�pO"�sʤ�2H�d��e!��\l������ض��P�����M)�=�
@&���0= m��	ZM��$כ_����5 ��VP�wɀ��U�iV�]�h��S��h��Y�I$\sF�e	0��`Y���d��</�AӋ��������u�xi�<b����8���+�*wtT�9�Q^�9<Ys��$G��׼<(�~��{�[��zB����{�ׁUeA�l`5�R��bkS؈�=h�W�%�Q�Y �1t7	� kO�,'fn9��Y��*�EM���&�����R1��˳@7Tq\�bG��d>�8�dr��`�q�ט����+���p.�~ڂ���Ȣܒ��WNLд_8ZPB�3���cŢ?�w-䙮k�%���rnhR��&�������՝�Z2$��#+Ba7rD���;�*T,g�������A�2�L��[����D �4�=��@�"�6�s]�xύ$?�� s�?ө~����p�P�.�Ȣ�%�S!��p	[���P�hb�ߎ����|�)%��#��097�I����O��b��1΄[�AmN8��ga�I,��>���~nh@kfi�F$��p�����c�'��|�YE��λ~`�����Ty������C�ɃN�K@դIN	eP� �z_Ă:��o��3Y;�qr�B[�����D�8�GV�%	�6��s�a��l�r�|�l���*Pr�� ���K��Lľ[��=�D�:�?�?�������'՗����]b��Ԑ|TO|�V�l��M����l��Hm�����tE��	��ؗ.k'|�u`�^(9�H.@�-Q�?%��d���
of$�}Ѥ�5z4�D�h]�������ǹ;�U�ci;�ʾ�xz}�jv2��k�r�@�j���2���ύ�"�C��`�&�o���0t���+w�t��=`ھW���FBe�BҒ3s���ge�Ir0�~
�nӥAc
���@���>�(Gc�� F%��l��ŗgS�ے�������#^���[�	S������.q����S�S�Gm�>�%w���-[�[����3��'��!Sa�T��%F#��������>k�VC�wE1�+q��d����9��_�f��Kry^>X�
�Y�"���i��[��:�K�ۡ�!�4����	�԰�v2�>|R4���8�c�[q��9�Jh�1��~�^Fw����0E%P۪���f�IA���H@$��7j�b �]{vǛA�`^Yt����D1+cA�3�01a��B@�qB�,$�~N����#��H�z�d��+�M�NQ�2klȦ4�E��lʿ0d�����gX/�k,��B&c&����6ٕ��̊e&�]X���^�l�m�M�tJHV@:���F�!uD�1���O���fm�Yy��_$
8����f�$�|�E�/*,^t���G��o�IC��H�B�s���[�*�kC�N������f|�S�.߃1�D�T#,%���'�>�����~q��hW��ҫ���'�6�Gp����9wx@��w:L?��?˦{�\u�����k�p'��g_TX�m���*~��{�[<�#���H3͗j;�Wqfj�o#�9�J�Qɋ����l���/���+�ʖ6�&�{Y��o-	��I�.C����xP.!C�5� �������ܝ�'Ã��?����<(����ٰX*c.��c6lh]������e�����l�+������
���4J�����o'a�Zg����m�C+�v�hV�KCp�GBY��m��R��~�z�y�^e��h��
�u��;����T����a���3g�0d��n��Μ��!b,���H���<	pp7E=H�s[崹��蠦츚��=!�Ȍr�&e��z;.���F��-d�6�[�h����i^T���{�0[}!Q1�Mr��m�-����3�j�|���k1���Va�HG�2���z��kf���3�R�7���o6W�~�=`�&��[�5�s�A�D���5�|EN	пb3����AuP'��?ub�gm��l�1{qUx�_	^DJ%�j�2G�:%����H���g�JmS�[�o�I�aDc8*�X<�U��+tu9N�����
ϼ!mU�sbO�3�X�a�����[�����P��!Y����e�b�	�Q��̡Z��j�Wǔ�Ϣ6��4���@kξ�t���N׽��|z��H�?��u�w�>�Џ�b�ޝ��U�����ܨ�QXD�5r���V�9�J�	cҎ�w����P��a��C����K�� ����s�[!sP�Z�K#����`�Ct��?!J�aD�7�Z�x�����0M��T�9��2�rS>�ǗŕGl�}D�1�/��q������u��J���3��z�-($��=��@�`�?8Q����N�Љ\�����^�b�/'��Z��u��r��LՈ��l *W��M�d��g��Ζ`�E��"��M��e
>-'�(Y�U}�u��,�y��e^(��̔s�8 ��*���0cgm g]��>�+/��Tc�cH�es�_���+�^hT��� $,�4B���`�~�_�����R�E<e��W�o�9�H�	��������ަ����0*5��ҁљqlJt��1�0��M�e:�z�sC�Њ�6��꒿�	(HbC�������JEC�BLcO0�J�38Ԇ'dT2���� ��2��y?Tơ��y�c8O>��x�-<�B��v�y8�D�!��bY�Wi�s�W�l�4-v��wxz�֓����0�Sx�Zj�~8A�/J#��r�ݺ%�0�s�0�5�u���x�yt�&Fm���~��D�Xc���F+|�{�9��2W�kH.�?7�Ҿ�"?B�����
Q?�QF(����j�Ϙzjč �a�>@zZ�1�
�b�l�)���'�����M�7p�p2�S,��ӊ+��Q���2J�/��m���)2�>�0<l��L��}3g���vl�������k,��z�Hj�ԛ���֥$���p2���䲯�Zb��RaO�_�0��B��t�N{��KP
z������MnN_��4����F���L�t��ZF]⊠�'ql�'0m[̠�vk�h�4���/e��� ��{��D-�!���`�a젿�8�I|-��ʚ"����P�0�����«����9 4:l��&H��D���Sq"�Z�Xu����Ç��j�F�ӁR.c�Z!��\�%���vI�B����1��Q�q���S�� $K�!(G�ty���0�u��}�Í�����#)� s��x[Ms/�M�ߧ��WC��z-A��(�������������|/�\�֊ �!֪Z������6�y_Vz��(�F�耒��ှ w?j��b�w�:����\b��)aL�ƕ!�_?��������N�����D�q
j�����)|�T,l��(@�Զ����L����}d8/�-)�ku�4QIvb0��኏�"j��T��8B���^�-٫��AsT�a�(ښ�{�$\Bg=���Kx��Â��X%�?ʕ�.�5�Q��Ӕ��!	jzd�vs�T�fq����ZX�~�2p�U0H���+�y*�#
>�O����D�Q�A�s�B�r��`[S������N�q�>�}5+wt}��#RMq���.��zG%Ѫ<J��iƝ&XO!6Gtm���#�Z�|��Q7|-��Z0�[ �����^���Ϥ��`�7}��}(�����. �O�X@+~�Y��HW@nÆ��L\s�zd�C�de�O��}6K�JD�+��*�� ��y
{�e��x�\K��w]
Y:<�Z`�!r�}厂��hP&R`]x�B`��V�mO#���67�]�g�~rؼ�X�̛՜� �A0�i��-,��6�-��{U5<Z&X�Y��A��������O�RɭF�˥i�U�/���^�G�!c8j��]-wsv���ҵ�-a)u��I�������y�WA=���UU*�$	in���A�H?C�"���F�JoM���/O� [�&�#^���Wms��� 1��,����%�Ԕ�|;T7����s��+rk�,��n�+P3{���^�u��q��\�7P��ju֫�OƗÀ��ސ��h��c��<lQ�����>#-�Q)}��h^��
dR��۔粒P��(߾��\@(���HV�-Q�KD>��K�]�N[V��:`�!��N|��m\�=���nȏN(s^�����F�t-�Ў�e��P�����5֠�8���j�4Z�*�'c���a��m�) G�0Bӗ*�p�����xI��d�og4A���s���?j.�gq���F�@?/�����n����	�Y��hD��:/!��;/{��ӛN�:ŕ*�=�/]?ў�'g_:w��&{v�o(��O������.j����v����n<@�2��ű�s�����%Fi���%��o�E��j<\�rQ?�NE�A`�>��	U��B+�O<�l�/�щ���]O���ȸ+�gƨ��XOQWےm�W�Vi~�~��,�Mٱ�q�sp�Cҩw��۟�k�l��a5��A�k��T�7<��K����N�q���UwV~Q��I�L?�؈�qT�;C�&k���Kr���0K�Ĳ���m� �0x�%�ށ����_���� ���撤�,�޺����9D�pE�s���a�	�[? �}�/(A������pq�Kc�y+̋aP��{W�Ӗ�v�j��� ��/_IH����F��s3%��w�����B汈O ����GS��pL~R4A�.򓃶;;P�2�3����� �O����!��5�1�T3m��"}��O�1�<�A凱�w/��:e�iG�����'Τ)r*B_�<X�ݲ��Z�'݀w�X��7#�=8�����B���gh|���*ʒs�Cm3e��Ё4&��'JsN2�A=�p]����ˍ%�-��l�\��4�\����3- ��QL㑮�K�\�;�pL��M-� ,j��F�Jid:�4c
;�CY��j�˱\k��[���
���Z����&M��tkg��i��Z�n<�0�6s���ۏ���7dt��aO,^�q&�ʰZ�P�Q�G���ॡv2a`j��;�w�m}ՑNGl+����y�X�}\� ��Om��>�W5�o�������r�Ĺ�[�:'x���!�	do�ĵc/����g��;�n����6�e�?�X��V�Cy7�S`PÀx,�J��盉K5�-0IF�,Ё�Ȏ
��7�t�Y�NkW
��q��p��3����u]�,6f�3e�-B^�y���c7{<k�����Q-Y���&a� �|nI'��a����+�%n�Q��(���������h��oqql,��;.�*K��JA?�[{�5t[$@ug���n��,ێ7�l[�2�-���>J��R����*�~x�t�z�X�&�UԿ�Y���Lu�)yUko� ���3��s*.m�v}|L�U`�8c�=��M�	�>z�j&�ܶ���������W"�#����2W��9��KR��`��d/e���v��LTv���j�8	:����@DO��D�{�3є$��VK�����˯6�_��oqo:��h��h�1�8L�/��,~8^	�݌�Pƾ�A�H����[:�+=��ͦ�`T�9�����Q��J��ߐ7s"7�K�h����
C}�v�/j'�ڒ,5��p�f�2tE~���R,�mQ\�����E#0�C5�z�ݸ��l؞	1�D=����#-t� QF��ꁸ��N�дE��Ymur��)���ŋ���h�XLc�N�v��.�x��S>�c>��ij,��M�(��N5�s���{V+�V��Z��[���}6C��@���B֏�iȀ1̅v̍o��+��MW��!���&�y&����7qc��*�+J$xE�Gl���UD廂4#5\;�3��g�{"2��y�|�U2w��F+��b�������q�%K��i�I��v�,��h���O�x ��05��ŀ��l�0B5DU]�ȶ[C�45Zz��شL�<��s��E�z�lf�,m���Z�������C�7bV�K�q	�� ���i`�u�O64�H!�R�!P`{�oB6]jC��/3b�Rw6V�9c�lґ���d{��Њ53r�}p�9�����o	�ঌ�'�ݭoI� ��{��
�*�h�e� qz��E�i��B q8Mhc�����b�;�PR������X7IX:�@Og=�
��F1��	ﴜ���A&� ��<J��}�wn��/ˈ����U2�� R�ػ���3_��;X^.x����4���ы}�k�� M�Vs���3����/)z��:{8������¾.rQW`���%B��m��d1�G^~�*�4J�L�/�89B� �w�}F���M�`t8���>�M8���2�X�AL�r;��m+=�7�g��{<�=*�d
����V�P�*qp����e�ݠ�Lo��,�)_����bo͜��Sb�q�����)�k�W��[5 �b�e��Ԗ�pQwMQ��%�W�&�K�K�c+�A�S�fe�-�*;G:�t��]M�]o����P,�~v�iC�N����������a�6]�	���!Y,�C�����kp�j�#�[W|��.`�*jܮD0��n�/�(�O�!����L�M��^$d�l����$�Y`�q���GYῒhc����i�^>�E?�,�&ǘ_ss<l1��G�[0(^$u�M��8b
���G��K�����6��{Y�H�L��ML�ǩz�Kh(��Q
i>�̕Ƽ��$��4d&u�����Q �Wy�$!��򣓨�zr�
>/Xq�@�����Q�g��&L������T�1�)��%oG�����xH�_E��nIˊ�+�7P�3�:6��p�~�<�^5Բ58����n{����~�PY�T�$ގ�b�l�k��s&ʎ�;��G�u�뒐���b��h��J nr1�:��fܲ�~[�$�}�?�GQ��9X�ӊ3,h������aÁh�$�U��)�����r�~�n>0|u4q�RHJq\s�/�h%4�ǐ�k~U:���U�`Lg�Y:Wj�10�֫�g���U�ߍ����Vq����G�o������y���9�>�UgFѓ�&ނ*��J��7S[8`�t ix��$O~G����hz��! |���=|�-��h��5��0�Y�gp5����m�gJK[�2
��ln�&�1c�.�Lԟ.�N�����&=Z��GAq�c5|�녍A��O��|D�ҝ�<zZ�����j`�̊~���`��g�j�zw�=��cʵ͆k�KM� 5C���
��Yi����~�|��H�/]IJ��@�
�B�S���N+B�X��& �n�$@Аb�w����	���6dM cD��]T����S�ʳ�U�Ț�QS�F� 3�<ɹ�r2�Q�*�=dE)g��j����h�����0T`�ڻC�M)޺2�cB����u:	e߻S=�����Pa��Xg`PIm1j(؎��</�I{o��P���]�_G&畢�i�ly�"oO7��8d(F4+Q���C���I=X�� v��I�I@���M�	����P�Qt��۷�Z��;
��U�L��$�|iy&���FNf�����X���8�@}�w:Az5�=�Z]~�Z�FXo�`q�6S����:n}R��]#tsr��f��)B4�.��_׾�F7:��F0~�l�;��;}.
�Փ�h��w��W�.~/�|)�2��^JB���p����]@x�(��rJ-
���B��:��R��V[�Q���7���2F⛀}#���$�ҋ?�ovn�&��t��8f3�����AC��C�� "�p�X���ܕ���S�a��߼��5	�����<D��8�h��aw#�p���:dnh��6� g��|a��*�m¤	a(<L��2�`�X��|nT৉ۡ'�b��-?�eFUm?�c]��|�gs�㚑�~��g6�n;�h2B�kC;4�,4Zr8w��ܞܠ���Ò26���A�/fӱ�A�_W��xo<��������Ku��Dk2�#�Ӹ��Yx�W�"�7�%̆�Hou�EK�y|AX}�-�����4����ѿ��3 �ʇ��k/j�b<��_���[3n��{8B�>zQ����x8(�����A�!�-�2	)[�6��X���kB���&IƄ�@�>�����y�#��d*4�20pdC��R\���}T�f�N�D����T������!��z%/`�Td�&�3"�[-� ���8��~𝷢v&��W�O{4�π�3UI&���ښ�4`�:��y,M��k΅������v�j*�3���-8�fΪKb̶@ݙD�3�"��U��I�mۗg�r��#ըZ�s���d6z�C��j�f������m���W|�u������\�i��$9��'�Z+O��"�8���!���6�	z��z�Nw�Q�\���lL��uY<�X�b���ţ����9�_�&�����$���ef��;�t@����0�˟z֥+�����n��C�ӑ���kY�*7˕H�%�/wT���:�b�Y*���xcLk[���C���o��yx4�̔0ȥ5�Z����B����q��w_iS�+��6c�����L�:ˇa�ٱjJ{�kK�._�N����ִ�^�"�m6��-h_	��q���9��*]����D#2�tAy�u
Ze�U�.���K��" ��չ�ZmZ��!����D�tx�:]`����0���C�ĥʬ��̺_��¿�[�2p�Fh�!K3�p��rr�뾩]4�EΦ���+�3&�}q�Hv�9���UC�i����+]`��
����U.��r�fdĖ}�Ѯ�� |H����q���6�����ep��w�XLC;W���L��F�	_a��z��)?�Vp�7�6����#�IfQ�u��v؁���v�4�{%��+>!��Kkv
�������+=4Q��ǩycc��h������ ��BΡ,Ԩo��
��*zȓ%^�z�Gَ �K&�$��>���W������]�ܣ-�3�m9cuc8.I��z�{Ѽ�d.E>�kk�%P,J#�
,
s[ 	�����h�]���[���Y�3��N�i��Kc��ޔ�%����٦ �[�>�4<͍���|�L�AFBђ����]sp0�J`ܗܴ�f��#G�Ok#-�;�5?GK�|!\�Z)z���t����M(�XB�����4'����C�#�10";�]ơ�m+��/4QR�J��uX�x�h�����O�9
��^��4`e*��}f�����f�b$�9�RG����h�#R��}��i��s��խ"��a��0�å�/��0E�(_�430T?dI�W$R�¿�s�hF�dkW��BX���(���r�-�.��e���R��B)���?Ep�6�!� �>,��C?�߬���|V�<�֭)A�2����B���/J����� pjX���s1B�{da�g帙�ձ1���E v4��T�*��F�# #֎��u�iFQQ[��򜭶 �^��X"7�ik���No�R��0���WaZE�f��Z� �p#Oy����?���|! ��q\Q4M�F��m7[ٟ\�ˇ�f6J�5��Ld�������m�����D�ʐ��l��Y"ѷ�/E6�Σs��}��O�옌��*��b��Y���a?rj b��U�^��,��h_c�������c0Ea����"UE`�{�	>�$��#�`�_���-:�Hx�;1>�����F}ޛ��F��5�P��JW�yސ̇���ڽ�E@q�7Qal{�:x�W���r�����^�����R�Ï1�TQďc�-ј<�eG�IrІ�3���D�M9��P[j�O�1�Ϩ�SP��(x�9֑XA�D�����2[��gV%�Bb1EA,A�6��e��=�XP�3�V�5�����&�%7Јn*7�p��w�C�9��l��������^؇�M�H'Ɛ�.v=�&�X�7Q,,�z�¦�9Վ��X�$T7kN
!PO�:<9�6�Ņl��G��[�J{�ڄ����%�YO��S
gą�@�.���&l���Y$� �
�R��gtւh-0����m�?�!���φ#<��A��U#3�����J�!���5��Om�/m��i�����~nՐ߳q�h��~W\�U��Q�!��.}V�Cا�h���<����Sv����%}j�����zS��!�U����1�ߤCE��:��^^�Z�{���(
Uo����.��7d�>n�8b`���VI�H�r;�5mw�ѱ1qg��nM� �Xwn�>}*-��$>�飐�﹇@��⢚����:�լVg�uU�f���8�#Z2\�Y�Xh���[���<3��� �O��������� �@coo"�@��5E5>i���Zz"����b���
<�F��߫{�\={�,�Z�3d6��I�+�K��"vvi5���s<�WV4<�^�P �!��!�-�kO�P�w���s2������F���P7��}��P�h�J�1��?|����J���J�&�c���L��	�xr�*�Hۻ������[ߓ�����S��%�A��S��&��m1m������=���E9~�C�QHN�I��7�T�6�̋������j$���.�`��`k\���ΊY��N�[e���A�h�Kfi�c�x&�����4�3f����
�٩��I����nt55Lt E,�-�����"���98��⩊��ۙ�Z�^�����/�4!K����b��C�Jw5R>+p��J<�θ�t���Sc�W�lإ8�=q�P>(a�yvH�%Ǥѕ{9?x��X��l��N<߭�2�Y����\ŏˤ�J��{ɖ�;f�.�#�>"���0n��-on%CR���ɉ�צ��`�P���'=����)Ǽ�����Z����/%�O�{݇l��u>�YN�i�pK����S��d�YhA�G*��E�e�  ��+��Q�L�f�����a���ʍ��g_=�Q�	������=nc�#9���;w�_t��(qP&�t��aj:=��jd��ӗ_�B��C2�/��z#G����%Ao5WЛ�K��SI! ����^V���� �&a h)��F/�6���	��G0�Ir�>�K�I�L�,F��;KY��u �Rv)ӕ�u$����K�"̎f?t1S��5]e��l�	�p�駛_e+�i����Budc!?�
��Hā�%��z�"Ѓa�3D-�&�O^�a���9�F��P"��ɲB��W��YpTv⽢�ne�c��D� 5�5�
I��,,��ٯ��u6�ࣷf�i��q����ECSZ.���,�c��Pz������:ʟ��mH��X���(��T���QN�� �%��g�e �c�~72�+N�g7~��*w�'~>� -�_i�s���j�LZ�04�u�Q�Y]d(_b���G|{<�.	M3�p�@�b�*7��"��>h艂7�``C��~d�8Xɹ)p�0{W��/�Fr�?����9����BZ"#
PD7��7Z	/;������Wdí�*7�����L�D�	1�NGj�if3lN16�B�Ig�e~��v�}0h��)���2=�����}��.8[�^�j�b8/з�4sYљ���0���v ���jA+HT���)qس�K�XϚw����+�g�H4�M�<,����J���F��� �3���Xw�:M��%y�J8?�j¢��2m��^����fc��zf_؛jR��%�c��^%%H.�":��VZ�^W�o�I]Wg�$s�;\uxS i���-�v�s1lD�"T��ȫ��|�7�v?s`��?Ȍ�˶K�r�E���4I}��.*�����`�B����h�Dٚ�L=��γ��y>��ۥ�i��,�jb�HT���]�l�q��k�o4��:��n���N@��[�6��K�d����EP�qۣ�sT<2E
sҼ82C�@ז�a�Y&X�S���w,X�C��
��/C4�bE�q5�$�+���>�b .��N�@�c����0kV��C�V�Y)Wi�z4�&QlP@y��]P�� ��B�8RK�4�߆�c���E�z�����R� ��ն�J�M�iDw)����߃W�O��T��f���.��6�.|Tm���Z��'	�[��ԡ��HS/�}�,|@]Ӡ�	I�S��N�����^�8���W�2u���`UU7k����d�F����B��ܻB�ӡ�����^ZI���LG��_���$"2��'�"�	d�.*�wD<�Dp�k|��)�_HP*�Sx��Ѹ���\�H��9�v�u��������A;}=b�a�������*bm�� �(^΍���t�w:)�{
 q<~��{ؽ+����H�*!l�L�=���ڍj
�ϚY��X���o�{���4_Bw6�'#����ÕE
+e�η&j����^6����Y�.S�N���Z�e�]��J�<�7h�pΡ�7/�ApH��Lf�`���*���q�WA��z�y޷џ���W���G���yq��+���v�9G�W'�ί���P�-�P��'��!���71
����B'+��@���p��yd�ţ�����������<1C_.k4f�#�3�2����W���H0@���O�s�W�T�*dZ�r�òx�hK���a���vj�[M�V�����-�n���A�#�µ��Z����E��#��Ѽ����t���>���Ep՜Rp��I�Wk�cD��-X�;l��{��6����%NbA~����|����˩V��x�;�q��3e�n����AtPX������M.^�dr�lC#K%�` ����=x�ɫu{ʣ5)��#io����q�:���]¼�L6>6X�vw��'Q�-�ͥ��1X�K���]�=z�=�?2.����_Ǔ����?p��ԑ(�t=���q��}^M�"'���yU����f),�/��+��2t�,��'m�sE���=��D�z��kϏׁ.�5�ib?���	zB�?��&����~"~�^JC7�+�O`+&����������Ё�|�|5��Gn�a�¬�5�������~�LPM�oI�K�C{���QD��ze���L��Қ-���7ȕ�݁�6��v%3����'q��~�Z��*���4z�����6ă�}��S^;C��ݾh�
��1S�M	�'��isw1dt���a��U����^|�s�^�`Q Zα����v�����T	)OQ~Ư��׳H��U��^�K�V�e�, 	��ҋ�z�<��S��˘���/T��f�M/����Px�{��%�x��m��;�5&S"�W��{��;3��Ԑ��a�0���yޘ�[�x\۴��[��{G�3$���_<?@�C �?jZ���$���xU+e�("�]aQq��X~�ƒy�JF��qg)W38�w{�5K����(��@����W�+^�۔���,�R�*���@�U�9�x*��R�CUz�Z} ���k�5�iF�ۛ�f�֓����+ j�r�)��htI@�����h*��ֺ�&�^(��F\kB��# E7��V|�PM�AN���f�qd���S��D;f�v�2����
hZ���<�Qj-��SD��`�R�Ҿg�m���V62P|���J�s���/�����ʆw��U�p���I�u�� ��+4Uc��W�
ي}�����:&^�:X�]�d�XXB��x� ��gmRhq*o�ˊ4S<5_y���t��~$w��;#�7�����?ZT�-�%@o��))�Q�2�A�ʵ����e]�'2WUf�*�U��E �����BWߪ��6d�l|T���x/'�y�/ڤ"P�)E�D;X�Qw$B�J-���
��b�i������1�����O�M\2XձA�DGe�EG��KfL��e�� ���bq�6ڃ801�U&Ҋ�%D7���}4�:�4�'�l	��ꮶz�U|�(MdЙ���j�߳�Q�dݜ"���a"�|�z���U�H֜������Ef�'���@��i�=�3`t"ѳ3~,/.�"@����tT(��,V�~B�_��i��� ul�re}xVS��bFA�>�y��:�] =JtO�%/֊�F-ķޫA��v��CnA�Ƽ��
�y�@NX���[�@1>�R�Ɛ�a
�պHz�(������8����ýn��H���q����"�լDM���*,.��z
�Mk�6�S�VT	6��&]S+��+���5|���"0(e9|�Ua��Kܡ�J�<P	�1F�������#�  f��h�q)T�a�7��!��c�s�,$��}���y��)����7��N�l^����ʗo7jg�Y^��Et�"y\���v~�u$�lⶏj�@k og��ᣔ�A�0=����e�H������:$9�u)3!���U���7��% �(�[A�s��#4&���>��Y�,���Pc}�7�
��cO�,�oWZ?��e��p�2����KOk��k���G��-��,�A��z���
��v\\��&sg��[���H2���^�Bb*;����YK*]����<�F���$8�J�e�t\��!�.�f	F<��X�_)����C[q-�Plc$O�A��Z�CAFl�(���;��	�]#'�������\5R���&w:�&��]DL�PƴN�Se6�N*�'����F��X��!��Q4|����}'b~�,v��rږ�O)�����l��E����P�ߦ�U�'�:�87>�"��/�4�K�`�x"s~ߢc?�:E��ȁy��PEa�0W��G�Y曲����{v�΍0Tz�E�jz�WI��s3 �/;�1h>o�#Sߤ��=�)��CN��?���'���-B3,O�Xy
a��&Y�hNs��W�g�[��w��!64��0U:@cC��Ⅹe���8Ǹ���;sK ��2za��i\�m+�KĹCUhZ�Rمx�"�v �ԝ�2�	�т���Zq�z�� uTGf�9�1 �s�MYF᫜�/�o�9��F'�obO0�olH,+
#-ͧ*��m���H�n��秭�l�w��WlTE�_��o����+:�9��{y�� �n�uP�d����Q�a1q��u�P\��ReTtc����t��iѧV���w�0� CnpI�R���Wm=գ1ze�p��`.pHb:�WH��L�ĕfY�&��'���c�F� #7|1��AHc*}�I~H)�i�d�q��3fK������O���W/q}=�C�Ŕׁ�V� �����v���j�-d��,:5�lrj�1�~�1��V�<c�G�����8@�:���
<P���	K�b/SǡJ�ϭ?�R��v�L�`PՕ��?n���b߶)�(d�a��.�hW�X���/@�>u���x9��\��%��x��a����BrC_�Eu��I�´'��v/x�*��'�D��C0��|��C�D��>Q_� 7��'m! �W�Ʌ�)6,��w\�5�?�
�6��y���R�`�"R:nP��D���@�6K��&Cm��{Is�5q����zRs��S,+��9�u����Ƕ����_<hpꌐX}������"��ڪ���G2��A5!�Qq_�����+6uf���/�1�����W���E�;�]B�-�t>�H����Њ=UFv)�$����� F"��Uɑ��܏���Y�Y��&+����7I�B��z^�!�u�S�%JrF���,J������%�ML^g|G< ��t"��R#=�Z0+���y�� /�c���^2�̎_E�~�@�Y�~a#"'r��&9ܗم�� �������4D�&���Y!ZꦰƵ�L<5j��9�ZH�jr
��j���dF��vuW�߮�YUq)M*3����~��:�Jlh��ع��G���(���x �8���ѱ�Hs�)2獧 ����s�^Dz���4�'h���L����Uqzn�U���U{�_�><�����=�a��.݉�#]� ��/�S�u<5O��������� ]8�ϴ�O��M!��͏�g����.�麂���h�B��D���T�����:iPqi��e��&:t`���/�`�Or� ��*�����RF�3��t������r\����M�ݧHh�T�=o�䐀F������j��%�]��a����E&f��΄�c��-����)>׾�.0���rP�f~ڜ�6a�_��|y��"l�9�;�o�u8|�����<��+�58��:m
���"�*5��F/8���w��U�@�9� j��ڿH����3h���Ɒ��pV�UGص��y:12b�z�j\T����l���Rϙ4B��By�ױm�d��M�I'H�!�c���V��%��2�֫�5M�2ǻ�&�$��C�H�?!0#3Q���nB���D��hg��a n�죳�tFūd-�/�8_d��b���M��q���뭸�`�J?��+#*����~9��t)c�+�"�vBܶ����.3M��]`5�2zS����������(�72>m��O�+8��kvV�~� ���l���Ѓ��y3o��a�5��4�-X�ͧ:7b�E�lE�e?�ΰ��3�Mr�	���~a\Bˡ��+���]I�Q�G�y,�
�����
rɣ�ʮB}\��q�i�K�F
A��Ş�s�E5'��XV�iB�p�*��[SG��2�4�`���I:��!��4�Y��ip�5��|.wRaD5��y�\�A��s�C����+5�!�rɍ��, ������CZ�N�%8ݐ����%q�1�U&M����¥��̽ w�jR~�=��U3b0�7�3����U��o+,�t��{`�n�nl�srQ�>,'��\�UX�/4�
	o�����)����`�)B�4�Z��6b%i0`��Ni��'�Gk�3k���]�)!��Vo�i���WGTִO�q�ئ�β[U�n��>�����`r�%�w.���d�G�$�G詿�D��jU�*�f
���i��o���S����SV+B���L���/��u�:x�M�G�B��:E��2���g�[L��qO����o�K�e�i;uZ ̤��-��O@u��F��)�ǀ�0�Kw�@8�f� ���'��m?���t�S���Px�_mTk��{�D�DKn��Kn�a�4(J���L	A��jJ$O���:�|���U]_b�8uh�)��H@�8����X�5�c��bC�Q�+pn���f�Ě>�e���"4-+����V{�4�tUC�c�2�w�[m��
��RQ���>���������w5�d]���h"~�ٛ�G�-4�A�@�P���2������p���Y3i�j..M�-J:�j�������|a2�����hޣ� q��U�<�Ӫ��X�?E�5S���a~ݢ��-~�  �<Ң��8p�`:n���V9!>������:~JPM��!����,��k��H�mc��Ėɹe�g���Q��&<s���;J��}يV�qc�*�����0����ht�+��H�Sf/�?K�hܓ��L!�q-TMY�����]���*!ow�T'�{�4����+ݬB�jv;�	U��4�'[�yMB.Ӱ"G���4�_��' 6�}�$-ZR:�t�P'�]�2�r/��=A�էI\�h�@��y��5X�i��sX3��P12r ����后������Y�y��ֹ�i>�և���6�
%����k<G�z�Z�e����-7�,)�')g�]46�TM��m��%���L���'�x=v�ē�(�u�D,~3�w�t�����Kf���r�k�
��_%kO
�<rEA5 �����R@ݩ�o�(��P��Qڱ�N�O��b#Ea*��!;��H`&T�xb2-V�2-2t��1�1@����B:v���FY�y&����Z��㌈z<�a[�T�X���.��e� '�"��>WƥCFXG4\��ql]43�4�G3�[/%^��88r9pG�s&��UìY���T�RvF &X���G��h�ԗ�U��J�r?��,bC���5$�?ǿ���&�0UA��	��<wF"�����-�"1�h_O�%���������`_W&r�4��ׂ��0�F���TM�/|����dZ��X~{ �E�B�H�����#�]�jJ�����J�iW�X���+z|=�!�>������Z�1T��� �Ă��
X���u���f�pM� �EL�c[W6�u�vP����!s�K�Z F�7=�iZ��"/O(�v�ڋ+#���X�O�i�G@����ݧ��B�K2k�F�[.6K�`:r��]��j�� ���%0 1v�ҧ���_�/+�������3Ƙ.��@�o%��S��(e��ˁ'2��19z��
n��ʿu�y�a����dp�һV
ʜ�]�B��Njͬ�N'�'w�lAᷘERѹZT��^��(���5Oou��t�����g������4�����4F4".9�9�+W�5๪	���8gEd
M�]ż:I��;��c�&m�����`�I�=�ل�$QXӳ�M����z�Q��g�A�Uq�Ӷ	����Y&*LD�����FWNu�RZS6�L�5Gȿ8Y��$m� �H#/�����?&��ڑm3˷s���'���fHk���Q���ת_��W��^w��0���;�����n���1:=H����ŭ��ј��A	��a<����5��(Fs�tF���4�.z��o��?�h��z���Wr�;�G�b2D�e�ܦd �`��gv��������Nc1N�`����/�V�OoG��τx�Y&�Xc��[7nS-�%��(���;�t+E�,1�Nj�mE�IH��e�݅.����B���4�3�O}0�5Ľi�
)w����֥���G����.�d��I0��xS�mK[]UM('S՝�s�b�D�3*��ⴸ�T�.�	|V��QU"���� �X����Hl^�EJ�h����GOʮ�Z��/&�g��!�7qx���9��X�5�,=h���Q�7�<}_�%�Bg	�U ��E���k;UB�g���+v��v,h$¦�(�g����"=�#�1�����@�ɈԢ1��ׂ!8�5���Q����,H5v�z=w8��+/P�����>�� ̟��;�E�{.��eh����F����J��[�ۍ�!en<0��Y[�� �<��橏�D:w)��[����On�TQ7��rhi:=5rv=��G@���/�]:���x"5���N�gIS���T`�����w�B� �#��e=u�Cc�y� �Z��Fw�S:���7���>�E�t�RS �+뾟l(�b�]$���J����a��U��i�N"�@�N�4a�R�-�a^q��!����	N���G��J������$�,J ͿJ�v��+��F"]~��Af�6��w' ��O�I�痘��P~���>�N�W�
>����Q��J	N���,.�E�;��D�߀�v{���e2̀�|��l�'-���P��bs�ۖ���Z�Z���������GK��Fde��i�v *m]�&�~1�����]����Įb�j��4�l)WSo�n)�իq�(�O���,���$m}E��2w�Q �6��v���P`�y#���}.�f����+H���V*�F=7G�A"J�c���cz4yB ��wD9��^����4=�# }3�sP���e����;�(+�|�@#
�L��
n.�řތ�3BM@j3�	���+1(n�˴P��� �D�H()S�n���lXA@��\��U_������0�8��-���]��)��R��'�'+VT�����᫾�}�)�4�7X�7t���8��:R�c�����WPiD�`=H��EM�UM�jh��VQ�SX��������sMi���f������_�F�|��d��C{���X���י��~��z^y1B�MR{(����CXU��-����^�[���%=^��q�_��f%!ͱj6*��[��z�)�ߒ���M�v�Ɵa��]�k5�L0�c�kY��%��|��qy6/���]���Nh/]f�rV1���������X4V�|p��\���@z���~���.�ܮ�M���aH���ʋWq�������J���/W�[�)�$�5|ƺ���LK���{8-J��V
�k� ��'�`+7��#�� .���2�:%�{ɯ���6�!aQ�ѺZ� ��:�Ы���b*��3�����Z�1�o�;�KDgt�W�5e��Q�&"�{?�"���!�0�-�*�c��&��1��²�Q|��+=c�����1s��=n	hM�A��11[�K6�MjC�ST*m���@��]�E��n����Y
i��A�\G���>����ig�~[\M��"w�q� �+	*ݟ�!Pݒ�+����қ�Ǘ�g�HǎDwb��|C����aq�z�p�:��S��B��Ur�*�iC�L&�����_PFsП,��6 �PSI�,����r�Ur!����j�WcH�/_�4ҹc.�1�2-���J)pJ� ED����|���{ w��k���u ٝI�P�e륹���������h����FowK�E��xIv��PNKoq`�%�`�����M��zt�V��I��:�`	>�O�����t���: ��ؐYQW�M����ӛ�N�����`7|�6!��4��T�{B%ol�M� �59ޜݛ�1DNK,p��O�|��;��~&s�[Q��D���8lbRl���Y�t�4�Ww�^Ǟ��=�Ȁ}qE�e�R��Z���ƶ[�R��y�I����hD	�)�@�lg#5�7]��Ƽ��@JZh~���fz���G�8Ώo��_r�'E/H�Yc�Fc�fm9����B���dF:\�_��ץ���|$S�	(��W���a����F��]m������?��x���=e�i��~�������u�����Q�
�0��Ճ�O�K*R��v����T�o�Y�?��`jP���ұ�HıC��A��?L 9��{�A[�}����G)�u8ڪH�nn]�`ߎp��5E�$��.AUt�m�P�"��X9+�;���ɱt��3�n���p��n#$&	�#��]0�"�����$?����������Ё��(�blҴR���w�-�G�5�-���Ϋ �T�Z3�=��$G�À�g��n�^�7i��	��� ��]����h,�EX �0^jK���s�z�R>����Km�=r�k� ]�&�/��4آ����R[Au�D;�u�
������-�p�q7N�wi{�,�*�����*��=)Ɖ�
�P�-������NV��} �Gå
��(!�F�pVB�+��8&�?C'	4��F:�%2��}{9f�o��3-��J�C�nnXJ�xr��2,g���"C٘>�5�/���p9.�݆� *S�BD��S؁������P��:�g���N�N�^Gu�z��.*�$��S~tUYv��}�N��s�ȝ(�o!,�$�"��HX�E2Y��m�O��l�t�H�W�)��<�/Hu�_=���"�~{�����_�ˋi��`nȁy�1FЊ�<22���q�%΋Ɉ.�b�oOU�ٍʨ)"D��/��9-:z�3�c�43j��4i&��K1�g
]]��]a�0�&��y/����xr〷r{E��㐹� #�[}��9���{��K�&*|�������h!�I��r��4|>(!�/���M;��Et�v:�/ѿ�{n*|[��[�-�dS[~����U	�~{o.O!ׇ�Xֵ?*\�2_
*�L��1��N7���˧=����X!L��@��ͪ��� t@�		b���:���ͦ�r�T=���ݵ��X
�Y&o�Gn�٪<��h�V� ����z�(`)��Ue}�[�x����aVsgi�浣2)�	�W�z�I����M��[�/A�h�TU =K[[m�����%��>�<��uQ��	,�z3��G���B����1b��0��>�ppS����x@.��V!vE(�8� #c���4/��К��O���/U��0��;����%i�S&���;�V��� ��#L(��
����S�'�\�`�ݏ�8�>" 0�������/��Q�����br^\����w�d�nΑ��j
����6�B*2��o���7#��2�#O�ө��w��y��^y��s	���Q:ӲL#�h%M��Iԫ052X�P��^�Vo��o�gJ�����ٷ5�M#5Ѭy#�"i�m���E���]N����/E�c�6M��ߎ��Q3�_���Ǉ�l��x3eRA����]zV����.�ٰp'�����$�e�v��<WUu�� �h��iL��{qu�bA{ycL��{����e����J��0^���[�t�x��Kr������*�Pt}6�kuR	;Uʿ��Mw���3�{Z���3�qՕ�h�p�W���[���0��D2t;I���>l����2~c&�팦���
��gt�&�z�	��4�^�V����_J?S ��mʳrbS�佫a���Y� ����ĕ����k�J>���W��/�>/���_>�7�J*��)\b�xT�{Xf�"Ϝ���ER�p��Λ(�,~��$�ؐ�(Ÿ�$�<��j�8�+��E���2݃K#�>@�b N
:X�Nn�H^6+�h�$>I��sug���i|.�z�E,���5�G6N:8<�Ɲ�%�G���p'��gg������	�:[���
�Y����8�R���K D�x����'�x�t�VYJ޹Y�Hl�������!^7���6/Ԗg�
�͍�dٗ�]���n-f�'�"��Mn5��NW�����;B�m�S��9T�e?�c�^2�Y����Z�D��E��k�g3������+0d�\��Tl��O ����!1���,T`�@y�ɓrZ�!3���Ș�O��	u�� 90g ���o�B
F%��^������1�@e�_���lKLu�Bxv%��������02���$p/��
7�l���Ҭf';+��e���f��9�WOct,hz�v�+{�7�,����Y*������Z]�����,Q�Y2��j/���{yVnK���"��-L���W�%���l.�r[=�Q`5���$~-O���[5��tQ�'mN���� ��4�JR�C���qf���=��NX�8[�� ��Fy�e{¿Cs��j�V{.�L>��K�_�_��2>��6n�c/��z����^^�Kfl������{
� Ua�i�9���]to=\0 ��q��⑞q��J����s]��=��_�a�ʴ��nN9'`Dg>��h�z�a~�v_P��ڜ�_�*���v�M����I�,�~98_ 	�C,�F���6�$�Q��7�sz���n�g�?��}�Ԅ���}[mgf�1��+�,,�΃�yT�SC��71���婒Ώ#�<ܛA&jn�N������ۦ΂8�����Y?���5���oM�a��P���I�ގ��[?dķ�H��>��脐���#	��g�"%3�@n��\qH�e)�D�n��z�|��R�&������+,��/5���HJa���_.7��1���$���N����+(`F[k-� �7��ߏe��XS��C8�3e@��aW��-sC������~�IjNX�\��]�yO��d�P��(�%��:Z�uɌvg;���(�������-�<�0)���KU/D��Ӂ�^��DeS�s�2��@P`V$�G	��W�,�|$I+o#�&�Ԩ�L�W�]�Y����Ԋ�x�2��4��[���X�ؘ��(�,��Gw0�����4S����#�-��d<�@&E��i]B��Eh0�ݡ�.ht�3y@��)������>����Ƶ��&���$H"3ПVD!#�������q(�=C)��OEvL]����p��	y�CI�1�-����<_�N�Jr�Fn�"� ���b��6BR�7u�n}�p�����|Y�.���X�t�m{�.����'�9�˰T�T ��"����+n�D�_�i�}8����f\5���']!��QB(vd��"e���*i� VT
B��O�"B�Uc~-=�'n13�DG�����)wq�U���C���&�d��A�%W@j��� '���q{&ͨ�Q�������;z�R�kSty�I4�z|����8ʙhx�f��T4��=�yCi5�ڪ������Q�S	�� 4���@��W�3�V�L�v+��\��c��I�i��cA�ʫ��g4�?i�V\��o�`�������O�x�]����P�6!�^!��P0���������a]�W^�UIRO��:�"�jt�}���H�.A	�#ޣ�b��β�� s��%��р���YYo
�z�bo�^AGz
@��� �����Ľ�3�����%�BĈ@_�q)�]=7HNE���R����CU�%N�&����
�<[���û�/m�����2=��)�;��^M�,�܂~�!�����'[z�Lo�t�l�+YgdJ��$��RTs�Z`�<�?њ��90�ϕ�IO�P��<�q�a^�6Hj����J�P���#�Sn��ER���U���zk�N摳4��/�<���7���#j�آx�b�a��gS�����	�
 ��<+���rl7�O���� ����X�t��ON��,W�.1(5t٧>�0S���?_�Z� >,���O��r������9�<����9�w�b��ٍN�|$5������nN},���x~�L�,�a�b��l�	����lY�N�>��f�	W� ���WUz���>���1B�c��{}�B#|Y��++aA5�t�W�ߝ�:'ڹ��.2�I<D��`����2ƙ���l���Č�d�ܯ�p��.ż�Y�7䏵Ɓ�&���Jx�Eu7͒��
�J����+'ը���<�+-���� N��5]*V���^��C0!U�"���`�j����5�lOx�y�1�;6ӷ3;5�W�4���D��	u�C��`�%�3�e��L�;L[�������gH�J��@�qNņ�>���*�t0�B{pq�`K��CpB!�G��ԡ Vx۾m�?9�B9��f4fq�Q ���RH�	4�T ��Ț�0_v�k���)�͋Swl'�oo-��{�sh�=�=]
BWߪ;�K�I���˥. B�B(�GR:t������S�m�����[FV|_���y��?��V�K�UH���XTS �X"�a�<F��E�3Ƹ ��I�Q� ��`�n⍧(.�?�ڡ7�!	":6݄h�F�6O�+�>�o�������5��;Gu/���lw�<��n�=�6x� �+?�0�÷i��A�[�ZC��D�O�$�u"u��k:�C��ժ�����` ��EyJ_�D���A�f�eU��?�.�Mҟ����f���0���߳��
 t�2����t��,2SJ{!�e��E�Njs�4r�>���>���'�"�R.�)��)#STp[=�D�{<Y�nS��ERl�p�(�7q"�U*��av���ĔU�r��c8������a�h0����%�X��4
�Xo:i�%��s���0���۫���c�ɂ��� ������8˂'&"�$C����V�<=��w�G��1}`�yp>�l���\�=,�$;�E�cK�^1��y�o���Ie	���0\�1�!����T���0&!��D}�rep��F����@O�7�S59���	In �O���uj�i��)���.�ܼ�5�=Vz��) b�''x�ޒlK��P�e�I/�	�.�K��<_��hW�����,�,P(ǩP|UVZ&l�̡/�ï�)��NY�]}�a"����#ֈ��2��*��B9�<E��x1w�������:��� �4%��a�������E�a�`��������@\#���v0L�Hl �-���NI'mmm���Q# EG�Iv����S;�ʬ����Z?q
�ƕ�~>��=x�f���u�-��{lƗoBGc��
��|}�Q+T�|i\0#�m.p�^�%��s�v6q=k*v
ie�Я�s�\��Dl`P����D��8@�=&�e���GSj���ْ<C�����|f�n9Tm�������H:������}�e�O�^Qs���oJX[�В�n��z�t�i��:m���]^��k6�u¦���ᯯ#<��M'qNhW�������
úƤF�`��~�DzWo_=��Ƶfi
��:zG�����7�{�>���Ic�d 
y���q�à����rU���cq3ꏎ-E�'<>��u������Z�N�;Е}�P|�H��9w��FI�=��X�x�֚->��=(D��;3�t�/�7��1�E�2��,�@�(+���լ�t���롰�w7'nO��d�9�Q�ND,O�1]�:@;��i�y[{ѣ��(�J<�`]��ԉ5����O����Qx����� ��-�g�",w�o8T�-���-L��x��}�c����)���?�ah-.t�#�e�G5�L�u(���;���q%̿�Psn8�y4^�!@E��)�uK����)ݷ?¤�>G��p�3S{c[�_G0�"�z`���+�Tzo��y�\��X���h'9�pMF��iU���|����7�}����Ҿ�8'hBEJ��h0J�1=Ү��o�[b���~��p �n�ш!#-&vт���D���S�)�l���{=]��sgS�������O�$ه�
ᷰLH'������-���(��J�o5��ƈn��7��a�߰��buȡ�����lL4�/7�l?66�b=�����t���NI�;P�ӑ��_>(��z|~��e�����E�u�n���p]|K�a��H<*�hɿHh.~)
X@C�إ�e�@|��77�����x�:���J�q�E&
���������xp�&\H���Ԁ�Aw/s1��tAJ6��D:��j��6���d����\��x0xǿ�kщX J���!B����ddO��*>��7�qŮ��J�B(ݧ����R�O���ea��4c��*�S􁼢�a @����"'e�I�H��
/*�9e7�����ק�>m�&}���"']�~�z�m񈡟yt�R`���F2���k{+r�6�׆���Y��Xsm�QfY�6����Zُ $+�4�ha��iz����.�X͹��̈́�O�|p������ F�P�3ѣL�zm>W���.M�(���H�<KTG������М��|�w�)��6�c�2�f$8���-������wX�)���:�[X��K�$���R�-�He��d��r��,O��H-f��\���Y0C^	{��=���*m�+]կ�~�-���|`3���8�-%>G"R7��p�/���G����~�$��a>�ޟ�w	��(�Wu��В�,�B�������^hpΜ(c�;,����ޜ����g����N-K'A!����&w�4?s=q�.�ߚ}�&=k��(8;ޢ	A]d�.��.L"�)߆�z�'���k%ZQ�h���Բ]Q�z��nR�a�ic���51w�ujǑ5������1u�q�B۷����QR�Ɩذkj`����cmɯȉ�iٞ����	W�l���z����R~4~E�<����C�'�*��wM7�e�F���$�x c�6JU�1�È�x��$sq�V��*=v2,�
o����BL�0S��].���;z]���A��J�Q����VZ��Tx���_8��o��j|(Z$����bP����W�K��i�ی���BP��ty9��H��<�M�G+]*�y E񲰤��ҝ���.�B���Z�/&�}bɅ���`orh����N�1�#�����'g��y$�٬ޛ�rԑ�x����y���)e-MLcAe&dS��w�w<U&�=9�������Tv����4�"Gr9��O�!�`�����'��U| �����M�:[`ز=G�]�9^��y��s�wWzc����_�`�c[�IG���Mq���[�IMn��D��ҏt��E�8�H���xv��v\���Hi�4[�l��5RB	����τ�
�������qu��fʻ@4$���D�#H�=1���ؚ˰r�e�*/�q�nXٮ*w�N�e��s.�%*�ZZ�n8�z�{����$�N{�q�z}b�R܋�h`���u��3��g�*�=n�Lt�z�W�I�Ea��"�H�/B`�Ɂ��\^K�� d�sA�=<t�
y�Q��[��)$�S�*�I��<��Y����f�h��2�w��~)_G|�d¹��L'�%�b��%���N<+�\ju{ ��k4���L7ʬ���&�=�A�'�<����[D��6�3ie��а����9szh��O�)�'<�Wϕ�Al������o��׿������C�ۮ'��\w<Ŗi�#��(�/��y1��.�B�@��t�m� �*g�f������{O�aD]����%����������h3�]!-$Β+�Jf�?Du����� #4:�*�E�e��~V�H@E�T�y�v9_i��8N0��
�������id��fXjy]�X�,�q�%IL��P��l*05�o2LH����z[�Ģj���u���љ���~�sp�9@�dV	(�P���Ze45�͢�zߕ�A�N��#8�=�/F��~�o�(7�G�f��ڲ�~ЊG{$j�����sU�K+#r����>f0���6kǹ�<w�=���Ɇ��U@�`}�V�e��7�MH�=�y?���-���~�{��K	G��y�
^+��&�	�y�~0���T��S1�
�~:@�2.,�"�Itڬp&+ziCX��[�#������K�n��NV�.)@0Y��8�
li([�oJK��u���Z�Y�!7���5�^�T�M�ȩL��Ļ����WG[M�m��dX�9o��A8���j��o�}�|�m��U8w�X^)({˕��=�X�-�I:��P{*᪦����"��jd�O��p�l�:ג�U�C�#����{֏&l����BrU�*ξV��ol�
A�(�|�k�[ə�� �`T��e�&nE��}ן��P���U�R(Y����x"��SlP��O�Z�z�</�Ŝ�k�?�o䐁b=�M�J���۸-RS���By9���� 95��Sq�����h��M��,A��3��3v[~r�p���g�!pw㫓A���=t�α�6X0[xi��smԈ�*��x�B�܈&p�0����Bb��qPfR�B$WI��3��[��+�.\�TN(���+����;(d�37{k'���?jJ��ps��\��1 ���M?�U����o���o�6��@�+�U���^NƘ�r�dĎ������#��5�P��j��/��Vw��R�l���劅�n(��Bّ��s��/�f���]�e�:�?���ԏ�s�@^�:���D�9��>�?�ɐo�/K̜PQ�t�TH�զ�m)���KR�`^��f�3�bٸ�LVUK�7��`�
�=��ʰ�-Y%�PՆ���|a��] �lHB�����P�;�Y�h� ��}G��翟�n7��K���A��=���P��FOe����7f$�����.�p(��<ƹ�w˟�jDf��D�j-�©���U��O���m#9:f왃���a���A0DBS"VH� ��&��`ɨ�5������\�u���h{-M��v`�'s5�':?���L<���	�	��U���ֳMz��a׆�]uFA��o<*/�(���Z�����>߀�٦_վ�{�͐�+�׈٫��
�:p�Y�e�x'm�4]&1/Kx�rm�#	���J�ڌ�:�˝�1��&5riI#��c�=6��>��q�b�D	q�e���
8;1�yZ:8 c\�C��o� t
�<$*��ϐT�=}��+ɠl�(�ʹ�x�
hs�'&�6&Kѻk2���ªҴ3}�����*���I��e��-�D�tL�M���`46��<%������lev�bii�}��F	f�	�W~�DJ�^�g,�W!p\~��&M��9-�\N�J\sm8���Ϊo�� �ud�w����`��
!{���8=�}E\��H_��WWh�u�[�h�E�@��������!���)�L`��y42ҡ�R�UB{6�!� ��{�[�{/�ܜ��m��(�p��F�+�&��3�6�!�������{��YE�ݠ�?�(�ڪ����]gH�aE�����Sk��2ͣr ��\ �_���x����m��k+ε�	��1�^�C/�wZ)w(�~>�E�Jz+b����r�ݗ�R�*?�Yd�J�(9�~g]�<0H-o	 ��a,���ȏ���%ݪ�58i")	Yg��]��~����1(���~K��M��E6�T[�z��f���$8�
��X���J�KZũ��P�-:P���~0 �.Y?v_i[�:�$�}+-����R��|tT��C)FlKJދ����	,()�)o���Ɵ��D�c�,%���]�Y�W]����)���T��;�k�j~1��z��?i��	8��&Wye�k�W������Z��|N[�P�lv�i�>HD6fG��Se��[S
� �v46�/��z%�hK�q����I�b����K'��=�gɨ�=~��3�燳��+8h����gVģ���w�8����qy�د�dLb��wڽ�n[�!��x6�]U��Sp��P�GíF*=��4p�V2�"/|cH���� �!�)$��Ŷ��6n�j�����X�H@�U-+t�M{�w2���Ô~М�mH6������AG�@b��: ����ּ�g��܆>Xs��ܣc�U�k��9k8��N�ND�)�)n�8m���&�Y�Z:�ˇ�����*r����.Y	��#�R,\�78�Hf�7.�h���Q�d���Q����eK�QE;��Iixﶺ�+��%?M�<�j^]�q#W-Õj��i����ݺ�Ss3��_�;(j�W͟�Z�b��o�Y���X�U$����D]s�ӫ~���=���d?�c���^�����(��V����{k�D�����if���������G,��R�����m����� �|S��wV���pΛP֞R'^A�Ur����4�W?!���i���PZߌ�=΅���,��Xy��Np�%�va�[ș1�dzw�e��U�iV`��uiԹT�Ò��c sF���8�n9m����SN����_��s��Gnb&N9�=�h��3���� ]�ŗs2e���Ǥ�F�u�%߲���p��8�FXgj�/ș���m��P��<��?hB�% X|!Qq�y�oX뒛�������V�����[�%�ځ� E�䶰�@c�L˺����'�D�u��Jkm�������i-��^c������l��@���n\��K�A���A ��<�N/���^�A�-�J���P��Fp�~0'j�qϨW=T���x�ݒg	���F��8��q9�4����ӓA�cJ�45�+N��4��$�����i ����a��m[�%c�����2K�[Ν�ѭ��ױ�0��\�c��t��y�^��=��»�5��;�M��7R��,u�WG*�a_f.`�O� �R�7s+��D������>����w�U�0�lq�o��0)�R� )y�m�6����=��2c(�8��~5�G���h�I�;��y�U�D��[Gp=��\�n2n�������#��׹�S�t`Y9����6'nk�*��!�n��?�+#a��s�2eǄ��dڋ)B.F=܅�V�sf��b1i�8°ka�#�`��C��xy[S��"�s���E|�� �=���f1�9��O4�m_ۙ��/&6��<Z�&\H�1�R,Q���7�/^b�������L>(BϤE��&K�B�į��:qw�b2k��9��,ďGm���Y$wޝ�H�ԣ�pB�,�txj���f�&�/'l.m�:ס�v<���!��V���8<?���z�{�klH|`YI*ܠ���'�,hܱM�l�=P͎CLw�hĒ~�ָ�n�~?0R*`I���}�ب���F'�8�(��	���c&�{�=���2��ӕ2 p������
E��t7}�Ϟ�&��4°[ʫ�䋯+,cC/];$\�!f�BH�ac��ߦ6%Ȍ�~x[u�I:1��HH(��$�rM�e`�\-x�'�����͌E`�ۂ��s�)H݃6��8��G��p�5A��P��+�\'\�.yLLE
�跂7���C<���]?mr���ok���,Yr�ϧ��� B�YTz�|�? �'b�&R���t��f�5�*~t7���F��J�E��S\���z9�-�j�`�aw���vf�������Ǫ���u��Y1]�����HN��Z%�$X��1F�-Rn�}���d{���u|;{zl��
�Sg�K����BߗA�)�1?a�#
�l;���O��E�I���q�m�c@�?L���o!D����a��ǲ)�1K�W��$��.�5���TOV�|����A��}R�3#N?��������M�a���~���1�c�#^����Hǳ*����xV�1���C1��r!p8���Nl���T�U<=�WA�J���Q��]����a�|b�t�p¾�!&5Kql)��ry:��<*�j�u*��T�|�G�k�Q��H�4X[�u>WM+�������mok�#�ơ�`x��mE�_;i�x�����k1Ԣ�q�MX�@H�&Z�1Y�������2v%o�]��������=�:�,�� V���/�M����]�tVD4Ԕ���a��o��)s��QP��RO:�n,��4�|t@�HSiv#@��~��8/�B�LIsT�	,sm�/�`ǥs�����o'�h���.��*I�^�Ttj����j����F(��ME����Ó2�
�f�<�R��{��.MڥeC#�� ϕ\���5�G�-�������]<��n����'1����}{id*�ldx��)������� w?�� �>LR�J���c����Y����P��Xh�C�ո�KT�p �-�<4꺇V��f��7EY*�oN*mo�gXE���U���֠��tV�`�g�H9��/��ٵ1Ot�ȫ?tG�T�������dH*�5���B��8
ގ��U��gcpc^h�*h$M��A��Pn@6#���2D���g�3xO��S�5�i
5�ٕ�Q�*�"?6Mhe�VR�a&'C�#|���S1�V�م�~�=��:]�������T�*�x��kE�)sbRT�>���Y�w�吰O��d�F~ 2�|2:7؆���r蛉�$��dtYl )�S8���/��T���������d�y�t��=�+k+�1ŷ��n+��@���x��_����*��)�17�^,n�g1������rK�+	/�'����&ރ�yA�2&[������-e~���g��b���X���ED��	T�%���n��4V�j#�,c��di �>9_B�z�!����ie�5_��O�6��W;C�%�h��7�z8���b�Ζ{��G�������F��B+d��689��&��`K<G�mb�b�g�w�~y��x$��S�c�J,I��5?d�5����k:JbE�0r�D)/>��as�w�Q�ZN�"E����GE��T���G��� <�������#7#}ߺ4����[��0,�&�Z�<�ң�JvL�� }b݂��F|$�ο�/��n��W���0�.~��:c+���k�Y0쪝�l˅�~��l���Cu��%q\Q���R 2�>�cR�����Jj���$���EC�V�=-sO�|_�մ0��.�Dk[�$�fB��*���զ��eH�.�Ih$�h	�e�o�\�̯;cFa0�$~���&�yNt)aޝ�}����;�]Ǭm������H
P�-��b�΃ˡ1Y�[��$�r����_~��_�Iek���,Ӵ�q�"���-H��/�����V^��C�蒔�MLgd)�ZX.�I�#����ˁ�-�s��G�ԓO�S��M�~��y�y��z�ã_�bvP�%\B��8�Q�@v}��I�r?!h�'݊�Bj}_��ܳv��1�-|��Ͻ�F�f����>�� "�#:��{U)��-��.em�jzŉR��lږ)�-��E���F����KE����lm�"K�ݪ���A�2����+o�p���r)4S�햩�źQ�[���CIj�>D
�_0�lv���G���t��*-�8���H�恴���]�jw'2˰������y0��~���u��WN�$���>���&�~.�!e�����G�&���2��-��0�Hb2<�!��jz�����X!��(� ���T+d��g�4��5�{���jW�=
��+���!���2�ctpt���G�@잂��ID�!�>
�d�YT���2�$*
�E��^0�)�
��yW�$�*�4SH���uj' 
@���`%_O�@WW�d_Zy�i�<�	���of��!PBrH�͂�&�ĥN$?_/�[T�9���&�4 �	���o��՘��l�BSl�>�C�Fy��h}�L�|N`�6~������Ta��H"��f>j��S�k�Ց
���cf6gX�N��eʞUZ+���"W�f 
�2�ZI�#D4�9�:���J���v�w�a#��wNg_Xű��
�^e�N����"9�g�*8g�Y3&���=�#�<�+dl��ْ�>l��%/�z(}�fYW�Y[
��uM/J�2DL����L<I�a鮘���ŀ�b���\���3͙
oؓ�i��^uZ�Ƅ"�`Ppd[��VTepLB���q�/���~bf�1$�@u9���p��¨ΰ}��=��è��/\�!�7�h��UJ����V���U�W��Ғ5�fr*���Eyj��N)�#$հM?�sڙ]Y�Hb��]Y��@t2�6��SRˍJB�t��z4�75 F9�XnF��<y���Ž��j�ͽs�]Yp�+zh,���!��"��E�᠁��{�,���������\��WR����o�
�+w�q������Ӡ��Tn�ל�v����2���O/͖V����(�uaU���ESc�)v`����eZw����t�'�瀓�E�$�paB�X�� �o���Pmn^|l�ަ�\�g�"*��0����+me�s�Q���؅��M����>���W9۽ټ��	�����P�8
�����=�m�F�o�?9�Kjt��=g�+�k58���d*я��
��2�"u
��|�\c��^d�c�)��	��B��g�l}w�S�D}އ��Mju�<"�k�ۘ"/���=��^�L�������w8�f64��K�i�W���J:�^(�
�.��{T�{V,,���ψ���O�S�oFk�� c]N&�ۣ8Q�
@��͝$�/0�P�M�j��W�/ pa3��4������.j��"R����� ��o�=�����;��9��+t?�e|��{�����3����W'+���rp������� �y���h��?�����I�RWF����7�|&�,�z$ 6��$P|-#0��ܒ��e�A7� ����>���pd�Ip���S��}ť���
������J�&=�*����(d��������?�[i7\�f*�R#�eH�q}��UL!���; �b�����0���Y��j�~;�2��V���p�����]�<6Kw��y%]��237�°�\h�7��_�,�b��܌B6�h¸�}������!e�éS�%�#�b�K}?j�j={�3�cX;A�T��=��iP����F��~8�EI�Q��G=� xxErz������>uob��2J�����vF��5�w ���I����v���@�f+9M��l��"�a&�eǠ2]f����=¸��|�2�˰���c��uXO�j��-��D����UEH�v-#s�F �ń���ir�Q��2�lΌ[�m=��Փޱ�����X�+��h�k�l�S%�MJV��C]5�}��5�d<3Fo>�[���Z�~0_%�K��%1 EO��n�k�Qø�ϑ�۩
e�.�F�U���E\���|o��Φ���ȊZ��l�3�J��l�'�R�j��D��Z�R�/�$c\/��6b �̘�Ӭ��g�R������)���3�IW��n���hSP�:�ң��߉�.���o����>Z�pu��8��i�c�_O`~LB����G	�)��H��Gp�aQ컿Р�
�q�9<"��OI���A���Y��JrфnRj��ZM��&@���C�G���7�I!f�6����>��ʅ�A�H��o��r� �8�1����y�ȂuP�J���;C��7~��� �Kᶽ����!����t+x����l���Z�*��	����wD�d�{&�5Vmzx4If����)H�
���l�6i��B�nթ��w~�v��#S&�\�4�V�~�)����çST�2?ciE���&[1o�_/�J�����NT<}��M�M��b�h�����_˼Yg�M��k�H�uԦH����G�����7g�P��a80ŕ���jK����������L�ŷ����$�IN8[�&�X�'n��2=��.;����;5
"�'�M���`��{\G<Ǒ��j�d�LǍu�x��P0�d��)d�P����J�B��������]-�䗏f���s��`���{�Amּ���ߘ���h�As%���QH5�ck��;����v��>Ǹ�G��f�|������-���풋�q4%�Tr��q:����q��a�O�1�܂��y�M�r�j��q�zj���/8�SЩfN!���kfS�[���6Ş���-0��d� ��-f�����rG� �e���@BzeO����w\��9�Ѥ@�+�2qC���NγZ��t�դ�M��x���(Qz�c8xur��$��p.E�)��&��Q��Yx�K���U"�`鶚�n�+P��]�)������Q_���ǲ<�L�|r�c�Q�μ�}�\��

~��<�N�Ѳ;I9%�H��,����,�O���(7k���E;�*d�
�wT��^�QL�ь��%��Y!a�s�
MR����k@�0�kL0�ϐ�B��A	ש�l�
_B�N�(l�U&���/�Ά�"�۳@��߻�Es��.b�"k�C�c-�4����I�վ�*��%=.�?4��E�?�Y�D}s5�v�Z��8GcH*�h���Kl� �x)��,_�+=���E����XC�`x�/$:���A�;���A�K��$l���段2�����@V�ac��@{,�O��	�bI���I�ҏ�D�A�������v�>c�*L��3�3Aǹ��F�)A�K	�R�na�#'�]H�(�*>S ���&h�4:Gs���V����n0�M����O�؀�|��<9��;�U��Ԃ�N� ��Z��щ�xLgr�.Ɠ��q� *��dQ���^|��q�C��,Ɲ�n�0G8`1|��ߪu�Ƀx��v� �W�k�K� h�mF�u�{���
�4-�;+`�����Y�my��mI}wT�Ջ���QG�~joW�S�7��7�T���.�B�3�����e��zy^!�:�Cj��[����%93��Ә�Y?C4�d��X֌��8���na#Nv��Ou�@#Gg|�8���5fA��!!*����W7�"3�l��Ag�7�G+���{��6]��DiF�1D��@WⓊ���^��������qk�ꑻ�@($;���Nl�k ��9����A�cLH�9	������Ng�C�k^���ڞ�[%9��p�N��1��y�jq]R^��9���?@�Z�"?`���kƁ�j�Tr�Z����<����smzSz�ŭ{x�`,�)����(*Y�,�p�9�>�3?5�!q�����m�]���"��z`.ۨ+Q�����9�G�M��@b~����G��Q�1���2 ��l�ķ0���`�O^�T��}�~��U��Ff�M������3u�������,��|\@��U=,=�z�_����H X�^eCU�?� m^pį�_���=	�B�D��^-������a�م�B�xuc��3W�����GTk���S4��¬⃹:��k���=���׏�h)~v�Y���R��VPS�W¾�X�k�P���xս4��rmLG�=��^\�<m�A`���3���d4��PB�M!�b���������%�^��c����vВ�_����%~�o�0��Н*
�W��j�p�?�:p��,F3����%!䈏e������r!�.Hőo���P��5EMx�ѐ!���g� �{KXT^���8Õ�	�9&�u��eM�D���d〗J5Rne^t�:�ö˾��5E0ƨi�N�5���kɷ(�8~�وҨ��C����Ĝ��S��u�q��ӹ�х�4��f��wl�wO�2��~���/Q۵�� �4��P��<���$�y�|Y����K��oZ�	��`������Ӓ��`	j��h��ugH�ĳo7���6KG�O�gr��^f��R"xff%������6�z%���^�M��mw�i�p�Ɂ��.��l��5��5�L�l�[�t��>k��/C��x}0ZH ����D\q�d9@6�[b
���b݌�p�Ҳ�ڿZ?��u5kN���ظ�Eթ�XYsyvh��P�._���i��������q��:5��A��y�jt1�8�N�� �wB������ؿ"n�pV=��b	�N0e��E����j"�X��(�I���I��-D4+���m��6K#;X�[���l�_&Ĥ��P[ş�j̤Z�����>���.FІ��lω�^���&kZ+]I%�@k�&M��!H�q�N��zî���X�E&Ӝ9`��{�83Tt�Ķ�צ��H���6��3��.5l2��F��ݺ�|U�ؓ[�ڌ�.%�h���m~98+��s#﯁�r��m��́��[+[J�� ���ۗk5�#!sN��3M�kB�$��Kd^�1j�a��}0�0��F�m�E�K]�X�����R���݈�'4�;�k���d
�XU)R�r��sÁY��_
��Z<�i�<�G�&qt_[ �ˏ����q�e���n�AW�8���fb�K�ɛ�����+[�)'W���+b1���+%�4�7q(�!��d�xn�/P'y��FCS~�Ӻ��$�	�uj]�ݎ����H̭�G�b�V��l�/h�^y+�)�R�Jj{|B���w��	�gk�� j�-�n]�M�*oXEi<V�;! {�F$.F_�7����t>e*p#� r���7:��,O�S������@4r�d�M7$A	�j�H�z�C�|���\N�;�'���?e������:��HD��D�K<1I�#�_����FĖ�dD5A����� ;���.��������a�����,��ѣ�'�A�����}sJ�ĝ�@�js�Am�b����\z�m���74��I��X��['`c�h$(��Iq�`I͉	�XnC�i3�;���3�@�l*:�0�Y�Ʉÿ�,����[��Z�"f�6�ӡEe!	��F�� @���$��6��0�=�'�/�_4d�T��Y��1������'vyn�m7�َw�]��~�8u�j�\��u�])u���ЯM�W�/*�|�iz̾hM�u�v�����Z��qݰ[BK!q\2�(�ׄų��-_�Ǒ��7�G��c9	�e�Cx�b���D�U�L��hw�Bɺ$��QN�J��ԚG��˗HG-M�>I*H�'�B|���o]��D~5��5���	���O�T�)r*mcZ����2�B��p��٨OH��Ɂ�P�ѡʳb����PZj{Bʊ�����Gղ��0�D�Oy&S`#CD�����q9f�i���Jc���(N�������):�3�%���tѻ�⯅�q �;��b7���,��^U��A\������~פ�/1�v�}�?D��>��'Ff��3>V+>7�얎�������Ԧ���&�����q���N�V���d6����;���xi���wWe��O�R�&l.��=I��ה���fk�A�)8p8yÄ
!�� �oE����~�p�� Ђ��Z���Ŗ�G�������,_O���v�E&�_�ݩ���L-8r�h��B.X�!��LG*	n�b,�#���Ň�:WjV\O7n���\ur��f<ƬU�B�q+��Y���OmOOB���D����œ�B�9ʍ0-w��n=���p$���C6�r�ZM�y_�:<83Y	X�D��_Cu{w�PZM�H+�u�����KC�7L���i>&ef�Kpdѕ�m�mk �2"��r�ǔ)��*�{J�H��W�X�a)�'sO��#q����<C�-C"�,�	��v�`.�h�vc�7�Tt4:���?2�n8ao���f%{�L��o��&(@Ox�¸�u>�"����"�z�o�|]^�ƭ�Hp\��]�<&V^ۙ���c6�M��?�C%|;r��	��z2�ߡ��ُ�7|߉]$�c�S���"&2.C����
��~��,��K�l���*� `N��QA�D�L\J`ԒnD�X�b��A't�$ۢ4�eg�~9s�o'����{\���9�n{��^2`�?��B�-n$1\��{ç���Dp�lf��KGy��r�_L�
W,k���_�Gb�p�~a�Z�=C;,ڀ�PGc<�VӅ��W����Νx i?�{Z%���l7�w�����%j3mg��ր���l���p~��:JX����`*R[Ϧ��O4����i�����Z���2��x"Ct�tk��%�����A�#_�*���_� �@�	�����Y����4��p�Z�Y(����:��h	:�O E��?��W�uk��~Q�7�S�����+Ԅ��v*K��)�x�kcF�(3��8ē��D����s��C�0��ݤ���<���I�@�`�z�6w���^.���-�>�%�bqC�s�y��vbFo�G��2��|��j��9L�E���g*�k���#�'*-/J$^2���x� 5��󌥚��K��/�n���(K�+ٌ~��p!"��8�
�i�'�'B�B�Z3����v���-��q��E;�5t�pM/��|&3X�5�=�-�ڬ%(t�k#T�	�����������7+2,���3�E��nDa+�4L����<C�{R��0���kB�m�����J�\���F�7�^�N�h^�Σ� U_F�&��6�I���D�	�'8��jz|ѯ��c%j������a�,��`V� M�v��:��Y믙�H.B�B*4r�ry $��r<�rk���*��R��P��G���~��4�3�T� 4�>�z-پ�^bf����7Fv`�2*%�E	M: ��������^t�DA'���R7By�1ih4�,@v�2�"�{��,����Kh�}~�a�J�\����5[���	ӆ�l���,09(�F��Il�Fң�Kb�+lLX�Z�T�"4�v�G���ey�:>�)2`�U���T��!��;�ӿ� ��F�����+ ���$��j
��*��R,o���K�k���P�e��sl\�_ѿ���*�o�ٖ����U]{�t��}5Bf���$�G$�(��y������i����1'c">3��2Əc�J�������෍� �9�ܢe������ M��@{��;ux�$7Yx@���6�)T�Eb�ƨt��~�~#�=��}�D�;���0� �A�E�՚���@9M��>��S���;X'�/JXa�LO���Ƴ����L��:l��~W³Uwi�rF�+�4㧉۟)����^~���y�TI����aW��#��k�;�:_���I��Sm�����͜�O�ro�Ydr�79w�J��&ܞ��7�7�q5P��֊.�?��w��o�N��x�3���QoM=u&��uY����b���M�-lcJ���_%�(a�>5�d�u'�tUO��9�7_�;M"���/M,�c��@Aם���-qox�?��j��He�'��B�h�k.�� �p��X�e!��E�׺! �Zȫ��/�t��S��-^� �(B͉$�Y�\���������fft��~�q��+�v��ѝЀ��@��f���kEm��E��f�E��Y(eɶn�;*�����+ 3�}�����]��������\�QKP&΀{��g���s�f�'��#�'�'�NV�@����&W�;ܐ�E�/ʞ��xLz� �tT��=!�\�Fi�NW����e�!�Nz�5������� �NҐ�h�y��Lmmp��֡c\kR���77�|�B���+����}�0��H)+�r���a[.�S�2���+҂j�-`z�*�~�h�j	���@�ך�O6;h����Ш��ᶧ���g,����>���ǜT<�\d�fL}|5c��$ҭ�����k�g�>�Vat]s\G.�����fPJ�s��\�P�4��[�0�x�ث2cP<6�:ｐaJ���o �ٍ"
[(c )U'�,�^_�O��� ~���N�-M$�� �:|�ֆw �~��1�U�4:��w�-�j'^=�N�ؤ�����'��W�� �Z|���I-����-�*��N����UW=
�=�&lB+N��͡�I0�r�iU�����h�7�!�ۋ$|')��dK8�n�=^��i퇧�N�1�r���>���5�ˠ��3@�oBt	ޥ�dF
��h�C�Sm�đ�bڽB�xfKG̾�,}1k��{�A��(�\�v��Ä����1GLoL~�����c��۽�~L�g��[�&k&v�G��V���.�s
a�X�jX��lp���t|����~�/�c��]�j{���ʺY M1����/��n�������ѾC9
GH$��c!.�M��6��?�}\���N�-��^�)y�	�4Ӿb���qE�{�M�}�.P��˱L)���ބE�����;\�φ�0B�} Z�{�;]1�E0�Ү�&2ձ�!�(*ҹQ�f��8�dMzbڼ�	�)��=��˵�s�k��w�U��6��x6�w艽)$��H�V�(�I�u��i�h%V	/7L4:��j�/�ܶ�Y���@�H	�עu��\��ڔ�+�Hs�ζ"X��O����r9��B����]��bȦ@@������7��� ��kΊ�DȄ�]�sa���:�k����3�H��r0*�b_
&MG/�]�-��d)2���X5�`�����-�)�Y��V��Ǵ�5�K�"!��a EgUe;䆱�}k�M��-%'&Ե���o
��G�jȜWZUK/�o� j�.�������+�(�$=gx[�T"�׼����c��D{�?W��{G����S7�����N��O��ţ�$d}Ek����(�����*����|��j(�c����h=`V9��!Q�'6���t7NK�_��:��P�ӚRb���J��&W��
,1T۱�3T��?ݙ�'���g@�./8��#~p��!�*�*ڈ.�5QAɬ��*��v�C��v����@̎�Yݩ��C#i��)�oWU�h�@)�V�?
��v�ﾴ�V�5��[���+��s�w:�����6#i��q*w���� 0�i�t�7N�W�r.Â|�'��_鴓�_|e�S0�q�j��p��%4�*n]P
B�Ȫ���N7�"o=��euc�6��5���x�Y���݄EB`���m9{��++�vr�i{�wh��������	�ٔa�q���xH�������_ăs զs���x�Kl��|��<��E�j ��)c��`х���;�E���U�=<u��䠁x:}z���'���lM�P�O\<�J}+wYlX���f' � B��Q��9�f��GxM��B��)�g�%� {b������j�]��m�����+dzo{�ZѦq��	h��X垊�ث�\�S��֕�y��G$�y�d�jihg}PZbc\��r&���?qܻ���2�E�$,�T��͕Ώga�0��gEl���;����9�~���̊RTz�lf��~��lp='m� ��5�E��-���Y�>V�3+�^B8�^��_��9�3�3�K�L�r�$aRɢ,����
f��*l���a�Z�����q�������0��S����i9ܧapyD��lj��W��A�z�Ю@0���;d��5k?}BE�!����<zL�O+�e��=T�64
;�v+K������D�>����M�hO�e���=�r!G�dQ:�& �yi�8E95xVD�f=ӑ=��M�)ڦ�k�]Vʚ�Xr�bW��_��{�o�(<��?���8z7�q=D�pN���N�5h���Q�z�j�K<��ʒ���
��D1�M��
(�8��a��Đ��`�h0(��-��)أ%���`E�y�N $p̙��+�<�J� _<詘��Ք��GQ��2�����5���Ϛ+�� Y�n��z��S=������}eΡ��bݮp��@��h��1(��EY'Mc��Ǯ>���/e�= %���+�9���qv٣�˫K@��%O�֚h���%���\��Y�!N�6\��R��c�IV���V��Ɂ^�IհnsI��U-�3`9�u�h�W>&�(fh�8���<q���N�C��L4�V$�V����j��ʟ=�r)/S!�g���%�#�o`�/{��c�>�-A��{Zߦ�}m�1�v �"�d�_߳�/��6{���~l.����Wt
_Z)f�N��l��Me��mւ �|/氦�$�իՒ3Z陱�^�7k��F��R5p࿕�*u��xI�P��e�)^�R�m�D���t�{~6B��L;�U����0�Li	���j.�Hl�b��ʥ�$O����;#�� �p�������5�D�֡����U�@��������O�^��M(�R���<8Vd���7|������#B  �޺��-RU���E����ʴ#��5�z��'9�s��^]�6$�ޓo��9���6��9���܃7���e]lxBj��{�5x�5�lQ�^��|�h���Ȭ�,1i�@�Av���Eg�>�E�e���� SʹJ��-%<�E�u���������D��d4{;��7������q-��h���J	�Ht�'�8�=Ha��Vh��T��y#E�̀�,��D�/ě��`�皿X�˹�0�����R`:	�@= �I]�>#-rQ5��=�C��
�D�(;�E�����W�'6�!) we�*�P��5�)�����|`P���� ���6�#	!u�,Q��09�Ɠj�X�z*���4�7��r_r��^�rTv:K�u���No�D��89jʏu��7܃{�*���ίr/�iP["��7���z}x/G+��!@4rQ���o'�
�ȵ��՗�#ŹX��h�`�P�3��vj���	?;xw�x-��g뾼�M}l\�#&���?ҏ��j�H"+�OK�`P�tAL��k��y������;��8�dBk�-��K&���N)���~J4���9SӲ�S7����Yإ�0����;�E��}*OE3�4���X{��f-)e�}�f�p��F��
u�am���)��'��I(T�q���x�Q�6�W���0	7ֵ�%	��2���gL8��ߨ�ɝ>?h;�Tu*��5�n% ��K\����۹�t���VC'�+Ơ1٘�n0�E�� ��k<���.<���zK�˄�	J�4������R�d͉A�
<�]�-�=�%���"�6�z`An��t�_���y+���B�Jm��_�T-��"�+$��{=�����ƀG����CƯ}�[?h�_'�zS�&	5�2����gof��]
;�/W�P�;w�,�˦mJ|� =�;zQ�_(1�|�r�veP�S)s๡wu�(9��E�ΨG(5�;��8yl�'��CZ�vلq�.�Ճh���\��xXr�m���Q�K��~�1{ݍʙ!����ӆW�Ο�co���5��A�����-O�?ށEf�.���n t��F�ϧ7}f�C��3�견���ݾd��|�QH�����\ϲ�X.�.x�{S�4���<�1��4������Duןu�U��C����f$��}M��g"��]��Sjϻ���9:ό�����1gS\�/�����0e��g =�����D��g�+�E|�j0�2��.�
{�ߍ�/kja$\�3YqI
�R�S`������,	� "��7���"���G��ow�w_�ոp�LV\����E��(bA�F���v䉷�?CtK�n�"�7���ia��3É�-��T��x���I��*��l�ba��y�F:��T��)�po��ue����C�������sM�s7B�����J�]?b.��;Fm��Xun�PG�"/�!r�S�hB�~�n:��Ѝ�`uԉ�{Q�%E1�i�gVn^�{���ݍ�J��Ӝ��k򄯒&E:�+c5��go��#�)�!~���3ݦH���..���ܓ��_�	����KH]%��'�6BL�-���C՛(}��hm��J�r���y����(7"*�dY�����N�:�� ���囬�����̺��卑juD>����U�n�ԉ5-���]5o��o|R��R��Q�+�@A���\*�`Q�
d���>�JdD����ڦ�P�r�/�7�`^����� �WP?�� ��ۀ�i�︫���]�fT	
��5�_��;\Ԋdpמ%�cc�?f	�;�B���m���^��w���L�F�(#�ג�w�)�s�������=n+O؎�ͱ��3�݇�I�̫NU��&��n�)88_	����Pf棠$�+��}&��	b��)�M��^�p`���i�ܸ���9�(��cp{.1eůr���N�`��A8E����A��b�4��H���P����IX~lu�صp��jִ�ab�rO�����e�O\�X�/�J�^����I��x�
 �mst2TSHa��2�΃�]�)�mt9�M�
2;���Qa��.@Z��{�Krn9����0�~�c��n֡ �A@й6?�p�f��y�3Z��.��-v6v` ���*�5�O��� �,pڇ`Ƈ��$]�4l����׊G�����*��m�| ����ʱ�^2BR� �4��Q�B*���I��b�?��'��IF=7P$}�(�N��K�%��*�G���$-0��RdP����f�aAߛ��I���i��Rb�Kω$74GYc�
 JV@���"�u�_,P��S{�D��UT�+��	Y�3pv���y�,�+���I�j��v�o8GǴ��Bǆ�v�$_O�v��'�'����d�X�EkEE(I��@���+B?�MD+��p�PB�A�����5�M��L�Z�=ӥ5B+�DK�#E?�x���'��,������ދ�Cs��Z�I��Sp�s�� T0^�����C�cW���3�%�C��ZE�(?�g,���I]��Ȯ`�ʓ�ﲜĞ����#y�0��j�"-�r��u_���-|"b���/S���@~I����q�{�(;��=iB�|1>
c�I|c��[�߳;
�KØN/���u���V,�ϔ��}cku������.H�-�Ƃi~"����
Ϲ�C0�7�j%� %�
�;�Vrr8����Rd�xkwz�ĺ��h�nٓ����U	�
U�~���S��<~�Ơ3��F��k�F��k��������uE�,5~�u��=t�ܸ��[c�7�޼o65����`<۝gfhr�����6��ig�<�Q�Ul�fH��<H�E��)�4*t	l]퀡�g�&����LoZ�җ�K�B�=k���!⡱Gu��d�>�I���j�lsonɫ�8`܃B�ٷJ��{�0�w{CfV��g+5-�ts� S��|������gc��A��	�����eh�,m��vo4jd�,�G4�A�-��#�	�r=k�ET=%�j��A�}0��V3wjX$Cm�G�>�F���v0<�b��g����vx6ۮQ�ڵh
�������G�Y�И���&xE��Q:@"C�5Q@��ǈ���*��731G��v��`(˶��~��xl,[R5�xq>��Bv���l����!�����~h�|AA�B��y���!d�t��+G��x��ɚ[x��^����a(Y9���ە��h���|�+�������$�\�������[)����c[�?m$B�i���P�r�:vm�}��#��e�c��*H�K��P޸pyP߅_Y���~��[�l�7�u�]����@X�H�O�� pE��ک���{�L�P��Ssh!-���4�f�D70xRȐ������ѧgT9�Ω��w|�՚�:T�����x�u{�e ��Hv�М�%mtM
�y��3�i���QY�(��WÉ���_8�nG�qP�$T?X��΍<t9��r�ƣ8��BB,F~̼ݮF��o��C�o�eDR�ԯ�1�oh����P�Ů9２�ĂD���#Xz����X�-C�i�a��+k��ד�Lԗ4� �_y�J���ц��V?�W��>C�#�J �қ��aSX���+m�� �2���,��.+�����5N�0����p��u���5���Ҝ�x�e�N=��v�Hy���b�Y!t��M)3�)t�q��FXT`�"-�� �2u���f6��X�q�RQ�P���c���}�y?_��E}.�G,���[]�
��5�bqVFe#eT��^|$JV.��|1�@�Ũ��l�"�5t���7�}�����;��.�ݵ���n&���J�e&J�L�B�d�vd=��5�WZ�Φ�Uև.dǽ%h�������¾����f�I��Jmκ�Z��?1zi�jֿ�r-#�vsL��\���>��Z�c���(�C��%˙g@ˉ��V'���'C�N��Ю����P����⧧��q���;kR�X*��l�+����ˀ(��G\��O����z�'��<3�"��/��.�.��XQ,��߭���������c"�����e͠��9�#H��y��x�!�l��)	I~Q�����28����^H�mU�K�r�1�z}Ѽn�FC�ωo���X0������ڕ�ee�)e:w��:Png�x��@��;)y�ի+��V�'Djɿ�����_ ���~�?Ra��äp?
��ϋki]������ٵ�ABX7�rG�T�91�[a_�E6�5����i�b9�9��&��0���B�Q#�	�HM|��I����I��N9��d���F/�(�����텰^Q���rP�`R�D(s��ݱ����֠��NV��P��
���`N��V?/�,�X\i#RVg��}謑y6D�z��U4�m�i���5���hA��>U�|�n�ps�Ik�Q*56���U�(P�6���?pG���*�gH�� fuS7�@�3����e�/",%� :Zk�O~6C����E�nh���X����HgV���@R����ק��z�M��I�襚s��h�M�}������t��&��m߁�����:<�m��v�ןip�hz@q������Qa�6A]�k�^�'ğ�Y{�U;�̊�'Β���,�d��y�Z��HBd]��Jx S���v�'PnЮC�B��F���CC�In*4&,�xT�n��L^2�d�*2�]؇��j�"S��x��S�t1��[{��43�(��S1�JL��6�ݿ�CQԛ�ý�6�Tli[1�*ĲHZ��S����.Z�5��_:�	V->.���_�Y�O�H�|БB"��O�⡼���a5o���>X�f�ݣO�Y���L��v�������z�g�׀g�j�J�!i��"�-�Ib֒^�J7�B��z�1�����c�_�CiNJm?���1�Іy��շ{�`�uD\��Q�cѱJ�K)9惯�q?��<��;�*�#��F�U�t{�sEM�L�-1S�=�����j#$h�Ĝto�w��HyyA!�>��L�
E<��εд�~�x�����H�9�ɸ�..u�/ ��|F�+�wV�P���'T��[�bq �<�.�ɤ�� �� ۱μs��{P�1gVƽ��B�o{1s�_�;�n?��@��e}��~����q �d�9q���?�2��p���K����fKe*땉�6de~
K��z�?E;���L�`��Z%�~@�Mg?��?��΋�1���Q�{4}�nzXn����bGը��	�S�-�6���\�璚G�M���_zD��x��#]�k���(R[�w�%�C=W�yw8Ŋ�?�K���6�P�>�aE�0v���lP�
L�~�#���zH�С	��	�!'动;	B$�ݠR�+v�fU���#:+_�>�~���}���-���_�ۈ��t���0g���%�^���R��-�a�xr��������
j�/i�	k�q�
��\��S�,��Os~X�Z	�-��/cӠ;ye�DѾFt4��Vx��&����$��l'�&-z�#�1,���z�k'�I�?�I��D�v���b{�cV��0d�.���Ŗi�D��S�O��8�b�3A-�NӢ��,��1�?K��g\�6o: ������M��	��
�╡�=p�g�d���g��
�,�\��@o?�!,#�~:'����іj�艒���H{�>ȲG9R�v;+t�b���_��K���m���m��q��-��(x������c��m��2;&� $��?
��LM��ُj�σB^��&��A�k_��4���:��{0���a�$
}��-o��L��2��1�������'�� }���W�h��[3`��N�jR�|�� ����<ټ]�TWӈR��!��	+[k����fIm)���},F�N�+3��{��2k������ҋ���Z�;\���
��-(U��*��эh^�#�L�|Uf���$P`:�p������A�]y3�����@x�����)���Q!�aVN;QC��Nɦ  ��n7��.sUo��;-��*�Š���Q���6�+KB�{�pۺ��3X����G��<�ڒ�(S�^ՋA�e�8W�J8�S������܂A
���ק~�]�ʽ�ɭ]0Eb{��0/Xӱ's����Yt�]��pA�x��$����(�:;���=g��c�qr ˯1��i��E���i�n��g�z%ۇ���R�l��]r�x��Bާm7�mZ�O�˒Ot��{�m����(D�T����4L��(��T�f�$�}��_w�t��1�������88\�h���Q�/�#lMyL�Y�R~0�ֲ�_��I�ٔ◙�l�>���	�j��hߖ`Q�|pm�۔�p_�>�!»��.2iE�܌Ez��f���R�R�I��������B�\��%:^��6N���:��4=�����ҭ"����9�B���Fj��Q�6��	M���Յ���Ng\c=�� ��pu6�_���q)|"X٬Kq����c ��mP��D33��ș 4�Y﯂�7}��+��q��mτ��T�d��K�&r�ZLƞ�{x�V��6�<>���h����Q�{~��
�Y��v��ڃ����OvID�}���-���7H hL+- ���/����zvg.'�|bb����������a��DQ�����p���M�D
�Wé̛~��0K����K��1��5ed\Ofa�2��Wͭ!Oi�+�q���іS1�����/�����zn�1�4���<��;Q7��
N�~�Oi��?�օN����`:�!џ>û��^G�������B�)�@Lo'#o����u�X�&�Q�m�w����>0��4�Y��ѕ�W@<������E��U�W!�r��ؗ8uTj/{2�G2�t��Y��[��¡R��/_u�R�!�'�Ibl�T`mEf���ɾ�r�����Ww��k5.k�N���g���n3����ޥKj�bI��f�#�c�yVB��9|e���E�s����:,E(���N��Y ѽQ���u���1% �/��x�9���*׹��L���Lr~�
�B�~Țb��ߤr���e�q���Uh�p�4��I����B�su����ƮA��zŘ#��
H�	(��M���X�������H{@1z��t>�����H���y��!!��wy��W ��H��i���.i^g>����H=(m�嗷I0� ��,M�I�}4=�ek|����Hy�_O�_zV.�Ѫ���n�}k3�$ ���X�ġ����v1�,�C�>�������qO�r����'�(3&~қ�R�B$�*��0���	���v�8�����AHUnU�݅�q����6_~�	�xZ��E7w��X&���_䲿�ҍ�!�5;�WT*�j����������c&��7J�s��C�	����W��vq4�eagjq�E���4�׃t��I�"-p ݈e �(IÏ�L�05G������ut��k��D�}�H���n����K��n�l�Сz�2�������e�&4�'\�L�V�����G�N4��QämP�Z����d����UJ���t�[6z��|�a&����a�Ӈ�3)�i���ٿ`���,���J��l�Y{���kG':\l[��c�\��r|��p���h�j ��tUF�CU1��7g��C���fٌ\�粑\�<#+��������:����<��J��K�;v:�9�*�G�!+��;a!�c`��aK^�5s�[1sV��~���_�CVa��~|ᛳ��_��C@�d�j~��F����"�F�i`8ٷ�;_c)'���]�I5N�YGm`Iyҕ	�F?��cd�P������uÜX=�ui.03���'w^XW��	rJ>R���j^m�
��\	�}��anե~4�zr=ht\ۚb]�u&%��a��� #^l��صa-q�T�A�.Rf�O��n��CI�^�D&c�T��Y�@�t�|#��p1��<�a��Qd��x����H�haI8]������ff���&�TW��-�g��4�.�[�v>����������o4���,O�4�U�O0�i�/y�l���@ϲ3g*�
+.���0KF��3Ld�z`OoH_E�E�$N����a�������o6/��9&�*���3�����@-��둗�	"=�"���/��?OQ�<�L�ԧ��-��t�p��qTe�`]V|���LCQpUB%�vi۩�O���㡲^�di]�^jm9p��K�	Z�(
צ� 3��$x=�;>o�G�Xp.87�߫UIL���Ռ��t�[U�!a`2'}��M�P���� m��_�5$�;z?�^�������	��P��:���7Y�ȿ1'!oxd?�c�I�K����W8�����Y9T,�=6�p�4,�A�r�c6k�ܳ+j�ʋ��i�p߈^i#b]&�쐄�)1�d��ZWɿ�wh�Yv<+�v����k�5l�2� =^銷�J93���N� z����F::�c:�
�#�N�\�"�jLl�L�L�obG����6�>33�?.׀~2�I�3��s�.~��8�M��6��Ffg��<��\�Qf����iw*T�=�5B���JvY'@�d`Ixːg�C��ɭ
��Ό�87�Q�bd��-�pQRk2!L���x�Q��/:�@�DM�>��A��S��,p�WC��F>N��̳X�2���:���`�8�S�G'�������iI�jW�J���0j�[[��7�-�W�[�bg<���c�E��~�XmXaM�>_��'��1��\��m2;l�͊/|�N�!q�(�����Ly�6��$E���	5���=�am�uk���#WE���C8���K �=�,�n�G���{tUέ�^�����<��%͂�l�Z��<ۓy�& ��S}^9q���z�p�`T��	0��;�B�>�B��9��y����ӛ3X̹AZN�U�j� 篎�`����{z���Fk=�H�3hԢ��d~Ь��lKdk�8��x��w�ME�+@R]�_HS��و��qc���������(��%N�k� H�*�2�X�eq�F���a:#�
������p�h�hP^e�ZC>*`��?��e�/-,������:���1)O�Ч9�~�HG�+m�п�߳ϟt�u
R�Q6�����s��9��z��u�����3z3���ds��!���o�WV<B���!	��̔D��2',�3<}�E�a�i�V5�J�Uz'P�(27�K#�`�"�)	].$�ޥ��iH��.�G�gk)n�4={-D-خ�E�eJ;y~�͢;��Gg���t����z�_���j�65+���C��n��A��&�Q��$"w�w*��7@����~������!�9-����a�z���*���\�#�X+�4��2Sl��,�P�����:qt���e*m�r��&�㹻�Ϻ�� t������%��Kr�c�t8�l:��&��j�q\[�V7j��R�`d�i5�%c�;�G���)���n�(��=2��p�Ѫ��{p$���=�n0s��� �Y蓺�_7�E6M�Jlg8����C>\����z��ۗ0M2��x�A?G쯤۾|e����[�)$�$#Ĉ}Rc�W��2t�;�|����[&�soI2(��C?�4�&���fZ�J+����8����"3W�־G*��8����Y�!a���"�B��x�Y�,:,��x6mְk��10m����� �>+ ����dV�#��n��!$x��{�A�3���]}������&,$���z���Tȼ�V��L�(Z��B�-�3�\ogeф�i�4jV|o{�w�����8��o��فc�G�����x5N��	v�Ym(R�m��bTHMн8I��Pږ�T
�Dv�Γ�E���'�c����(o�8��$h��A��	9Wr��S���9�MuLh.�0�)�_�6��e�n9�^���,g�4WTmL��0���^�[�Fe|ϭ��@ԓ����pM�
=A`�^�L|��YǦ'a����vC�ĞrFEPƞ�JD �7��U|2Yv��ϯ�0�R�AjA^�]�:�����x�(����b��.�~(�>Lsg�K~����Q�
Zg�:�fC\&�U�WS}�f�[��q�V`�?Z���9����X����S拁��W�n�6����Ǜ[8�sIs&���D�x�D״�(�'���N_FC�[��V�K�oY�$E@KN���>�zp���u�!K*�v��F���U9�C�@�O�4B_
�,�h�/��>����bX�K�gg C�k��!�<��6!Um���B��c��D_���I&+�q�]3��ܓD!�L�pj��x��ư����hHq��
=���;@_�G��vGPޑ��V�jĊw�`�
_f�?՚b�z&T�3����MN��E�d��ws��7BL?�.&�_6z�<D"�s�KØ䟡�rP3N�ȯ.��hH�`�����уX������"� �G-�.��2�G1�t�Q�`M��������A�3��B3��X����J���LE�<��BT��i��XՊ~�p�n �$��J����|��k��]ֹ�RoV¥�F.��ܥ,dN����-���@��¨0�©�]��M���k��s@��$����s\$���������i�i�wS[�v�}��X�ry~R���o�NLq� �Qk��5`�#gVi~�n��;�B3���z˅_�I�뚸',u�(c��ɐ�'��9���QJ�Js,���^��@�S� �5P������&��i�u���C۞
*��eӋt��`^/`T�f�s�Ƞ���������唟)�W����w��j�%�O;T�;� ����re֍婘���3 :��&K�ut�����8fcB�V���=Se�N����:3<]��ō�裟�VcE�\��g���G���vɀ_����~�ܾb�_���o���"���ԟ��4������Am�͔Sw�=�A��m0ЗuL�8~�*�6�"g�j��P�R��4�G�Arib�?�`hG6ȷ	����ww�����a-c*��'\iL�܁���%D�ki�I��O�4Ew肓��V:��e&�5¡D2Hų�K�f�s��y,)��}���t�ޣ+�������T��{|I��S
�"�&i��nd�޽�3�G�C�_~z�[EP��CP3��>�."}����Zʔ��N�im���������i�]�6�%d����K.ё��O���o��f�jΉ���G��-RԽ�8��'�J�XР��DB�5�������Xp�B�@�w͎,&�h; &��B|�L��"�� ����Bڥ�xqiW�CZ|�s�n�� ����AA��C�ӭtL���p�i��8����|g���#'�Mo���Lk'8�,>@I �GgR%�k�T�4�wQ&\��j�2Dj>��`[UH]�Y� �%���K��Sh�n�oRs�G�m�fn�c��;ܩ\	�~	2DoO�Nނ�>%x	�&�-[�/��؂�G1�Չ�P�� ��Mk|e4|�T[r�����vaI�:��e��U���riBO��O�0L�
�����;z�`��sT����y#���b�����ٛ��	�$� ,�8���#�Eb�|g�&Zi���<M�}֔�$�G�
�d�n/�jd'�(�T�'p	g�̴�x��5�/6)c�h0I�7I�b���~�dݣ�\���]����������O�)�������j��<�G�^�ɩ��o�c��~e� ���. ،%ƒ��ۋ��7���b�������b7�7b]//T=��b��(����Zz';�X��y��̭���(�f�12������ʲ�!��㒹>\F����}�^3Q`���� И��TB��+�%!����NEl24�.0O�C۶3��53�p^���T��|Pib�� �4��W?K�lbq��40y�c�Kp�s����p�S)<�~��r���|�w�����s�T�H{�	p�Ԣhy����9����V[��eH���5 �s�}����8���\�r�q���;L��5�C�V
b�G�C#�B�/!M�D��.]����� ��&V�~~]��p���e�K'%���X2y�E�r�؟�X��+�t�����}<O�G[��G���ǧ�"�f� �]DD��F+�������Z�d  =>C��f�>�����&�ck2�dm�09��(����o�K��>�^�	������Ч����b�i�=��$��]�UA�Ǔ�A��D*%ޓNn��io��N��ܒ�vdf	Qm�����?- �K�;A�l���#?�K;���?���Ǭ��9�?��k+�|cA2����%�mE��]����5��g0
�~N�A�!'�������Yv�p�Y�G\v=G��1��-dP�$4�?A���t��U+���;�9�Y2�U�7�Au�[�X'4�m@�Q��kTC+�F�(��{���Wڴ�[�sqB)�#&e�1�FL�,n�PS9��cFi�-a|���z���xtͻ
Z8Y�:k�J�,�Y�}qŁ�5��O�s�85[SjE��g�`�o�>��������vt��3A!
�Q� 2B�cAY��ڎ)���!D@�.�>q3 f�F��J���b�(~N*C��t�u���q$[��7t (��}��(���|^���'R��y�i���Z�
�(���I�[��X[�$���]���Q��E�[c)�JfW8�&�DS�E_���7�Rĵ]6u�Q498dN����A���<��Bi9Z.�x��>��|i �D�E�Y(~�����z�����R)t)r���.��<�6�ћ;#�>5DO�)�EQ�3|�����oG�vH+f2��*��5��)�n�e!���[���d�O����x��&Vx�&Z���'?��oj��4��~��՜:'j�"��,NY��)���e�$�93�"���d�π�h7�Ti8k9`H[):��"��g�
D�J>�
�� qZŌE�ow�@|�(P+4�LL}��i�aLUL&,����Q�Ar9�;��5;��V��<�F=��p?��3�0�_�)�����o���o,o�����[=����&S��A�}oEXJ�[�Iji�$ `c}�s������9i�[�L��\7U��8��H 2��1YZ��~�������
�A�X���;���@���e b#jJ��d�=N.�51񡶒�oDl�<T�f�uD�J�^�]��`�V`0��º-1~�+T	�ve��s$�����}��+a�#���Q�*�^�X���k���#V��G�;u'���Lim݃0H[�|\Bk��77x�V� ��E�>B�Q���e�>��=�4T���tC����Tϳ|k���t�.�H�ʔ+)���M�W�l�NV"�wj�tԥ�c�^X;��v�jP���ʒa���қ���N��B���
^�K�#*Vs��?(�ك�f���|�@]&���kw�o���L��S������5�/st�L�tp�Y�<���� �� �������jK�7�7��SDY���M�&�O��R5��I�����uQ� }4ø�?�{i�.$������N����L�+q�w����_�Y$	�x	�@ąZ���a�FNL�-��J!�2��F!R�)��VZ���m(2�psX]�^Y�y$·������{���q����gJ�p-�S�¶����Y�Opz��b�c��-��f,ϬGoe�β�_7O��[��nb�v�����Ж�)��h���~`m�q�`���{�V�b��9��QX��jձ2F����c�Oʊ�7��Z{��"y��++�G�˨^�����$|+ZS�"�3�c� �e� ?��oI��3������N@~P��M����ڒ6K8�z[��)���Fݲ��n&�}r��u�.i�2�w/��[�y�Te��*���}���VD�g�¥P{N����:1O�p6tމ���8����>ܯ#P>���L*��hB���|C�.��y�'Ti�ǚ����|Z�b���?H���A3l�y5�g�� �P�Ԇ�ftm��<:'r{�Ɛ����F-@��:SlMc�����^c:���`�&+�o慣"=ow���3VTR�4��㘯���Eli}�{T��}�u�֬r���& ƺ%�p�O� D�W,1e$p-��g5*���q�9,x�z�aɹЂ�:��e�����3x�Z�Z��7'8?r�<��G2��X�^��h�"�ۿ����;j1�pq�K��ڿ�@��N����%�+e���.N����Y��n�PMu��LBt���@ڬcl1�b Ͳ*Q�8������g���B�ƍ�}漢)xA�Z��Qi��2���Cs���$��*
�+g�� 99a�=�(2���$��:~Q}��R�8.5f�f�Y�
>m�v~>g@�<������q��b�o��G�����ۅ��
�Z`\5` ��;ȌÞ* ���}#��=���K!�h�^s�v'�S�[��/M��ʅ.g#�C��:#4�˘�A�M=k*�u�?/��-��������Y��g8C���+��	=���V��įӶ�"�bp����k�I�����vm�9�(�/�:G���.s�޼F`�2�[᳚ޱ�� �sc��k�QB��q�EJ�&�/<�N�O��2����1�*�}@f��Qޙ:e��smQXbE�U����oaM�_�b��k8�A��c�E��ISG6zZG�����-E���nV��7CRdU�?����"��د�E�x}�ĉ�ʌ�!�Qގo�0"�4����^�e�������n:d��"e��Z�ha���	�JY��G�=��=i��]e�"$r4�S��(�J���<��F�M�S4�&��tK���xi(`��6�*&��n(LU&ɿ�B~�qoH�zf�Qu��	d���n=ЋI�q�&@��*�5F��\G���H�0��+P;�꘽��i�E��<�:�,�uϘEèa���AM@�[���C^�HN�j�߅掚�s�C9�=��:N*�g3-��T�|���?�>���蛟~�X�����{fU3��BbW�-r�	���:��$��٢��D�vO�Q�UX�hT�!�9v�C��3�ρ򉍫��k �,�jȓ��yF1(�aO`/��~ZjN�x�jC����zN�C��3��f�̲H���i�r�����n�`�$�q���"z3;n0�R`h_�nߋ�	BHa����֑�d���qj�5T�e�9���(�;˷IT�F��Z��v@�c+A��s��.���o.E3���7��S]�!P<���f1�u �m]�iS�%�B��c������!�Q�H4���kq/����g��A?���5�|��)Pk�?�!.��O#e�9�l aF��F76�Jv�K�����_�����JJxHCxԯ�_R9;�}����C���_��Zҭ����)������ۍj*��;��<|�_[�~\,�����w*��N��6.���$vZđ8�&Ԧ���� ���(<�K��?�i�NWb�s��1u_�vMi���U�3��BR(b%�f�ۯ���`�-�GJ�=��T�r%���s��$%^oī��=�2�?���E:��[`H�*\$`r�ؑ�-�崺�)0a�:u���6��jR���l�i�]
׏:�h/�ƶ�?�M���W$9�+��p�;�v<����۵�t{�6�-�j�l�
�-p�����KZ���Jqx̟/}G�.��9+q�U%7�拎���/�lz�� �گ�l�H�(�F5ʂ��xu�E@��tX�d��*���3�[܆些1�?��\��;8�	���*N�ө��N�w��s�_����� ���Ϩ9Y�b�����[�)�r��FN�f����H���W�cm.*g�QZb~Hɀ�;�I��"��7+b���G����T��7�m����DB�0�Q&�L�A��Jȹ���;C�<}7Y�#�zRc�\=�~�(�/�QHB��/U�jP�6�;�"~������M���(ZZT��!��+v~���y��Df4�#�,Fo+{7��#�x�z˭'c��_�� pau�C�P2x���%���
��S�,ތ@5Εd(On3Xe�XGx!�
z��y�x�@�#��!\+O!p��#F�SG]�KX)�j��Ǣ^�"x�=��+Y���G�jL^�t8�O�G�[.xdKإ&EV؟�0<���:���]\�:Zvu�'��ˉ�d{ ��<���-�6��)��P6�7*q�wϸ����5$�nS�������p�l�.�G� �k`��9o�����K=NK~mn�_.$���}���B�ƽ(�}��Fo?-���+��,�G]}�ͩs4����M�/��ɶ�e�-2)|����:� �t,J`�屨̕Ip>A�x�}��o;z�ՙ�Y]?�̟���I]��Xb4�}�_թ���$W��6�B��ۭ�?E��D��,�"�<�9��?6�YOu#�޸!�rP��s���g:��4�B�������	��:P�q~*�W����d�r]4ݴ��5�w���)l'a�A-������R�O��N�A|"��iu"U�(��N�Hv��Hf��̝���(6�P�d����l`�mQ�>5է�$?�=����n%D���9�s$�QI�h*���d���Jpת��m�;�Ӥ�\����T�����ZN��-b]�'��M#^��3�m�G�S�V�w�~��Ë�GO�֝���M�ɋC �Z����(|~\�.�PٓY�!W+�M��qg�L5�-�	6�:�<Xd;�e]�mѵۖs!t�[d27��j����J�(|�2}���X�[t�4�K(z5�Q��]xΆ)�ߌA<��O��%��컞�bjLQ�\�B<�}������>�
�Ӣ-�+^_;h~�a��a��O�LvO���� $O�y0�PGN3���,���|0���$۰�Z��j�����x���D��ӕ�q���i�J���"��V�j�����!���2I��Y���G^.@�:���;0�<���<P�暺����4p�pc�,\�BuJ˼y
6���\q��+ e�+���?�9���f�8LJ:�Y��[j@Dm�C/��1�x@���ZB�2On���tH[��h�b�X��*��+�c {w
C�e�T�^��q��o�x�Y��R��B�����vBV<{Vs#�|uir㭨g�c鸞�fQ�B���VpD[9�O�Q4"sw�ׇ��X�+�U�P��=e�Y�[�&	�tn.y����&�F�L�����c��b֓O2!6�8	�ߪ�T�/2"�w�l����2`�f�8�R�V�.�n���_�bhfn048��_fUݬ|��ݯ<,SÂ$��,�4�.yMI/i/���^ߊE/5�Ҕ밞��Ư�l���;��	��%���U�F�>��؇B��>����\�6"�W�-q��|�p����o�ʮ������'`AP��'��5����c��6�0R�K����{2PD|po��3���W.���=��m�(�ٷ>�VD �}�	air�-:Mz��� '�z��[��}��ה�D�c����*mu9�����@t�,��qjk��~�g|���=}���1�+,$�č���\)���Jd�~�{E��xð�_��Lk���*XWP`�_zdV4��$,%R��[����L������L�p��!-�k� �5ș��")���o�6q�p�/T��-��gwRQG�{���̐6A�>j-e!&9�� ��ć	kl�U=K�A�)��7���{�S��h�}t�ZNsK��,��n4�F�M�����Z��fŕ�".�0���lIͲ�d��R���M X�0Ӟ@�fc$4�Ρ6��"��E ����y��L��RL�{�1���F��L�9�`9�i�=;dӫ_dJh�%y�Fڌ�h���ɧ�*���t)➪�x��]Z��(�N��Th-smۀ]E��q�8��b����: ����+�$QK��]��a�D����"��s�hl���tq�"�؃���|V�����:�H�q��@�JL@�H�zfa�E��ʄ��b8;>z�l5�Q/:������E���ܘ�TC�Y�(����
%ԘT>Ba���,E�b�*�q���LG'G���-��2w�>����K��i}��^��L�����t��;G�P��>�$�Qe``5w��4�d�z��ޝ�7�u�grJ����i��y#n�21�c� Z�5V�t2���;��3�D�I]����8D�N��R�<?jz�P�|���(�c�\��4�tJQ��1cuE}�(TY�GY|�ϕ����D��{8 �~�@�3\HV_ <�r����D"�|Y�O7 8�R,����J����[��;:'
���ÄZ���Z�`��O9��k�>k�t��3���H���>�S�
H�ʔ߅<���mS .NK`l�����V]��|�n�g���h����'�|��$����;*�g���= .i�r*�"\�RTʻw���W<w3a��!ݭO����R�}vf)B!���D�F+��]��,�Nn�����`x���[�]IyC�Zc����R�����!K!=5���̺������`QdC�h"�8��R�桚Ԑ�ǒ�¿��L8T�(ǃ�4����ؓ����գZ�	q6x��A���oZ�2ng� ���7C�ah�O"2x���q�	%r�д���*h�øa����ׅ≁�ӕ�\	�\�i�9�6=�[N�9�57��=TO�o��ŕv��U�B�SկKt)C�n'/S��@���:��97���r�A����C�sW3=#2��E�`��)��-��֐�$3���sM/1j�����}@���CA����b�:�J���Q`��P�����v���16#4c@Īl�k��6���Ҋ)��A��Ϸ �`5G=my[��۹�0��&�(t��پ�l��*�MH��a)�;C&s����nK'�T2�f���B� �܍����������{���Nx�p���P\� ����[�N���N�f��ͦ�n).М��-Z�_�шP�è�<Q�-�
"��t�f@�C�q�;]%.��z�U����B�[�^�	I �zs��j�ԩ�5(Jq��;�hy�������xb�j��%�oT�Ꮢ=�%�
J����о�2�U��DêC�
��S��p�]���۳��"v�"����^��ܠ�-�ʖ�ȴA5���9d7L�;�ad)��@J�W�+ ������R8��%g�ˑ O4d ��A��ә��<�G�N�U�S��*+#����, �p��e�n��L��7�}hS��@o5�֣�	��]�ᎧyV&�R�,��\δ����e��Okp^3���zZ(�e�����ou�,B���ɚd����2��^6�*���|$JO�+^<2e$>H-��2AJ���p16��y1��}�[8T§�9�V?��@��2!n����JIY���ë��!�eX���Ȗ�VO=B>�t����/�}��(#��w8]���)�S���y���.l�V�h����Lh�����@=��ٳ �Tyٚd���%�7$�z���+]9������YI�v�w���dl������B�|4�FzL�jn<��* � �.iB��I;�T|mn���9g�MI+�d/�1=���V�a��n>�U|�fj�	��|1���ؐX�;�$*U`L��Ɏ,�y��G����~1V�($V)��ˆ��9E�ǹ�����~z���Ƙ����rRT�o��o��hŤ.z����c_	���T��تB�q�K��S@���t�%��ޥ�T���|��,�8;���@'\a��Я �z�qhLL��),�r\@�8�v�1�e�C���7�&͏��/Z)\�Q
� 2�/��z��Zx5I����m�%���X�̬�ό��08�D"�ie�s�t��WI������'��U�@B̶��d��T!,/A/��y�PJ�-6�p1^�#@~{^]ʩr7j閏$tw�=��?|�9��0q8I�:d��7��)��-�f����'������J��{�T�������'�G�]�1-pF���{��2I%ݎ��B���L��Q��#l���K�R�T�� �(%�1Dk)�!��J�W��f�9����,Q5�o6[d68��L���B�
#)��
��pF��w�0�Nw��Q}Z��9� %$Y�Z���-U~�z<��0��N����r<G�*��^���$��vm��N-}C39m HF����4��W�d�W��4g���I�y�O�0���H�:��e$��Y!����},d�4�g	�k�u=8Hz[�W��Y�>��^[X�Xs׭�]�w�57:�X��t~���[2	T�R�(XJ��C�	�d��҄��K�܈�ѯgՠr��s�T���4��2W�|~��I�6KYk�4>G9/���Mʜ���@ť���g/�]S=�4�/�������c��y��^(��C��j����u�W�r�o�������*̈́x/�ݹE���oV��{���%� �z�N�ڨ�Q>��vg�9���]�'�w�:ۯ��+���u"�+j9�n���d����|�9H��`-��<
�മYJ8SV����5���n�����`HX��g]��A�b�����9����7�ބ����) ,���u�a�y��^۲ގӰT��8<�@]Sba��OL�/�*��4�q�C��$yj��oU���S�M]���V6��i��fct09 ���.�:����L���6��q�=I�7�+W��2���T�mB�H�}��M>��X�E��O����
;�e�w�uǨ������P���gH����@�h�h�H�a��<�g�l���&�`c�I,�����(\��qsk�_ׯ�0_���j��Iܻ�s�O)�a�U�����ǔn��S^M�\>b	J �jo��C�$������n$5���'�;�2���R^�O��'՗�B�[R
d�($�h�KΌ���g��(��2E�Zt��a��3�/����k?[jC
|<�E�#S��W,T�ND���P�ޯSKa�r`�3����ZA.���l�=V�p*|����ӄu��z�9�z�R���I?�Grɿ�@rY~w�(g��S�
&+G��̬��8Z|�[;��	UO�L��7�Z�4���.?�HDT̛m��Yx��"����,YSL���~ܚ��	�!]9>@�t��#��h��79��.�hJ52���|�er������}(�r�5hI"(_�3���F ��}�ŝ[l�b"v�~�0Za�ת�</~v�	R�Rh5�r�pD��x����q��n_P�t��u����?^�7�+�D�IA9|�{��x�Y�BĤ��<Nk�(��z�7�r�l��aK�̏��A�
�K�Eb��^�G+[s�Zt���G�c|j9���V��1���)�KJ�i~d^0�:��I���!���e�	��$r3�-��8i@b���G#W��;� 6�ط܁g£ڢ7ƙ�697Y[~���%�Q	�ٽ*����7[4�m�,�1��W�C�0O�U���f�l�{�2���\<���l4�3�[�؁�:h���@��փp���VX�DQ�q(���� �r_&V�S��8q�r֠{	��`��B�����л��ev(;P�%�b���g$_�J.�����]��&���&�I�T��F���ʹ)�,*����8z2���go]=�5cx�F���}��|v�`����B������	��)B7�p�#b#�b�}��[�M�'7�`"��i�i��)�8�x�>״�����tN�B�r����q��]q��e��6!���0�k��EC���yO����k�����L�%pd�p�@�E�y�f�[%@��<Y2=�B�rT��^^>�)��_KUEݸ:���^�^�{ˍ��2���6m�c�k5�H>i{��g�S=&���Dc��_��]8'�18����k?��`��sg1��3y߶�����;�Y��d>^W,JI�X�n�,[��O���b�U��/}t�a����uXW��dN���
�CG@����Qh�*Ќ	���=��5g6�� 0Fi��
�f|�i� ����j_��GX��M���ƙ��H�y=|�-݀�W~��U�8؛Z�ܟ�J��U�nc���q&���a��E�Ֆb�z����jNX����]�B�	�&���ꥱ��x�?c���1m���-$�����U�;q�q0�
����%+~p\�H�D���H�;|��#��!]D	*�>�ԫ��Ɩ�J�{�]���~����FW�_4t�XG��x��M`�~Y�yBA�4�R���ٚ��,��Y5h�}�)
���6�ˈ{ ��gt � ��6H������ce�A>�J��u�l�X�jűr2��S�0"�u�`��_�śR/K���ش^���+�Q!0�g2���D.
8�׸>�gh��
����.T]�ό�;P�+)fqr���I�Z�p�A^�6Uò�����r�\�W:XY����
>�M��i�w�$�0Q����e0~�}(*4�C����8v|l^�J@{�D��po����IZ ��+a�㳵N"r���륻��y,�i��-����	5����@�0�h>�X�@|�|�sgLѡ3V�t��Up����=�����A�`���X�W1)Os�L��^����ng�hO��
�>�ĸtL*C�'x�pm5���ʻ����oC�`@��"*K$Vp���\��Т������ַ����D.j���gL-xtߌ�.��,~�/žq����`�=5�m��j�k�q��P�#ۡ?�K �<.kVV�!���0Z�~wv�Z���Z\˿�b����J�d�U�X�)006���3n�5�
}P(-Y*䜃���W&:�:0�?-(�%٩�\6��H��Y��� 	Ϟ�2��Zp��U��0j:d�� > �<�m�ߍP������+DUd�8Gl�@+b��p3�'�M�xI�a�˷�; 1j�TC����OAb��x��G�na��`�)c�]��#�M�vv!����E��Eo����W�2j��q{7�>�d�4M����������YB���	2�+��[D~�᭪��E�M���J+��"�2#��ddg���{���U��-db=�W��3�P�`��ʆg�:�f�n�A�]��i��3���%#$Ue�L�|�����)�J���ܲ�P!�9��-�`02[��o�9���(4z-ޫ����2�E&�`����)9���@���dGY�Zįb�}��~
LFr>��
|� �K|�� ⁲���%�1���%$v���Db:��A^isZ�4Dv�<�v�=N�P��jA�D;`�Z��������[Tr:do	o#����b�k�z����0F�3<��=8���pnɅ���?d�O�F�+�&,�*������Ec��k�����Z��F��pG��E���S��k���K{�x�f� ����3Ÿ�y$��C��b;�ν�������|�w)+b)�g��r0<
�0�ɾ"���^��+Q�ޮbc¶j��)3��@����g=�p���W��3�"("���`Dn��5+���@�VChw���u����U�,L���:�h��-}7�K��S6>�?�X��Z��ޗ4/��`N,�eA�]�NK�'�;�s��z���'�$@ڦߨ��7�9�u���w:8���4(�����~�-H�L|"+��^E�*�D"A��G�ϩ6���Q����א�t`�j�z�B�x�%E"��$E_�4�u�:}L=r�0�(�e�6e�<�ɹ1*�\��Z��Yݎ;�n6�M{p�]�a2���N�0<_2}�@��A~��$S*Ep:�~�0��i�|£�c��$C�䛖�4@7�8�S�8?�_�T�rMz��U$�/�{���Ӈ95^�\I�h�k�9	�k��lf����I������%��X<�����O�k�4x����y2���)֘?�׃�È���x�%�*�U���9l�c��U`
1o�U�Y���bI.k��V��
�E��j$а�?8R��?y`�Ł��U�G�Ih�����;�d���~��j�@Ÿ�<ܶ�æ`���@@�C�����e�6p�F�HOgr��|T���R�VƧ����Ȇ��J�|�Ȟ%�0/���͋y�h����������b������i�S~6�T��a}�mr��L�U)��ً	��M�Ҡ$�x��"�Ҋf����BvT���+�T�)|<�g�y�F@��ś�1a[:/P��Zv��AH�Vl;��U�'�2�.�p�����e��?Of	[�����|Z�H��g�~��v3��M�xp>yG�\��:=K�z^�Ս���<��r�9f��牄ZJU��tx�`>����H�q�C��3���Tn��������	�*?m�j���;��4��O� '"C�D�D��و�M����`5SU�j�|B�nNs��2�`@%��s�LO�拇4̯�����PH)k'Ik���2m�8������.����b$�Rn�G-�e1RL�EL-�_R�e|��V��.guX��մ�+V�a=���I�ͪ���31 K�73��a�uhy�b�Kɂ�B�V��N�Tt�-�����P_t��3���,��3������i����M���9>m���{U�Ѣ@�+1����Oᴤ:]��=�ڡ�պ�U:����Ŕ8�z%%J8,om;�,��i%1چ��� ����4,
�[�D�ر4%�JGk�'��Ӻ!��s=������X$�m3%!��uϒV���!�����:a�1�Z�\� �Յ�o$��p���)�#��	ٔn���x��5a��<$�F�X�US]�}�Y����Y	�KR�	#=b���aaw����Q����c=_�:����اj���.0���_^�"<��u�-iS�2����@Ⱦ/J�lF��?�?�Y8¼(%��;����������<�G~�}k�ӫ1=����3��έ2�#H���խAKvȐ���u�Ѻ��ׂƀQ�kS�[�0Ӏ����
U�`PG��w�'2%����L��ڧH�UbC�?�&#�2Y��'F���c�9,��a�@���P�P9�Z��O�ۦ	̈́��>Ɉ';?�~��0��v��Ik8];��L��РM�#]c(�T�|�����&��)���q�n�",g��iHC	��0�ǛO`3a xз���L�%g�����&DK1��_�ʮF�"�=�˒څӤ�/�գ�^��qi�,�r��X��������B$t����E�m_ �aUn���M���͆��{���]�0i��#�'�d��� ��7����[���En"�>oro�ΐ�|�A�w�*2g��\b��QBt�i�t��H`>�mr�g:�#i��M:�;�#��@GT<t�O���!�Ŵ)J���+F#�t�@�2�'ۖ��ޟ��<���=al�V��B���������x�0�S�ɍ|<R�S�f��Zɇ��$`?���6���P+,`���;�0cl�&n�R�ݫ���U W�R�W�/��.��FŚ�TC��Oc%�|A�j���@����T��?<fˊ=�1���Ȼ�&���9\G��q^�+@Hd�y�Pg�hw}��� A�]������ڧ���ߜ_���a�>��P.Kzƪ�`!�׼��Q�����*���rV�"�d��f���ܑYn���k��sS:��ॳ�l��se\�/��GH,X��5@��'�(��~<����jx��
ɺt��U��/_��|?���$�������A�M�(w�?�����8<��:�D�.z�VrH����`}ɉ�5d��b��
���6��R����S��._i�hB�W	��Y+��F��瀸<����q�^4Y��6��4� R�����t��d2��D&�+0#稒&�j����r�&w��W��I�4�b)�OE���c�}bfyG� �ڝG��˲��ӕ�3�5B�i��R)"H>�X���Px'Wi^�*�s�~tv�����+Ӄ�Ȼu+��a��P�B\��[��[��x���)����c~�F��7�W�WF��o� ���G�4ݕ�U�;��´���"k`2o��"n����<�feZ�l2����W�(́%����IǕ���J%��PFէ��'���F�xt�|G�U�E��
���v�QB�, ��W���Ng+H��,�܇į$�do�@� ��nk�1hSܫ��E����%N<����<@Q�������PC��nL�	u�..��^�ۢyy=X/�k�[�}�$ʫ�;w�9��&}�
�出�z���}�x��=�#v@��*G���8(��*疳�{����G^t+	�6�`غ.�n7�ٍ0P�oZ��R�e,��{���2�yw�t�%2̜�y�-\90����/��" ���$���Nኋƞ�y)��
��p��|L�������BL�I,��˱�	�����q����$�" F����q`�'�b ;̍8�S�V�"J|��I�w*C�a3r
�Hь���3��lz�E�h�mTJ���z)b��m&�i����6j���>�=������͗k'���<һ���?]�P�aΙ2(B.�.,�!�p�K��@LR�����R��pF�
������)1"uU����;���O�ѪŚ��د���j���%�B4WG"f����_&,g���bpLN�D�{���g�w�)f㣽4\1�DC��3/�D�u�A�[�X@'I�3	��c0���u���3�@��l#�*���!��Ja_�W�d��g�}N��]I�.�����`4)��՞W�(����?m��q;�Z�<J��h�#��?̦����y�[Ҝ�x�#�l���su6ZWCP�:.��"�Ob�z���5cے�7f��t��,�::���эK/���O����a�b����)�i�vsʄ��	��a�1;Yf�Ζ���z���y
���G�����Q�>�X��#�̏s꽖_�E�{ck	�a�b�F�E��ݺ������[gM�2���Ɠ٭���P����H9���j��/���n�)@6MA6��S �[��r�8w�,�~�_~o�OVwh�O�>���2L/=��Z]�^���|���\�h���լ�k-ͷh> ���%A�W�^ -Rl��?�+�:��l���R\�$��KK }�J��d������ow:���A���c�DySYA��J>�AS���w��Dr-Ų�G��c+�Jyd��5k̝�!{��eP~��8^	�l���;���Jw�. ��F;�����(�a�����K��5����1�B�BJ����d�����ո�;�O�Λ���>{ђ0B�H
���Λ����o�@G�D�-�O�)���*�Z���,�ǥDȵ���W;����&�G�zɟ�S5��x�}S�2��Z�M�e�N�8E!�G��w�w�.i�aee'g>-�Xc�>��9jBg�y5
"�L�^�ub{��|+p�)м�8SQQg��]���B��Bn͡��������;�WpI�4�t�&dI�-:{�V1��忳8��r�v�@�'u��)'@ε����������^ΈB��8�I�6\���[vi�����>e���b�$utTX�mz=i�^�n�-�
�}��9��t;꫃rڸ�L��j�(?�UL�W���q����)�.T�w�8�/���_p^��o�V�S��֪D���z�TLV3%$����e�����V�'Ź����$+��w\M���5M�%�a�F�d���b�L�rwK���^U��˗�66������8��΁aԔ�����:Cq<�?������/�`�Ԩ�t�l|�7A��x-x����{/뚙�:E�Nů�P��P+0~{8�p!�Q(����\�8CH~>�P\[�ޝ������o������ 7�c�b�����������<�^|T�(2$��d�H��p��z_�*���;����Kq= w���F� !��ڮ'f�e\�g���t׾s�f�>Uk3��eB��L����$�jA�.�����~�?v������Ay ���y�nX��$��
nҐ��"`�i��;#�6,�p�����ݺ8��RX���zA�a<�.z�yZ����!�03v_=h�HYm�4SS���1X����=ZYi���	�} �IF������q����FްַdD����B��G0���zt�D��(Pa��G�M��h�P1���ݸͅ�p��@���[ƋĊ��2������TZ��Cl�%xW��`��ı21~�����ټD�([��Ц]�L�i8E��ƭ�x���R�PzS��dl����q�w�|q�B֐e�!\�,�`���g�j���E`��꘏���'r5���?_m�L�{$��+�J�	���(�(��<��R��5�jC���a��`�#���@��e��P�^�.�C�I�q�Sà��3�V�EEU��Q��\cΗ�D���X ��6���p}�#�����l`z���g��h��^�W]jx�v���4�Z�S�/��Җ:�N�g�� nzьD����3=H�o�z�<S�ZˊCA�_3I���k����H�f�򜓻���Nr��uK���\-���yNa���֞�Ω�.Wi�0"y�գ��k��Nl��9צi�Ԅ�A�P>��1e�Z-�m�d�l9�(�?wQ�m�ö3ubIiN���{��"��d���m�Au߉;�����jk����e�y��<�����Ja��Y��[g3�9���]�����w�"�|g�=��ݛÆ��[�h��i +Ǵ�U���#%~X4'���@M����-�a>�;�7��Rj��+H��� ��cC�K��� �WҨJ�㌺ʹ��i����fS���~)�\Z�ON�H�h�������F���bZ���R+�6�&�����R�j��������f%��#���@K?+<�-*�Ʀ���C���h������A�ҟ�-8�=���BU�~,������OVuw�������>�eDmi���J��3�?f[�!���U�ψ�KVPlᘊ���R���L�^�ͥf��!l�j̼�9{#s�m�v��|MY�v��/z�N��_C+!��خ��6<i��濅D�shx�
5��#����f4�9.�<��//���.n!���x`�U��;�i��L��J��9c��WA�*�%/]�*X��}^r�E"�$)�&D���'���Zey��J{}�����Xߍ��:z�{���E^i�6�H��7[J�(�K~\޴�cY-��Q�����!l?�3����M��z�*���lghC�'���=��ǜP���7���liw�ﷁ�}�[S��?��E�l��!���K�6�9��ip�V��e���'���IR=��Y\�")��G�v�؟�G������q��Z��c�Ӕw����P�tr@ʿ]'k�$��I10�$[E"���T�>�L#��&(@��}9�	 O��ӂm�g��!�;,M��n�� �����4�����|^v@�UA�x���\�u7S�N�^~�����x��K{Pfӯ���zg��=���Q��4��$����!�$��w�#��^`1D�������u(C�w�8a��=_LS>vf�������? ��8�U �_�iHz���a���<Gjl�Q�l����>���T1���A@ߨ��*䜌�u�:�-�y�r�mr��F�a{п��`W(��36H��l����ϫ���؈9B����_�>�d�kc^ʶ��4/i���D�Ft�=��t�4�70����_6�q@��������H�!T�\��R�w������vyq40V~V�VKp�p��[l+x�ik@��?� ~L����`���q�9��O���@Q9;�_�:d�6j4������;B\�>y�ǓA��H�~E���2X�CA?:��8Z*>$~�w����t�C�C`�>��oЂ�NK	
��G��?��)�����oK� �_�L]q�a�윥����P�Ӎ�a��������ι4.��g}�4�� [{'z$hD����*� ���bigv�i7�r�������S|k��X���9zF��Y��L.$_��|��$������'�R�f�;V�aWj�ky�)]{]F�0��b_0)�vl6}}_ú �EY�z��&J����5X'*�"��;`9;�B�2X���uJA�*��72��aTP�7�f�?ۼ��|%x��T�:�V����s��	g��咧�{f�!�Ķ�g!Q 7��x�P� !d��K�h��%r��6���=��.��~jq��܌v �.�Y&5��epK���<H+����=���	�m$l�uh<�d���Z���)��ɮ*p��de���>�{�"d �NU���p��o��N%D�}ESR�����[d�̔ҍ)��`l7)����T,�����0��		��V|���LO
ymHk��8@�)!JG�����ͮՕ��Q�y�6fE��"劁�^�F��݌���,�h=>2�@�+����p%���.F�^�{�S��Z���[$��^1���cWĶ�;n�b��K�Mޕ�:��>����7@c��ti�X��]ܺW��{4� ��U+�1�'�󇆈 B-�A���⣗PB��	B��?��3�B�Օ�x#4�H�K$�Yl|M�}hU�jC}:,�ӷ�~��)�X.?|﷋ ��������Wm+�~�v��v�~�����m�(�������|˸B��%����Gfq�v����D�RpG���E��l	��dc��1��T+Y!>6db�b���_��*�~�u�(?ٴR�{��!V�%��D��E��2�z��Z��N	�g�Խs��'��Hi�
��A�>*����+��lt6�� ��P��Z��A�#O픝c�0E��p2�D�D���[�|��S]�_��g��T��,
"Y���{��?cp�x�5�\e'�
�D{ '��O�z�x0�b�ܯ[�ԯ�!��i��-�ե	/6i�'���U�_7�˟f���!�Ke���ԛ�1.���ӃCB;�]��`E��9}��?���1O�c�c�$b)�wkI�ִ���"&Mߣ����\��*��9�E~��m�_��Ɣ�$�&��j�V��ʽL"x�L��Vـ]�����}�f�fI�a��g��?����תM���+�Ԝp��<�W$�%�>��#_��Z��xJ�أ` (u6��ڦn�:�*?'����{��W���m���5ݎ*�'*ޭM!3�??��;�v�Eđ:=�L�*Kw��Ȗ�;� {P�L�~¥T�����J�	�>m���~B�
{&�A���o1��A����O���k$�ڷ�t0݄ߠ''��8��sw��Ȳ��x����Z��tG�$��|oM�b8�t��-���0(�D�gX��UY$�\�/�;�Ԝ��;��f�m���5�����;[߰��!CU��S��-�"!e�	�~j:�뤕p���X�EMR��0T��a� 2�P�1�oZ)%����G��1N�r���J�����Q��_x"a�C��`O׬�64l��I���!1*¬�u	�2���9��L����y��p!?�n�-�����~�o�2��->U�n�1�FyU'��@З��+)i�w>��l=26��FDTF� ��aVS�.Dɧ�3���/�N��.�k"�"�+��Jʙv�5'�ת�t�U/X+�]�����&��Ȯ>����b�<6�b�t��!P�'�����t+���9?LY�P��A�6qf1��*0�#1v[�����%Q��vO��< d��i	�*h��hv�Ʉ���Ǖ&l��\�����2N'w������䵱�9ԭf%�ɜ�n1K^�E�(e8R3h��q��~ �4��I�V	A����eha����6���6$:1��և]�x�w��yB�
=	���P��zJ�����Pm����n�����V$�j
&�`�S�[#�z�k$(E�ú4~�{|�%3�ݔ4�ER���8��!���:O�'�(DF�9�;�lH"��u����͙d������˶��C��lIqn���Oi�k�F��3�z�ٕ,Zo3�0����r״���)�w�͊Oޞ����T��չ���U�wA1��M���o��1�e6���a�x��aZ>gT9&-j�<���ozx`:;E)�s�Ϟ�L���A����X}|�8�A���P��-&��g��Ѳ  �$����\S�R�0Yޤ*ȅ\Sh��6�l��&��jv���LV:�إ`�Kky�VBi՛)����5T�Y��X�{��L���ِ�@d&���?Q��b���iX�>{�.�y����w6�3mTZ��Z�C5%c��eGh��϶��������gl��Q��e��cF������l��AX�PA��E�~:�ӡC�I�`0�zvΟ���X��ש\7�:��Gs���I��x� ��2���X�D�_�Ĉg/�=�`�҃Z��� �(�`SIsR8s��/���"2괫�zE���0��E��T�@�4�5�	F;*�O~E�K@�[X��b{�l5I&%��v����{�#_p��z?/�\g�ry����7��ZQW��ڊ���y��П�7�GQH�x!��r��E ���`^~�tKKRИv�N�����P+�&,�g�*G����a���gՖ��)$P����O&S�S�V!8��ދ���e�_2>��Ⱥ��!ru���I��!�=~hr������_5����I5j������_�[��ի�E?e�V�ر�ꚻ����Q/�t���ك������C�&}��غ*�;���)A;6��7e�:���]���

�!���(,4T��I׿�d;4E�1=�U����O��!�I�=R"Τ+�z�'7{&&P�O��m��lR� =�{�nϙ�\&�=^%/Em���%t$�{ p;���6d��'4�H�7�"�|�1�j8Q���L�h���@�^ND�tPC6�0��3����E��FJܪ:��pF��1&tZ����'ڕ@���x/�����	�XL�e���.�X�nK�J�4����F�3��^�^'�%O/ې��T%q��l;��3�J���I��H�u�y���l��He-��l.:M���*�J@���8�O�1U)���;�|�$��P��Y���v�1�r�V���S{$�=#�T������87r8���{��y5S,�N�4yS<�"����_H�EDwX�Ԇ���D���������u�y����\�؂B�jD��Q`5�xN�I��A��+�7rɧ/���x�I��8h�j�l ���2%V�_������sL�_m��8�$��/҇��m�4��m����j�,��:xgg�,��7��勄��r����6�_�:�>	��͚�Kj�j���W�kHӇ�h	�@4T��sD�c�T��`��e�Ă!٤����3S��I� ��v!W�6�h���� W�[��c���n3u����5���&����S�d�������E�����Qط�p�!j`���2�5��T�'9�3�V~n�R�k�:��c��Ps񹚂��V��,���©�"��_�1�U����� tȡۨ��bҟ���Wڈ�+Uwb���.�v/�fXp%�����B�Y^��3�.�Hg�gd��JV��5(w�#��3j�2�N�Kv�O�2�N'O��+�W\#� Qu2�Eeb���֌��j���J�aR�	4׋`���f�?L_x��3	���ҨHRYɘP�r�����J�]f���)�lk��bG�.��q@�o&����xo��n���=(Q .�G��I���ĳ�p�����߄��87u/����!�A�5\Ә�\Q�ڪ��Avaۙ�9��	����n*K��Ԥp�ȔR��D�<Jļ�r�b�+nb �h�-C8����6� =��Xk�XL�ňex�H�3"�q�	�c6<�R3�K��:Rh"6��+�^����X:5��Ƥ�9@%��kZ���Z�T jV=Rm���-�J>�ƣ���˝(��r>"e� ����,f���C��+ξ�#����If;���H�M��¯�L�}	yϿUW������'�S�/?�@�(��f����L�'�V��Z�mp���`L�A�84Y:�����7,J�O�<S����<�r��%��o�^�]zy�g+����T8D� de	�B��*�ml�K}S���ܸЄ՗�6�AB��3oXLZ��n/����������=R��VX��w�fO�;
�dΌU����J��
�E��%�锡Qc����+�E	<�D��'����Rۻ-�-���dn�3���]�[y9B��)������IX�7E���A'�6lN�[0�"�0��!Dq�:}�/5h��H	4տg�F}{�'�ݓ,+����C+�I���q��{�N{t�1���,�Ř�M�@��l���E!v�?ۗ7�JWGS��&�9��y@6[.:i�#��o?>/����`.@°�sEb>)܊��"}�(>9�4͒<[g9��Z=��Zd�}�HH��� L
kq�0�����%��1�5��u�����V�ӎ�L0*dgadxM���µ��P����YM�����_7?e�����μ�q�g�ʣ,ͦ�E�Y���tk2I�g�����"i�1	�`@��� �t7��`����Rc9�Q��Έ�� �vd�Kb�E�QT�UL��cX���ͱZ2�v�q��5��%z�tI����ҩ�X�B4�.�Y��kp���?Qh(�!(b��0�j�A�\{��6�(<e9]��5�dG ���	��|�/ڼ=�����ƭ<�]��4{0[4�h�Y_KO����~�6��.���,v�&9L3���9$�	T  �ڈ@��яf2o�\�JI���$6����4��:�;���Gw����\����v��!6}�Z���0KL�o�]9�5����(�\�4z`w�v����3�
�w�CgN?�HO�_]bJ�5J���mƂJ�3�J!m��=��3�{ս�V��=W�p�d�b)t���L���e���FE���p�R�p��K�IN�̒�1��ϔ̿���$e�3�w�9;��&aޱ��n]u!"�_l�D��zz��h<�� ���g$���m���[-	���'����hQ�G�˵sm��(�Z(�,�W�V
vΪ��r��I_�зX��e����b�BK���F؎��s�)�M[p�]e=�X�^TռôIb_�#b�X���jϻ�*�fw��&����eU]q�+�0k�,/�_�P#�I�����qy�7��<QQ٨����U�7ȧ*�~�
.��ǂ4~2L�R�:�����"Z2w��·�#����)Ӧ�x{�^:�;ͯ�6���9��b��$�)�tr�X[��9/@�,H��q&s˔fR���R;~���V�u��[�FH���k��|�RȼR�P@��B�
w"��2�Az��V�#O �ڨk}��
��<i�LY����O��Ù���P����(q�J
�D$����w��G>rR5��*���j���
�,\��7��ިSk�ԹXC�8�<+��2�vdU������r�=����A����,��Ԉ�.\�Q�f�zJ1�B���u�ਪ�֌k�����"9.�h,���W%keo=�Y<p2��$�J⳹��&���c%ڻ���*�t�
��>�)���ٛ�Z����5���L_'�}�������B4ʟ�jv�^�)ˊW%_i.~-��-�"�:���(c��a��4�n�q����AV%�<�lVU����K�!�P��|irl�Fd`�o彝�h�OaOY�����B9?�mY�Y+��|�_I���Z�A��o-##oխ;pj����+�Y�ߎ�3�s8���t�/�'�A����,>0f�yǚO��?���v�iu�@�k�����e��k���A
�Y �Y�}�S~���L��I%����[e$bH$	/)kpE��6��ľ����	��sPtb@�i�x�f�l���l#t���`��ۙ-5u��nl�O3��h�曱Cq~G��TRl� z&���w���� BQ��a+��k�W8qwu�}˿���=y|�;���Ҭ��[�_h��;p��`�*�~��hly�6��v����9?%�%�����CS9��>j0(g�����IߣO7��.�j��,p�&en�*lo���Kz�;�w�]��N��2��.8�No�5D��;�fq���^G4��]v�ڭ�! ɯ�f��V����EO]8I@\N�+25�M �����=R�2���������%tś���:�w)����u%�}}�)83�!R��7���>���7R�&	�����}X�O�eC�����J��!ۯ�5Ŵ�%E퇩���k�Hh�۝��ʋ���bjg*����뭅�MmԈ��Us̨��0N�|n��v�S1B��������{���x�^J�&R��Z�7���p�C���?Pe�Q�#R�!R`��464��c$���4$�����[��]�GD$ f%�p���ܷ�7��x�k+�	Ȥd��/ȹO��wp��"[秎�7����Ο��B��)���\�@����/�/CS��zK4�uN0T'�R4`k!ǿ���Im�:D;�s52��ao'h�?hH2��&? �{��Ɓ���_"4ۃr�ó�p�Io�MT:�r����b��aA�;Ɏ�_���㠝�}��1|76��u��3� ے�������Lp��)���?�+�����ND����X�J��D�5�v�i=A��0�Po<,b��(�`!��Hg��Ł/�̧�n26�Y^�M��1�ǽ���2]�Y�-���0�SlTۃvepk׃i�����~X�"zfKV�yќ�$C'O�q�M�&���u���Y�jct��7>_������tz�5Lx�*��?�]'�;�"�7m�zptu��ƀ���������̆�VB#���&�T��KՖ���^q��X�溳�X���EZ��S�J<L��{��d�R�XE���\�@Cu��<� W����vߵ��Ǯ����|uw�7S�Wʦ+VG�<��)�J��R��,es�I8����"�������3�$�hØ�!ʷ;q[T$sRR����j�1&��p��
M�~�uz#�i_����!�=��k�����QQ���s�-�?9G�_����8���Ɍ�6}C̥	#:�H����m<B�!�#{��U@Ş7��`��J�7��7�ˑp���Y۟_�D�o��>rZ�8�v�4���Zev#�¢[�~�����]����K��a���g��A9�=��A�n wu��Q�hoK�2���ft������W�6�ݛ[�h>��xen�M������.ŝ���i�#���4Q�)� �KOR�I�8���X.}[�@ߵ����� b��/T��A��5R A��!�?ⅳdf_cN��qd�C���6�U�����������+:��O����qk�7
�Yc�&���o���mFL3��Y�4Rm��T��z�!�j�N3a�#���74�,r�M���d�[Z?��+�*�+���PUc2��:�;j����~�'sR`��0�u����W��}*aq}7�K���KO�W��JT���3j3�׆~�Y߆�q?U��+� �`ȟ��"-u�	�s���}d���9��u,
�y��'�޵֔'F��~�+�p�	/��z�"�xQnN�]~�	(~��������YVR�|ѐ�.w�	����t/�ʫ� 7E�m'\�oY�fi;��Γ2ZK=����.-�����ÍЗ�z\V��
R�N���F(<���)�� p��ʟ:�L�.���3u�~pC�(���޶��X&�v���H��ʆ�t���"=>GB��[6��}b$C9��wyB����@�H��*	0���k.����]���}.�{�1}-�
ɝTC���M\U��sk���|��^�A�����Vg3Õ��
�b�E�<��R�oe8L��v��k�'��2��_�L�3g;��@!�D*7�²�V�1nO�,w=�&@�G�S�$"���X����AM�q�)�t��Y!��	�S��zg�^��O�Cb�S�1���X�����r5�X��P���wdZ���q�i��IId��UB�{�օLt����4E�Q�J��o뭛ĳ���=liQ�hp
Aq)Ber=	*M����P���z�#�BįB��렷k�zJB�ѡ�6�`D�'�<���1�͏uC(�hi�����v��)�e���0����W
��n�`�	��	&Z��THj�$e"���(��N#FP�3V__�h|��^�q�X��ĪD�������5�3IW`͖±��� l��ai��eL�V+RgY�����TeLd=�=h�=]�x�jp[%�>+�ǇU�{g��ҽ��d�B��B�6���l�>�M����.>2�p�D(��'$�,�5� -��3ib�ք*W>���|V+8^p���餧���A�h!�	�1c-sunUe��R@!tۯOP���C�;�*͞��[F/�����-.����#o\�W^r�~��߈Hk����"����U�Dd�qz63?e��oYo�x�A�`7�
�����2�l� mm��g�F�P �Ł�b����Rw����o�g;�F� ѝ�ϡ���kq*/�R�(4���X�Z*�!jF�P������}��˾�u;�� �q{X���N��7%��'͏���ǲZ�`g�V�{m�2����zO�+YElj߸��č��n�y����z~��_�F����w0�n�Ґ(�wĤ�ͱ��֟A�xl�`���m"/(����i@���j������h���x�(���m��6�����!��@+	/ĻA���+��@�3��RFC�\����9��ѽ�O4���u��rs�c0k��ؤ��f�R]id�n5!���l��z]^˗d�	����`�q2*���A�"ݦ�Լ+'�����S��JW�@{r
's�:�V��֧2��e��G	����:#yZm�eG������%�'�A���5)i���v��*>cMP����^�!��HJh���_�6����d)��z���6kAJ������(����
��8��WXH�>�9��jZ���ϲ�"�V����R�d��0�H"p'�z�k���@�4X����O���e16�݌g��?�VDC�aPn˂�ؗ�W�)��(�W��Z�D�E�c]n0<�mFصod�x۶v��ou��&�ln��%H���r��!I~����ȑ��h����TpJy�@�Ķ����fYѱk��H��N/�&{���_�>�7+
%��i_d�$���U��^�&�W��\A�.ex��e^w��6\����C2Hq��qF�)�B%<��5s��xCL/�1PW�Ǳ��绨����J��ν"�#R�}<�$0�bP��!X�ܦ�+1�S�Uj��O��,���q�6ث)�A�l#~��?s��VH����0�l���Ҳ����n@��2m�fr\-�I�c&=w�ٸ�Du��C#'�����%�\ՠdl�k��T�����6t
?�ZAoZ1�� �4$��9?�~�+�/�D�f�6��K�y×9�7���w+����ilh�-؂�����/8<��V������JQ˷ɝ9<r�Hf�3+�MF��QF��w��������d f9�վ������
ܻ.	c�i:�[W<&4{��j{[P�%ap����^��S�	�y�T�ʐ����3�:���[}�P�]�D�j����ʹl���-����O}�V�F�&�櫄"�����&�(y�s"]���^xE�{��R����&�ο���6i�z�n瘩�:iK᙭3u�@���d��}^(lO�]��!K=���}���;ï'+t�2���i2��"�o��PW�{��U�-�U��I��He.��M�u�g�o6��c�[���銅�)k�2�Iɶ�N������ँ[�w�O�!������H��8��k�u�=�37��"�Ԃ�;��N1c��N��L���=.�R:2u�{���o'(4�s�rB������y�X����]7#[���=��G>#,�3�gj��Q��}$����Z�\qZO+��E4O��
am���ۼ��'0�|�����փ%�ӑ+�U|����D����zin;� ��7TK.ҝ�F[|2���i��[ݙ������Ձ��z�z�����Q8�/��lG3���X�f���ݕ��>�>=Q6�@~ew��mν��%���<Kk��Q.���=PA�U�s��ƴk6�~�JQA����Q�HN�u�[�����FNE1~|�&i��� 1 ��N���$瑳�*,q�^p����7�& �ç]�*KA�d�$�'�~�+o���%�#i#_������1>V2Z+��xG;�zX������l"��b~�@h^?zߵ too!�л�K8���ӟ�H~*��Z�<�a	�}��ˏ,V��5N���>	o��F$M�H[�-3,N���Ë�96;���r�@.{q���AX�i����fT�I����:��iB>g�J�3O�r����SQ�ta~���v��.:i�N���0�����Z�IƯmi��k��H5J�G���[��R��ԁф�����<�GI��Ny�9����79��D�4s5a�8��q%�#�c�/Hzŵ�������$ۉ����GV��4������7�}D�*I�Y�t����Ǉ���#�)o�Wt1r��,�]���b�g���c�#��Z�,Q�t�f���e�T?қ�U��� cP�����?u#_�Y�L� F+k��c�%L��uu.X+�7=P��Ы{+������=� �L����kZj�mГ�Ǹ'|�_��($VfJ���MU�@l��"X �����tZ�M&Mj娧B�D�� �,�麉��������>6���\/�{tަ���2c� ϹrB�&(����}����[�6"@�R��o��)Aְ7�T��
4�Z$U�c��۩� 
:�b��9�t�s�h8ȧ$\R����T�n��|�;^��*]�{�bt�i��H������W縺�=v7�jh�y�22)juẘ(����~_�Bd���h�7��"J�Pu ]�Ԓ��CL���LW��[���I���v����A�~�ʸ��2����P�y�j�����
*t����|�
�ۙ:�t5dQ�P~�ø߇��'�n0��E�&>�T ��q�R�d���j}t�ı�#�`���ASd�VR@�y"##�(I���g�u�qI��I���Х�Բz���Ϗ=�c��N��A�h�K��)ج��~��x���V̫��~u�Ҭ��=��e~�{��_pfwpd69�͐/po�mӬ�w)Q����]�L�^ϰ��6�$#�D�������颳L�q�v�T>͗��U8���N�6�%Sp8�6�_�e��Ƌ-zf5�����z��J֗�9d�U[���T�n<R��W�5^f�f�o�f���"K�������ԹC�HC�f�6ܓ���N��f}�B(G�e�X&���r֝��خ�~���B�w����/7�c�As�aARM!�l}+�����,}t�N��Z�w����oU�N���=�6	�qae�r���F)�)>Lu0�=E�^/%ƼP����������H�D}<�K һ~+��\	ŊƹJ\%�~g��q�dS���ƶW�dbvg�?p��'��9�+��&���劻��kZO�I�\�'��+�l��s�'�
I�0�M_�L}6�VM݁�2�hzg��HԇŔ���[�X����cTy�z5��9*?kj��ʨ�%J�u���Z �t���Є`��� ^�Ϲ��Q��3˒sՊ1�i�D���[�"��JV�|奤�y����{�$�A/�c�8[��ܻMe��|X�9ެ6�h.�#2���\��c���f��c���(�j�r��?h`Y	��e���\W�9�II�%�d+�Y")��' ޸4�{�s�����\ɏ"���诔CL�,�L-	o��͢�]\��:�z�������(��쯐�p��ư��a�+�o.�lP]��-��gJۗn���R����p֬�X��(�����B�c�{\��e6W��&%nC��T*|��Y
��4;q[b�G��J�m��n���l�r�Ч?�0��2r��KY����R����4�%�֪�6�?�}��X$�A)6�O��@]���S%K:�����$���zm���J��3j6^�̃��ѕ�}|�yd^�e��_�J4������P9�Pz`�5曧x�ɀU�Խ�/���:a�Kv�֓;bԥ}m� ��״&��z�%k;%P\'h�}|�Z&I}F�pݬ�"ʟ�q[�?4�bd�ʃeТ���;zrz��z����� ����K-g�l��PJ=Y]帨�1���� KD��C���؊����m@��2�v܄HE1�N�$���Le��v�__���Βi�zEQ)3utj	^-�#���^
{��	�qoZTo 1@���3x�>
�d�R�w�Tz��I�SJ�7bx+�~O��2��;��S��������t�Te	2�WE<�a:��t��P��if�fq"?�Δ���z�m��bN�u�k��U���G(�_28.������*�p�#f�mä���a���W��V��ٕ�-l�9#�p�����p��к��}п�@�?+��%��1	� {O"��!��noe���a����e����VM���Z�~��B�]����w���yѕ={W��h�2�Uֹ=�B��,~�M�B���Њw��9�.���)���>?��զw8��JQ%�v��xC�_v���}������j��&l�+�Rw(�W��Kk�A$���"n�3�2yZ�x��u��9������WwG��eub4R����?����2�ְ_���*_�����cGf�ՁP������+�,A|fI��
�VN�6UV����x:���S�u�?����B��ye	���}��}�4���˹�`�U���c<U��1�D��� �]��}2�t��������9�	��K��*A]u���%���{7�픪'@�'[3c$�Q!�F���!	����@�r����kF"��<VV�|��@�@S�nj�!M(L�3QQL���7��C"f?t&�jV=<8����@��1�N[�:e��!��{�Y����Yy5)��U����ك�#��%0h�ݡ�D��*��x� �����(��:Ww�@�F�t��R[�r��F�󠸄��)7�o�syw_02�
Ji�H�J3�K�+>�"����h,����^�Jj����z��>�ɉ�M�:��	�K���.�c[T�x?���I��*�(��l-�䨲<n,�TC����K�f{܏q	Z:�&�{s�;L|�c��a�Y�����63ءc2�����G��%����(���z������<=�jܒ>�k��7Bi+>��,c�1&+N�t��>\��%�[�b��u�v�6T�:[�ذ�F���@�����3-��y�9zS8y����'�0-':"���W���͹�0�?�aq]sw��I����9>�rҷ/uϒ2��F/krnݶ,r8��Э� �l>V��-�jrv~��|��9�&��9���M���k����-���io����H�^'�O�X<'Gёy�?��`��>��{��s�_��[0o����Xm�U-W�y/6iOن����n��6�Ф�`	v?d��\p�ݾ�=둴��X�s-�ipȔ�8Ǒ��� 	�9�Ѣ7��s�׷�GN@y"��X���Y�u�7$��_�>m��_�h�oɌ���f���c�+.��y���/�&p2WSB�s?9n&�X+�u��v����2��p�21!<资&<��~*�^�sA�|pyC�q+��Xobɫt��Xm��#��-X��ʶ������*�!C��n�#�[����ϿZ�&�R5?�g����'�+Cw�\1�ؾ8�	�+E�$���f9t�JJ�;�2Y�u�-�$�{$%$�>n��E���(�&ח����3��f�P���'���?��H��#H�O��i�����NĦ4Q'V�zM�FN��I˥
4>U~�����F�Qu�����˧W������/�ƁK==�*,�L�c��cE�(���~!���8{�.G��qX氼F�������Bȡ����(�V*^j����2ʺ�XH�Z�0抮��w�[��ޡ��X�; ٝ n$	��~Jk0_�Ryr:H�P�od�_x%���
�KRY봶�{��4���� %εѩq�܈J�S$��͡
h���o(�h�aY5ڦ�	���aeԡK�ҵ�\�'c��"��kg� v�����AQ�kTj*�}í�Z$^F1'�eSܘ i�E�nBʜW!��O�����TWW�!�j�ow2q)�4�%�8���;�՚����m�
��|{|��T$��Q5_7�0��� )9�G4��9�W�\IJ�E_ ��i2���2���}��U�<9�C�	UVH�zf��_7%�`�eT�����﫰^ukh��'n*��
�E����}�oWe.�~��_Zn���E��5K�FoJ������	P�� ~�YMw�җ��ֿD=h�O�G�L��#Y�c���杷*�'_k�I /fR4��8��ga!k�}�QS$H
��َ}�����q<u}jc�֓j�{�����I#+R#Y}a�^�<�i�_��d�w=vmU�nw�(֡���Y�z��������= �
��Dn�(!	�X� s7V�w�mkEh7V�3�k.����Y*�����Dӷ��n	\V��rXG�};)�xm���&BHZvu�~e��e^�cr�U�_G�p� N����R�lP���T�>��X�����/�e=��Q��k�C{6�9eF�~��i:Ȗ!ADa�g�GK�}?UЉ���R$��X9u*фs_X����Tk+&�����{7е�r� kZD��o3��"z�e[T���~�̄q��U�Y���f�#i٪��h�Ĩfҝ���L��M�7��g�9c�������u$ƂQI�M:]ـ#�h�	�T��Gz�C��D�ӽi�)K��R��r�U-��oh�T��z��QrC��s�:���g�;H�C]�Bj��_�fk�SpZ�b�g��ą���=���Ou�@�5�˕=�#�(X^���muTld��Ⱥ4L0�4��wm���b!3��[o�� 8���X9f��3cQw�>�}ryw\p9�O��f���g`_��¡`e�gsL8�q���K2dH��� ��́�m����ncxF1�������$��6�lJ��M�\��J�aU���h)��/��;�Mq��},���rV��NM��>�w�זd1lX���}l�Qʥ���JI!U�J,���a�$�_GF�)�U��h&1�L����u����O=d�����c���B�D<�^�5�M,��f���Z:Q��V�q[*e9{j�:�0�~����kʁF�&�9� �O�C]}b%���gJO�Ԍ��r����F4��� ��`��P��"�ƌdp����{�]�m~���Y�V�6T�b5�y��^�M��	VL�`Ė��p����.�	G&/��gy��!�{K��2Y�sX6l8�P�s����d<���D�d��<�-h3��o�"�=���m'�o�Et��Z��r��V��ru��^B�����r'㐴��҃3������%�#��:���^4f�㮄=�*4S�_`�G����t��#2;SX�h�>b��xڙh(���Cۅ�<?1�?�#��LzHN�_�W7P�����Ä`EK��f��N}���Q�`w�A�<� <����X� @h7:l��&��K9kR����]����T�)��v8�޺��n̤41/�
�G�O�Q�rl�H=�e�X���QTD����D������4٘�Ї�i�l�@8=_-&�&'��<�oU�c�D����-E�Ͷ#�����3@]�N��f7t+�@8�91�\a�P��uxM���{5Ӄ�W�a��j	��nW���?����BwJt�
�eFïR ��gDg��9��N�q֋#��߉Ԃ�r0��
2(s�(�S�/c�工�z���L�v��&EA��7%�8qc�&1�Z�m(Љ[]�c�#�w�ߦn���[�Q\�a��\Tmӈ�1�M�0#��{�kn�RN�{��B}�K?�E��e�D$��,F;�~M��:T�xj�y�|��qY�����N�q����HK�����[I���P�=K|;E �_K��(	}\��缺0�Kld_�4�N�N��øm��-��`u2~G�~7����B����q��[x�w@p�P?��%���p`l�UES��mtMX�	C�	��:#(N�K	����r,�v�Aj�,dز����jƑ{{k���S2������hN�y�Ezl8 /r�>�Ԧ�����+��@i�Ci�$y��1�/��z����]%pA`X`h���um���n����	l�N7���y�����'kA윿������7]�uQ�&>�S
7����VZƴ��a]��U�w0uW ��n�4w���bh�M���au�	o�T?c�}x���<�C�C��@��4������Ο���Z�z�A��xn6�!�W���F� *�Wm`���]����JB�!�����d��0u���@xj8*]��!��������Om����
I�Y�g�~a�_
������#��t��kH �(�B2֤�r���8��C�7�}C'=c؇�M�
2E�Qw�)�@�]����D�϶15��I��gKcĆq{1��J�$n^K����n�I|�r1B��[ ���V��n�)L���?��c�-�<�*k�nŋV��#*��+ܰ~�5w4A�]�jK`�w�+)k��G)���x�=��1dl$bI�$SX|�/���\�5��t�N-{>�S�)�ЅH9�ň��V�}hd��*�T�w�V�� �:ߪ��U��<�ڙ_z&i�i��������D��[e��X^@�(��~1f>�F�7���zb�l��-`�-� �u��\{S:��>Qa�5k�nz�
�%�a�뺿�T\�$&ھ� �fO���$g�}�Z�\���3jqJ�k&��Mh:�x�6�_���ImnN�
��|���<]�Wb�<~�R9_N�ot�� Y����D	7ĸӣ���E�|3n�Ę����~�	/}��C1�+�*���;����i1Tث_�� C���m�i���4/���tm+JE�Mzz���n�S٬:aRK=�6�>�`"�M��ev7?BhN^)H2?16��2v�5'��R'O��Y���;OiGځ�>��_���j���¾n���ŖR��À ��
5�jo}���X�n�-�y@*����E*Zw����1\4	�ۥ�$��@�d]�l|��}�#�&P�1�;8�r��SS�@`����|��|>]�a��I��<:/qg4$����U���,q���C�±!�a��[ө���7����剈sm��C��V�a�5����k+�Ejr��׽+�$�w:sD�P�Y@jJ4��Q�����OY���� ���d)� 3��
:t�*�VfêTk�'j���g��e
�u����9=Zd+9�[�Jq(3x�E�W7�"}J���Ǽ�y���/�d0'�CD�S�Ԡ��;�.Q`S�=Ϗ�Dtg�W�M��×��q��l%�OE׭�n�4�I{�L�ԓ�]>R�-���jrw��$
�!��(
ɪ-��"c<š
��^M����pa)k¾���jIkcϾ��7�͖wn�+gH9e�!�9���Li����J�%+E�nuΕ���ie'�,�A$1�o�b�c �8ԍ�����u1�U(N��M��DC'��8��J/����-����U�B#�T}�S9D���M
����N#	��D��)��J)@ѧ���:@�=��7Fw���l�V s{�9�l8�ϒ��U $E�rEK!/Ojꑰཿ�!�ǾEϸw��&ߵ"����I����k	(/�q~p7���gEֳ^��h�bZN��KVJc  +e�Y�ϐ����5����n!�I�-�7d�^��c�$d��XV�i�4_��N4�N8���<"Э)(���SMg�9o^���N�I�����8�"���lZ)����|nA��p���
��KvkS���D��$[���Z$����MM8d��6`�d�� đ'���3Ax��7�����8+�?`��m�5|/�{���\�=�mE��dU��)j
i��Ɩ8���Cb�&��h6���p$+��9CB�wO�8l� �]&�B����m�LZ1�~* ���,��m������Ԛ�_n�x7j�}��/��(����>�w2'�� j�NT>siD�XrcXl��:���eq����U��%ѨiI*���O����e�eh45w�_�NN��tg��Cim)V�iq�]XN?ɡ���."�R?6+��P=�o��:g���hx�����[�"��Zvd��6�>"��3���!��P��K^�7t�����ĕ�k�D;+���9;��gA�����^1c\��Y!0�ģ�h�$e���1����4���U�F�ꐝb�c0�kΎ�KW��)�!	61�mӿ��-/�k����BQ'��߰X��z�z�J��]X��!�.��P!g�~���PU����t���Ҿ�J�ڪ�/��H��E����C�\�w��з�IW%��Z�:���Y_��z=��J;� q��ܵ�Xd�+]�u������8>G��J�[�����n�\�������9�]K�İ
������\�Ү�=�2��ѳ�P��陒"V y?���u�N"ݴ(>Ad�k���U���$���vM�AWtd��fU�EK2��w_��̃��E�r}f]�c�bJ��ȋ��D����s��V��9�Y�'a�#Tx�8�&�$�'j��R�}���~�Z�c��:�q@��S��pM�j�����D��ͫ'�~��z�l��U��euŎ�y��~��w=f�3��č[I�����}k� {Q�I=.;`R�4~9����4�,���l�����@�'"��׀>��2��n�>�^��1�F��۷<~�`�I}�������C8�L�c�+��W���z���r�Ch�Ʊ+M�S�Hf��Ǐ���M�$p��`/��u��#E�o�_)b@�m��W����M`��@&4������&6��X����)[i��N5�'&��w�uvOO��E�cC�U
E~��bɞC��;�*�^y4�NK��z��Jf�EH�"U�v���y�}�<��ı��Rn���7��e+�L��*�,ј� t�Z��+����G�IZPbށf'���W,��1�o��U<t��}M����p��S🇨HM:'g���<�%R�0o￾5K79=��jo5����ye�	;��t�靼� ��w�0�0�۩6��2b�8�a[@ͬ��|��$u���֣&�Lu�
n���2�R�Kzd� I���E(w)�T�Gh���'�X/��44������)�S�E<����V�_4vI��j�!A��?k7ON ٯ�<+4��� AҬ��V{dD���&��M���%�a���Z�Y�b2Q��!�s��yR�^~�qK=-��������!�IZ5��Kع�5�|
�k_ƓT�eS��\l��'��j~��Vq@7�|�H��J���Q��
ԝ�mK��e�F��������hh����V�7d��v��$5��av_�p.a<�\?Ux�ȗ��Xg���E�����P�P���x?�'��g�{�js��t��q׵�.T�YH=w��H^���M�肊�F������@ޒ7�l���2-���=�L+�2̫&��h�_�D<��E?��c��l5��t���!���{��[Ǉ�N�+�6�4�AT��Y.a�}~��)�Hi��(����Vkߖ���#|+SQC��[<h�Y<a�2
V��$̆�`�.��ɗ����=��u���ڌjW�:Dmo2��B�Qk�e��MY�$Ĝ�ri�4ЀKJj�΀%)�L�n���I�C^�sK��ߒh��獷���X#[m���^�B�����
x٢u�c��� ��I�▋D�t���LkXf�h.�j������4Hҏ{�*�E��$gͰ\�j��N�9#�"�����q"o��v���Fs}y&��*�A⌐k㧥A6;�MH{Y��h�������s/����ȸ�yL��,�+�טrxWѿ��2G����E=J?��fi|^P���}���=�=Q2�ׄL7� ������i��x֛�՜h;�gc�~)��X��[�5�8�Y�r��mC���w�Hi��ɨc����8���#����B�9�(<GP�]t�!�XҴW է�.�	<��=�
E3R�VE��u�N��sרb�[��(��d��?��Uq���uk1N�ľ,fX�n��ay�	H�FB�A��+V��$_{��a�ǌ���+�=�̲������H�]a��r!��.ͼ'k/��T�Y7ǇL!x�����&Q�8���4��/Tշ0��QU�q"���g���T[ x�_N������<���v� h��i~nL�^��q�V_ԫ��B�f�[�����syQ��։HE'm�mA��)�sK�p�$M*+# m�P���њ@[��uK�m�Պq?���+f'�6�*��*��b�ZQ��{��)�����������=�b}�!�X��AVYU_=�3��+c��j��\d$l��VW��یa1��D9��|d'#P���Ĵ�ጅ��[/P�>���g"��iV�90��y)j��sIR`�:@�`�'J{�q.�m����K���p�4	��#�v����!���_+�J5��)�K�0U��6��>�1'*�6�v��-�����Ç ��-�m�T�4�^p�+'�����+p+�8�Q?��̠�I-pf��b8��5�4��VЭ�}��ک�y5���=|9�}(���n|�����M�+а�'�Ŀ.��)?���'��&�����f��2w�wv|j�@K����&.D�1�C@"�pܙ5nP�EG���=�Lh��jJ2>Z��Ę!5�{xl÷	�
���)ż�.m1V�Pb=1������H�6xc�F�v�xU�cO��Jï]gol����&Kv�.`tte�[�>� 6�^rѸ�J���)N���&*��HM�;o㙍���A�h���5����J����� �
�\��s(I�F�&������oeʴ��D^iZ폥�	�_w��>�g?z�[���u�#�Z%�N��X�_+�q�H��-���q��nw���I�������������ӏ[Gڢ�_��\�_�[��?gk��O���l��(8� \h�7D*uz��N�����ܞ����o���h��� ����b���@����,ؑ !���ؿl�[�j�~�g�=��9�Q���-�k�O->w��15��39��Q6���>"B`.��G}}�le��8�Vv�A5��/��*���.�l�?tI�B��� X�?ڶ?���춠���L�d�8��12����b� ��V�Sܷ��-
v$@CE��� �����*MȬ%���H���@��B��C�`j"�v@ϫ��};�o��~2H\|��u�1�d�|^�	�J�� i���2Ď)������^B�L��h�/.����3�?e�r�o4����D^���b:�\ ����^�<6���d��C	�תnBv��ڋ�ʲ�Ċ�G���Ã>��Lh஡�Б���t��� ������B\)�C���$H$�gp�M�,j�	�B�_�Β������C�}j[E�B�7��V۠	y�7G�KU�~QYS[�&�������KI�h�M��ͤq��m�b@Q�Ws����Ib�ȻI/A�5]�sryy�Y����v�X��D�[i�~�;J��[���Ivl5�����=[Q� b5
�4������C�g������¡U�����Ju�]��90	7��b��?zƧh_:�G�vT��,�k�� t�$;C�����UB'Z,���D�^��k���X�f�NF�M�����(K���]5�=��V1���[�.�u���"vm�n���6PE{E�訤'�ߝ���>YK{L�;��Y�YN}�6�t{�ۋ���z=��{���l�F�]^��
[��3����>'?�F�l��Pv���FW�m�On(��`P�����G�_�4��X��$��z&�T��K-H��cѓ��j^e!N0�������9Ô�����?��<��-Ƈ�M����c��֏���|�%�Ҕ��@Y�ܒ���\'��Y�T.=+y��b��z?S�WĂ<UF x�/97�^tɑ�p|-ױ�<��+E-a;r�p�{�(�Qh�ˈ�4�4F#l����(F�K�U��-_�O<	�-���ۅAX�A�m79 j�Tt/�k�0���\�~YU�������1N���8�Xڼ�$q�8�Rfq��훿R��+ئ/�����	o�=�U}�
��G��T�+/]����4z��@��d�J�I��Wƍ���K��|oU��ntى�?%"���A�H�x<(EG��-�Ō������T<��-SJZ���� ����,�:�v-���[�#i�xS*:���ޟLg�N!D�`�a�L�ܝ90��۾h�V9i�������H��a03t��Z���p���я��?�И��Vg�Ǎ<3f�E��sX������Ѯb��_O� 6�1 ��Wl�9i����^��WI�@�\(�p��̀#̆}MƄ������րye��$k>� � ?�{�\�|0�L�ְ���������phɕ��H��p�Ɓ��H��02G�?����%��R�n�X3�w~4b@�c������x֎����׉|��T���O�M��;�M�?͑d��5ײ������/�ԍ�O��l�Ds�Y↿�!��"����ՁxLh�����OǯP!�+``^�G�F�$�+���.#̡�ƫ��j��e�LF,S�2;~��*�go5�k���|���Q�=�3R�F��]H��\ޕf��%�s^Y�#�.��v"yb�m�K>��=���#�-��Z]ɻGq@ma�t����C�����YfL�� ��]	z�D(��
Z�9���Nյ�i�n��8�!4����q�EUTV�5M�ѵ�bv����G�&�P�(Vɢ�S/���
,[�w���i���iDx"�7�������]JS�^8[��|�����h�d8� ���nR�-�4㬳�r�=e����p\Cw����3S좵��ԙFU������i'�W
�G�AoAoX���gT�~�x�b;�l�e���3H�^�PG=���z$�}K~�L?�y�{����R��m�ժ��&m5���W?}l*�)W�	�B�o3tP�阔-5��DߐI��SU��W�`�����XښB�|��~�䬱[�&������zZ�ƒnt{�Od�r��Ƞ�#� �F6���Z!./�MT��xj�;V@
_U�T�����Qy��s��'��y81��!���*?�=c�:�f󢾟YՆ�v� ��#Q�O��k;>�.�J��i��0�	i�Qr8�rӠ�����p�^�!P�7A�fv�ENA`,��{�QW�ɷs�sosE�t��垒>hM6�5��T��7�$��w�vNq*fQ"+(i?�����fq���BuBAOF�]7`��c�_��(*�62
{�%�|��q�`\�h m�⁗9����^2"������Vڐ���F�RG�RLU7�`��M��**��Ϝ��wyv��3�!A��8P�v���u�����yJ���j��8>��[�MI��xY]�L�oׂ��QrT���UM��BYp.����������Dz�ju*hP��]�
j�Wq�9�t[1�M��/'װ�sy��Y�?�e������f�ġ۸Vc�)�Ӛ��3�A2z����R���~{11�믢��Zn	MRƤ�Z6j���Wr��:m����gj�N-!9���7�8��g3���nw9�L���k�v"?�D��D�#��n'S�1��«>�W��wF��T�J<\Lb���'\V8������X��{�$��Z^򭕳��ih�����U�
ʁ˔�NV�
�"P{�P˦��z�b�4g�CQ�"I�3�{��$(l���G������}YZ9�*Q ޒ3�b���j��A0�Ӥq�����R��xTe"^	
0�he�����	���)���a;���@�>��Wn��m�<isZ��䮬�b��ʪ���Z�Ex��UV
=�K۽aZ�~'c�)�Ʃ�~������ʋK�q
��Y�J{�K��)�]���ɀQ�h[�Z��c�Q���q��K�&��G��/FJ!���"���DI0�B'�&���7޼��f�
K �i�p[ ��*i	QJJ����Ek�~�P?��	�mC�Z�F4f?Q�z�޽�z�/g�~����A�e�cŀuS�;~&ra'}@�Kk�����otg�B	��e��U����L�L`OCr_^>\��f����C}�D�U)�����G��p|�a^šVu�IU�v8�P'D�?6	��5E��w5��N{�㊰�฾֝�4Û�Bn�&���[n�?G$(������DuB��s��/ r�����e5�>����Yl��E��yni�|`f|��Wq��t��ע� ����SE_\���`���/ޗ�ǒ/�-��^A��|7˰0X3���"���5v�2���.��-8:N��i�G�b�3��=ej��}�8�`�%򚨶:��,�Wn��W�]����v�IW���~}7Ds��6�C[-Ƭ����+��m|����拽�]}��U����c#d�<�W��̧8W�ww�leoj���"�
�ۿ=��2���J��/h�?�7-����F$��/���%���8E9:��m#�s����574�+��h�����կ��<�H��@�^QF6�ԧ'��k`�ܯ�;p"�5�/@jP�� �~�*-��o�禄�:ފ:���Կ���U���=:�]�؛�@&l%�mܷ͜A(���W0�4���8�9�A�-h���� ��I*,�<�Wxv�Z�{|4?�Z��W1��(�O �R�F!-�׏�"�\���vn�CW�L��m֘�{�M_��x���v�8R��DJsw���l_7�B_f%��"ܱ,���l�r�[~˝�
�0���S�%�ʊ�����q=D!9*(
b.`�~b7�҄�(շ�ի㺂����� ĻͲf�G�2/����9Iv�<�~��/����:|g�du2r'A̝����,j;?ş�ZK�����-���,�\ifIr|0Y�2V���w�?>@f9�χ�z�����{L!P!4���Id<7����A����������D�0��H��iC�K̹�z[���$5��(�_n�܃�5y�u֦��?�U�p���uz���W@Yo��C�ww�����vE��^O����>N9�A�{ĵ� ?k���ɂ�cal�.�a�U�k� �u!����V�W�]�5<`�}2E��t����w	����g���i2��(�xH�%�Z�El��<�[�˥��7J���C��#�G�3���z׽B�O��k�����^�������	��4�W_��䖔����oR�;ibk��m���R�U,ǋ�~�S0�����M:؊N|��`�+�}�b1���A4�Oưq3����X�.�	G����&]�zIO��K��Ć��%��z�vx��w�,��u��b�]�Ak7�MUD��H�Q¥/���p���<��:��x��u.C�������*]���	h���o�i���)$v��4���_��p@��}�6��┓��;�T� ���`�4��5?+T'��=�'UO�H=_��$�$eX��E�=aΟ�v���\��̉�~%KyIN��uڣc�׍���,�b]����v������I�����~2�f�交�4 `�X�E�⠰�~�C�WR���𯼰�c�z����/~�׼~@�SW���u\^�G���(���B�@cp|2o�(p�b��M@\ƃԏ�u\���//��1�$��R[R��,�~l��`qx�{V�H�'B	��+��س�P��V�fFY`��RƔ�龗��vo�䪰"���a�E'�NC��k
]r|\�mN�����!O7?O�\$�-��o��=۶�d�уbc8f�V|��I��Rx�#m���2m�o]��}�>����?���lk�:�;�)�\)I��(�O��PQ�9l֋3֚8�|���ii���EDe
�%0���G�6�[��t��Ǐ�ͺf#�P�<���<�������
����S���r��ދ6��-��"t��F'.c%EF��3�-�w�~��[�ۗM�]��'�3�l4��+ϡ��ޠ~�U:\�%��f{��X,��ǟ�%�`pJ$����[�#��g�,W���洭�$�4=!�j�!��z�����"X0�p-\�NР� ʂ��ZG����Ǹ��:ۓ(�2-��V:&f�a��0�˦Ti\K�4m����<�9��|��B��O��A�Ns(1�/��Ӓ�v����~L�Vȍq����6&Ha�#o�f�0�
���K��tC?)'B�^X*��_��.rG�����i�1<�W׿�͞�"ڹ�(�0��=�q#h����H'���M���@���YQ�.,6�מ6{�YH��k��zY��Y�8���N#�ڡ�ְ<aX>s�����]od���Q(?k�!�����	F�˹ kʑ��9���?4n��4q��Hzc0�Q��{Z^#,댊�u�=X�_�a���kg�7����)
��w,��d8<$n��tJ��d%��R�`en/IsL���qr�7�tG��H��,:i-�!d���a~�Q>��ٳ���<��T�F�~f�5�I����ot��Y���Y��9՝��$;���q@8g���鏡߻���^*�N��#�mXA�"��Q�|���~����,S3��?`�OU��ػ^}y�o���P��,���6@� �F��|*V����-����x�^n�1�k�I��낻�E&13����e�%�H*��+5n����B�S���,s�$%��J��>H8
9����saW��_�0Fz�e9�2�_#L8�H��8���/�u�h�Z����e���M�M#�wI\���ԥ�y���!���G��0i�SC4�_vzYP���u�"��|�Ϡu�(2�<R�i��)ۀ�l��S�hy
�1K��ܞ5Z�#%�2���W��\��`���%�������}(��ۚ�Ts�`�/��*:[�}m.�3�淵�+2�jo�"ٔ�rX�L��\�+3�˰pR8��;�þ��m��u N9�,p��q9���?-�������i���k��P%�OQց��[z��(
��I�ëi����d���i�;�h3|bg��1�̯�_����\8Oi�X'�D�"ۿd#$�p���7|Dn��/�`~�6��z6K,�@������,&����>o}�3�������H�P�.9m=��ᒂ#���0�����r�r'���b:�(��s�q��C�*�ij�OY���w�?b���z9ìxh�F�<z�=?y�i�2ӥ�:���h3���Y�geҿA��9�dy��-�p�wn�W�A ���G�_s���2V�^Aq���,qZ�����_��	C&d���c����Kק�j�`L���]�D�^u�5������3��I(w�����		���@q�t{�΁����1�ξZ���j�����ڔ��#+ˤ�ѭB���޹�奄�td�kp��J҇�u���qz�$�ד�x�W�=�Bj���i�k��E���F���d洫��Ƀm��@ߍ�l��j���C���sb��+.D���D ��9\�'��Ry�9���|ʭ���>9:�]�<����L\�}��`?��[�N5�Q'?ҳ�[}�v��R�#E#���B���Nve\_qv�s}}�^g� $�M�D�-F�~��v�f��:?���t��'}pCW��W�a���دTb�hLO*J���]�!�9�O���NPp'��L�{($O���V���R�x��h�O�X���bt�b%l�<O��Ϊ���r3���^��!~V��\=�����I�w��h?!qF�p�;te�rqN;�UeX�{�H�9��,��5zkB�*�Gk��[y��,HޝnG��j5�]����s�g�XT��JU���C�����_���8�ي�
�J��V����hZ�NA��#!�J�˴`���=��>I
v��rW�r��n$+�9�+/w��S�tH�mW��.HB{����4;ؘ����Z蚯�^ ��&������'SEfSCh���t���	�!)�ť��� �d=U�$��������"����Y9�������)�|i[!җ�%gg�ӳ�o:h��jC讴M��N���Qn��B�]�!�Xf�Ψ//���5y��i��y��:�ٻ>�C��:?�<��ǘ$�C9���R�vP
�T[�1B������|ot����ұZ��ݿX'����ץ3K�g���F�r��s�r7%orv�O�ĭ�+�1���Ÿ���;�����qD]�s�q�_�Gc��`���G�N�,R�3�ofs(���>����]�m�٬�`�UG��^&k(�:zդz��o�?1I''+m�P���F��R���r�a�Y_���< �,r,��#�W
jʇzJQ�p�o�ڻ��,.����o]&�\J�逴.c(�u}6�%�:����F�m�u��7yh���B��������2���O���ؾ��5��<�^uX�����q�U�&Ǟ4�~�|�p�\�>�GY��۲������/!U���)|� N�_��Eo��	S��lk�8��<��{��c�f�`�J���~�mj�H�be�'s�s�S�'h1o瘆�Q��S�t�s�_V�z������uu[�O�֨�T4��[A�,V,{��$�����C'e���/j��WFġY��u������!�_&h��h��fR8��bQ�k<�p�s$����O��,n�]-
��	��'y�3<��_�
�^Մ��B�H���$/��,��fw��Tڵ�sB�v��KuZc)�U�a�b���d����j���Di�,H��d�/$����>��`�T��-,����L��q��[�sNAC�-a��vߦ������w�`W��/��!sGH�N� %�N:0��N"������J�v9�,�*�	�a���zT�׭��	���uR
���ܻx�7X�r�#���Ps�p��7H��RDv[�=B�.	���F�������l��nCLt�}A��q��Q����>��>������ L�+�(�[�]:�	�y.�3�W��8FB0c  f!@@a���9�eov\*y��^��m12���1��e$n�j��T!��QW�<]6�FL��=���e]_?Fa����I��·�fW�M�I_�}�I�)#��*��!��f����Ӑ��y�K\��<�!��|W�Bxౄ������M8�{� .<I}�v�j�&U�brS�*�P@��{}�����ʱ7ޅ��h�xE^0d���A����Z�g�M��k(1������IϺj/IK�l��_P�5d `�X_9�\���[<tT~g6���̙�v��D��m3-8(a��d2O�~g��Pbq˵�2���1Y	A�E��X��p��?a�J�ykdd����uE��Ar�c8��IeN����w:�p�1�ƾ�M*pp�,h/�
���W"_����Y�b,�$��ڋL�16cQuU<��	���w����;�t+��n�;Lw���&w��Bș���Lv(
�i���{���,3?ر�"}t��<\O�����җ�u�&f�����ۤ��Ky3�º|?�>`��:Ņ1Xc�}�9Fr`���5jaC {��$;|��C�Ӽo@Sˢ��AX��$˰��oXԫ�J�M�T�AS6����� �郢nӂ�$����QFn���iX�˗�Il+v;��N�J��������]�d��T�nP����>oJҐ�^h��~)��	hL�Gr�T���e�&��]���u���L*�rb���w��ř+�bf�`��Rnm�Ư�.cX�J&��aeTq�?�B�VI;�\ǰ|�s���~&N�Rʨ�������m��54K���y4�"�]���>��O�qnF_ª���Q�ӳh>�nVƶ��������k�ƿ�����9��!q���ݶ��&D�*Ҳ�ȯT��-�ဓJP��t�g����U�}�t�kIW�u�	֧p�n�1߯��I�{�~
��L����va`
�'��iKy^e>_�H��
�S���6{Ut�3��w�gO�b(xj�݄	ط�N|�Q;=��'�, 
��$�L�~����� ew>4
��+����ˊ0!��p9�S�O�Y�6��8u|n/c��V[𔇣�ɛ�u<��vV��nˣ��b�+W������7g�*s��A~��/jg��q����7�����pY��2�BrOlw�vw��.����t�P�Ufrz�wΆb����k���Z"m�����?�dZƄ��*ϡ����*�L<͙�L3M�yN�"%5Z\ɽ-�db������?x;�4��3��[��S� �0�n�C��D"XP�y�����;c�W��݁�Q<
ɣ^�0��N�]��첖F_u'��	SSP#Y���;4��� �e���
��4Ġ�5�!K��@+b���FqˢR��E�G�.�+�$�ZU|�\���(j��:+�EZ����d�����rQ<�B B���GzK�(Tm/h�����f���J���5�Bm��J�9vy��y@r֤DJ�D��o0�Y�\"��r޺LDEQS���_x�|4�n4*��[l?�)��6�M��ʢ8���R܄�� Q���q;��(십���b8"#t�8i ggۉ�`|��#��iN &�	��[���p���v_j��Vn��p�EWl����(��'y5���V��'���iT1|���c��\�tڅ/J���L�T+b�쉽
UC����L���0�VǾ�H	�p~�x�����g�;A���A�<����R�y�L@���t�:����~av�(�6�����,v��531��+�1#��� qkr�74��b*Y�s�`Q{���xB�m���3�d����J�c`5K�A
�L�?��3�z�bxk����e[��m�U࠭z/��h��H^�=��������Gkg�,�a�wa��Ae^͹��E���Sb�E�pcc5���G2ǖ6�
�7efzy@�"�L�iM/�F��Q�xWv�M� �W��A��x$���+.�O�ϒ�uZg"�������[��Dߒ�q�i-h���j}��JC���3��\ʹ�&�<?��C�Փq��q!%��]���l|��g?��Zrp5���x/�o�Q��~��s����OT��h�(�mT��o�bo�c����{�=���)E2�n�f�#�FB��%�k�Q�j3'"�S��=���Z�W2��T��U�~��E�c��_�Ud�$Q5Jt�2@�bA�!�H��d��$�9<{���v�dM�<���J0����۞�)�!��ਟ?m�t��M Qxz��bY��Mw������0��ʛ���R|��
����1�`�x����A���e5�-���q�$��R��eQ�Uez/�_�*0���X(h��D�\�/s��F�zy��r���/���D�A�.��5B``� �ڛ6�U��&�/Uv��h���­ ;o ��s�ڌ���Ku���x;J����g�	z�~����U����]�'���*$&T*|�8��+���Z�'D��,D/�e��e��'l������k���[OMyeH0�Tp��A�tȝg�D_�,�E�2�|�<�x�asan��V1�لb��i	��S"��U����}_����̱z:�[OnIV��}$��V�d�t�Uu�S-b���GZڸ��`��:#7�w{�r��̜���A�Y�?�NAxo�k��K���O*��yؑA�����-�L���O��"��$�l�¦L����)��e	���iy0�x%�w���x� �B�y�&���8#�N�vRB�ӡ"Vf��tE#?X����n��7�9і灗��K�b(�h���z㮡�����H��������,�*�S��Iw�D�j�3��$����$����MN�l
�?*�+m3K�b< �i����ȳ�z]zD������w٘�=�(�*��46/QR�~��U�\��pL�ݏ�����[���3O*VVf���~�L���4���xKG���@��hs\eu+~}�F��4���t֠�?.��j7��Y\�����Q%�	"�H<�1��c�?3�ĸ��	8v�݃���������]\����Y��OC}�	��{�}�-Z%x�ʴ��IO��K�+L�s���V��Yp���Њ�+��-�_�N���r�^��i(5�F�y��5)�0��c,6�R!�4f�5����؆�ҿn%{)<�۱�@���c)��x�S����R����ϫJq<uŕ�Տ^�
��h~��wc�x��u�7-�z�دH�F"���:��( ua�S;���\��j�J3�u\
�L�:g��і%��\8�0"�{Ԍ����(���f��`�)7���I'*��0T:������NX8~�^��[Խ��L9aĭWr�X��3�� :o�u8~5��uN��)��� [G��D,�s)��&Bd��>�$&_n����`�5]M5��{�p癪���X1%�C�!��P#x+�B>V�T��	Agp2ރ"�cdDoh���Õ�qm@�d$G)=�U����S��u�Tð����TP��;-Ez�V&j���`X]�d�b.�p1mp��53�cgdq3���b��䞉.U0��g�0�nc*d���;� ��x���Pr&�H:-l�9�&a� �鑿����o,�ۨ��#��wCkR�ie":ޣ9�I�|���tҦ��8>�c,�E���_ݸ�vı�/#n��&ҏ�y���LlZ�|n�[*b���9K8�&Q�Uy~ A^J���u	������0�����W���B��DZ�hP=�T2� �3t�|oB�YR�q6�p�2vi��4v����;�
�u^Yaj��0M��Ԡ9廛>"U�Dk�m�5��o��.M@���s�}�>G9�T�$G��CfMd��[���k����su�W��$<�Q�M���m�r,�V�_4)6�K����Rq���Kyh��k���Nۙ?O�|�~��RsX���/�Eԃ�� >�!)|�7�b������_༉p�����i�����i�fU�ظ~#���oK�"L�V�uR��2|��jb�dM�`�7hL!L����c,���x�'�ٸ�f�e��6�4@��0��6�����)��6w�d�#�3�D��L�׍�(Kx�L�8�t�P�%�Kd�T\�Sp����!bȦ�y|��{^�$��	� ��,���N�r��-�}�LՌ��āA��[!k����f��[�״�G���2"��+U|1$i��l��7l�+28�J(��Q�>%�k�p�1R<�WuR9�9��������g��W�AЧ��&��.��Tɠ�9�ĠV1��us��6������u�Ѹ���sZ���9��2�bľ�r��D�����3oIU���5P�����E�������8�CFpc���[�[Lr�tΪ��g��O0����i�f�p]Jzמ@�dw������xV�\-���i>�D?�0�hQ� ���)2��E�/�1�%荢a���
�2��iSS��p[G9�IDA�E&��P��s2TCڨ�6���_��@XJ k�2�=�hɶ<xnBy�VL�uH�"S����Ȋ����
��U��6~���-��09����/�-Y�2H��Γ�O�T���pT6�5i90�&SO���RF�ͺ�:C#0�L-�VDq���-���Da����_��n���u@��E:��5���IN������ ��v�N�晴O,�Ό�􇃁B���N�}u󢾏�?�=��<h��1�ʚ���<A���sy����&�����w���phQۅ�ac'b�B]N���T7�(TG�G�_4�,Ƴ���]��Ө�̾`���\����3li�4���k�
�>/f�����JR�L�Z�2��5�$"�F�;_夨�2�x��o�l�U%�|h7Rm�{�H��V���$��x�wT <���=X(�ۦ]v�*�O0#�V ��˷�s]H�3�V�E�q�T������]g��D��!XR{�]�f"%�&�<�\���ȼ�wV\�8>Ym�C����Vf8L�?�j�;�=C���{
�f�b���BrFU��q��Ηa�Ė�{[��%�[q���i���rk��ի^�b�^B�6Z����#��]-�*5�3�y��ߓ��j���?S�S��s�,��+pF���U�74W`2^����.)���ڵ��E1Z�%B7r�M�������m��ߴ�6_y��R��{��S��e˂�JLu�A�E���xx��d2ϫ%p�$ɐ�S���ؖ���DP7͠����Taz0�(��D�+嵺2勒{���N�W'-��$��d����� ��x�R��1�� E��rQ{�U��=�m���ʒ&�y����.mU�}��P���Vy16\��5CL��	��4��9�V:M����h�0T��K��ћ[K|��b8([+�qi����5T)��	��b�v�S����
�ֲ�ݽ �pH��?ɴ9
O��$���3��i�:h��5sf�"�L����X�+�9�P�+ft9�w�L����=���k$��s��z���2�QWu� Kє�;�uRH3o���ʔk�D�֗��GZ)#Ī�zn	�Nᐷ'^�*�nUk��:����"��5=~���W�c����2?��΀������E}��q�a����5��&߉=� ���(�37j{�='~mcO�Z����*wu�I����&-у<v�z�(�g���`�q� �D���>���Xzyg@���K���5��v�� �esZV7[[z�pm���R(��۱7ps�bX�t�̹�n�@��-���d��cR��@�	?�z���Mx�r��;Qm�~�C����QP����U�+���H��_����z+��lB�#M�xzc�n&!1�C�	؂"�97������|.^�x�N�����!��+���1��Z����=����46��[�L��͐�,�&��6��}�s+��8vyEfK�W�S%V{ئ�Nxd�q6N[�䪀����CTG�HM��2�	Ebm�c�6�I2ضә�z�A��ʖ���R��ߵ����v{9paG��8�
�暐Oj��D+�R[�[ &q��k��ާ�Nw�?�ǽ�#r�2�@�\7.4[KO���y"����P���:苮�b���Fl��_��zg�i�V4-�B<(ٷTc��$�� y�D��ɹ�J�7�(�H�] ��5����CE�nؑwڀ�!jE/9��t�b�냗aoRe9]�{g�'8���1�k��Ƽ��i��[��H�C=��Fp����R�D��k��"��������4��p��2���LP��A����g��ROŭ�7([�ڏ�cg��JahW��9��x�A�~h����e��>]Է��+� D��I�H�k�ï�,��������5���O�`zP���V���źOv�f9#KE_n��걨z>��.!���H����SN�N����0bX2iz����h��:��#��F笲�d�ѭ���l7���/GPj�����0���w^1����A�Jkã�>�����%�+�N��n��1gH��|q1nN�`_g��%����r	MHtgP��z�tqW��s3Gb0�ı�sH�y��kX�$��K��P*(LdS��w9P�&9ElG�/��3]�)��Ϭ�p>>�(�rY��"�cd��@
�"�D��������K��jA:De�Q��SC��O-ĶE���[�TNC ]�Ębd�i�f�s�����h�=n,Gl�
c?���rV������hɍ����:��~K�n��
jۦ=U�� &��1�3,{���s�P!g�'=;Zpf	.{�;Ҙ��tb�H}�bEvHl� u����R�c�^�%���&rS��;����ߪ?�<޺>��~�`���T����x�:�)�ER�����t�15����LIR�ՎTC��-�b����cT���|�Փ�P{eB3�F��s��t�ⷱ	&�K��vnS:K�y�q����55D���lV���7����({*nr�y\q��g ����u���û�r�q����D�f��d���%� LD����FGh��mjY~#��yO��Eb�#|��U^�˄%����p� ��9��62_cr|[(�'a��?c� r��oY\�G������:����֞O'�~cT�)��3�U�)A&��0M�ǵm�o�3c ۬��w��4����L��s�fu�zj� �Yp 
D�к6�����l�u�j粓������Y�jLv,8}R�SB�S�,|��S3 P�iH���8dl?��Fe��Zuٳik�5JO��|Ϙ�m�zaB�B@P3�9��a�x�����e:9:��e[���hXD���N쮓5�c��B�Kn��f�#F�cVR3)�ǹ�s�r-\iu�N�I2���<�M� c1խ�@��b=�۠]r�L#�+�ƹ���b��M	�%7!�g��A�5m�j�U*��Xf/�g��
-���T��N�2k$��s��	�5�'���ו!���݀xi0��iI���@�Dcg���	O��H>(-�3�}����dQو��d�n<	�����.|%���*�PAO�^�Ȋ"n�ϟ�1���Q'w?�I�YvF�Y�n���7�8~�o]�R��aX5�̕�Nçdیy:���C�Z���[��w6���	��a�n�Ů]�U�@���a�Jy�H<B� �i�8���XoW�\�k)OCV�^C�XF����&��5��.d�Zq\��d�tY��5��U���O��o�Z�/K�=�)�}�&&�к�aͷ���3����F�څ#K�g�������Ғp��,�-��e�F&m~j��z��=��m��{��Y�J	޲�( �i�w�U���TA��_�HO{��s������r �h>L-LRU�e+�R����h��;0��l>R�Y)�-���0�:2Y����-ГO���GmU���7&��Vd�
go`A[�iU��Еk}f�ME��Y//Xfd��y���RZ��5/w�1��/�4�|Hd{��r�>�/�=H�� �Aw� wp�r�k-.�����*b���#	/��IX��]Į�U�����G�����=�"�e�s2���_���doE�o����=�qŞ&��\'�r��ȸ�e�N����mo.!���l�&�*6'.��i�����Uc�"�k-,���JɨGpd�8<߻:�o������jME��K���������/��؊�,{eQH/F��lX��jH���}X��d?�C`?�w��T�!F��)k��_�ث��Y���"�֚��Y�o����7Z
6&���b�;�@��u��yt�@7��7�� R�{K~m�����ʇ�	^%��z\5��f%�Ī��&66��ўs�no��ϓ$�֖4��M�������T�i@�����ˏ(�b�?�\�>��hst��x2��/��C��Q��t�-b�� �����x���Ov3�5�C�_u`�N=\�s|C���a}����i����D9N>ۂ��1Y���� ;v�g"�	�Pm(�G�H�+��o����K��
��	V��m����Cq�&���q�<����ɲ\�a��N�OW'��UQ�R^��$w�<)�9%⤨��J$�(�:m�[�m�Xx,Au�V�:z�r��Ӥ�� jO�I��˿�.� F�HYs��>�<5�v�BA���K�A^	7+}`_�d8��Ї�vϐT�]��y��4�b���{r���ĺI�)���c�kH�ưF�*4�-�s��`���9R��iTs�]<�;S��w����B�����:+g.S9�t��o���":�}Pv�󑣨�W2ݝ�q����Ae���A��õ��"[V��b� 0��[2Vri�=�!7�i��k��<fYbL�!��*?����X�yڧe-��ͺ�Q3�����5]I:ag����q£	��Jl�k��ª�ұ\S�}+�.`.��0��[����z�nA�zc9�9�5��9��	��>��oZ'F�����kL�]�ơ�.�-ӳ��v-��K����jq�?�fG���������e�m
�1 pl@���D����L��^�'{O��K�垷�Z=H����5�������M�G%N��! ��hj�G�ka�PE�#��G���$�>kތ�{G.��T�g�I�9��Ĩ�{ȨE�SZ��Y�T���q*	�5�S3�2q鏦�E�ܱdt�1����t&�@\����&;]}-�C��qw}rd��gf^��^,�,Ow�|��t�Xqs	#��4lM0ѩ��˱����֪4��01�cI�_�bĆ�g��~W5�a��w=^;�%���e�Jx�a��}8:K�8� �"�Iw$�g�Bp�y|u|hY���L>=�f�]I/�j0�=2Pl�E��e
��Y��7�in�y��S:S��~�; �[)��r���%��%��cU�c_�g_:xӎ��n��i���RK�?q�x!�;�./��Ŋ�yj�r8�{G�9V�

D���K68��&^�D\	��S�VM{&h�ܔ%vh>�����r�k�i���Ok[/ȷ�K��M@�o�o�n�+c[Y��������V�N�q��ZE�3%��,GIb���y� �mK��wƊ����0�l�e՝-֫�zm�O{�OV_���w��t~�Y����V/_LѰ&��{�ʪp��t�0�`#�X�As%�A��K�~�b��G�?�����0�ݳ�V��琤y@�4֤u�ն�	�
LS��	;�wm�ly�»W�ȃ��>�����%RI�~?�-��Xw��Z#����9���܎�g�Õ6�$�\���r��J��)��S�"4񑱋:�z��rY�gٴ�A�Q�kY�N��Ʋg~i%d��
��xd�O�1(��T�������\��/16���f�U������6���h.w�,�3�d�7E+r��a<,��&
d�U>+�@���k}�ǎB�[�ݏ~,�O48F? �7g-�A�$�L���+�5���˨�,�h���;���d"7��*�g�/ʭz�s�����%�e�ϮYgf���lNa���W]��0��#u# ��~Z���v]���kv����s�	
n�Z��_7 ����m��x�}dx�{ߨ�#q��7�^���5���QS��"�jm�p�Lz)�v�����yR76������X7��j悛�!L'�:/}(}��L�o��Fr�Un�e�����*�3o��m��s�v��R�9`�#`\��%S�d[��}-_��B�	y����L?ђ�}G�쑅#Qm�Wl~�������>��fd-��4o� ���� �߯�:�-^:�Y��|Z�ߜx�%����a��.Y(]��(�WZ���x�>as/�0��U�Hyr���]N�$��9�1�D��� ��(����}r;p(��"Zj�!��НI������;U.�� �c��oԵ<��7��ˁ�Kc����*� є�+)�8��� I�4Bd�\�Φ"g�NH����Q�\Ϯ��@��UI�XZ�j��[�2��Cw|�Q�����GqWtSb�Na�Ȉ��R��߬m��M��D��j�h\ ^���Γ7Ѻ�%�����9erT�' d��n�+8�_��Ӎ�c�efm�����6�%G$%�n%/��:,�ʗNL%%���˻$�b9�@�Fc��v�m�؞�|4�2W�5����'�!���ǠxL�C���k�2�T+!�6�/��+�m=�U��ǥ-ę �=����⌛�y�x�+ɮ�]%��oq��[��4v�Vn�mf���-�ȫĠE�f��J��j���UxgO8�4bs�n�!��u�`H�V�	RM?/����;W��r�mD@����&���>���}�2���Rּ�=0_s4�@qN����?*sڐ"�wq�D(��bz5hG���6r��K�\gM�]�\
k��/Y��;nf	���uH��_p�ɣ�.���5���^|Gt����3�
L�E�}U��BjuI�����"j��!{{��$��~�{/Y<KQ��w���/�U7�E�׮+���Is�j���Zv��
L�%����v��6�DL p����?|RV��sպ��j	Յϡښ�Wy��n�L�d�vt�>`�.A�AB��ɗ����q��Dq��c�!;�������#��ʇ0�t4���\������%�\�	��>:�S���[k��m+ϱ���rɸ��^'��*s_D$55Z��t@m�����"���'��l/|����6 �9�r[]p#�:�k���?b����'p�����pᵵ��5�j�M�E�G���Q���4�?ܫC
���CZ�������,LP��Z�=��VqDg�A�\��̳Xݎ�&�`kn�@~�y��r"���S��O��Q�LǱ���QѫľU�g )f�c��^�e�X- ($=-s��E��x!�8��B=߾Ѱ�:U. �=�6�Dj5!�����pI��d\+��j��v$��pc�Y�<EB|8�U�u��:/y�]�GQ��L����;QS~��Rb���|ԗ� �28���t
Q��Eܓ��+���)���C1	�6���M��{���`�gA����X��ج�yl�\=� ����l�$:�4��δ'��
,����'գ����|,�CG\�U�=��f-8�7D�!�]�I4~�l��G�A�c�Gϝ��X���|F٘��$�ߟ��Ȁ�R^�'�Y����
גf��D]�3ߚ�7s�%:tעX�@-�2�sO�K�O����&��3�?��_:=��p?���^���G�\��?A�8��P�L���qi�k�D��/E�#,��{Y&!�E�a�lqW'��v� ���2�;��:�F�o�ް���P���z�o5M��Q�h�bQ�d/�^Dc��|�bƑ�H}8mD&�&�ySd�Y0����0�D?f�>�Ȱ8YTN�-���*���T.�\�[8���9+��ۥ�lbJ�;I����!��>Q�����)�⣖R�����@���j��Tn����C/B�N�y�j��k?_�Ө��M�Z���� �R�2�*�S��K�T���+rP;�u�8Nj �3�K3q׵�O#���bi��Y��V��oBmf`�a���7Kw䶧.�2������p���-�M�&�5B1g���3~���n��7�����}<Q�}r�Z'�L��d��d�2e�_�3������LXN|��u��KB�M�3�6�1�	&���xO�
�o��D���|aҪ\J����`���g�zH�W��Q����@�G���h��0Փr����r����So��HLKb͡ȹ:M�4ބp9�@��7l-����ra�6��=�e�ɓ?QX��1Ü�Z��,�-�Zﾼ�J(�[����XQ�3�)����#�c%v���A� �_��k��AyFo7,�*C
I�F蘵h��rV�/�<�Ʋ�ĒW:=SL.(w���|���(D�@\�}n��j#�E��x9� %�I�9%�InR�Q}wQ��i�:M0����aD��`�{I��&iTN���z�e�c� L�����~N�.$��>����;��`Q�mO�xP��ʙ�Oa���!����~ "�2�x��r# �C�*-�=�D����<u�qGmz���Ţ��Q�>�֓�ԅ�v��,Luy���;JcȺ���_�A�jtն6ޜ���$�������>�H�X�maj>���/��@)a�|~����f���K��g�}�!Vk�ЎK"(Q�0K kV!�"VT�!��Q�AcS�V���p	#�v#[���Hb�����j�j���\�Q� Ђxņ ������q���8����]�3��A���Q�6�A~�Cs�*cy�`ݶ��/��N������(Y�� �>��0xA��PE���y��h k�B������'�;L���aKbĉDrP��er�h\λ�!�����ͮ����upi����R� Xw*��r(�;$8f-����c�31ݭU��	��� �u/����}W�	Ж�g��2M�#���8/���Dgb�x�}��7���R�RT�&BO�l�W9s;=���o!҇���[����u䚼�<��sI/ļ�w@D/W�W��(��G�G2ă���/�kzJݪm��{
w�숪�5"�L�U)<6)�bE��U ��
�H[];�-b�6* �N���[��H>v�N���Y ����ƾ��<���z�q�?��6�%�6����p�5a���19��)��L~C��a��_^�c���.��o=�7UG�� ��41R�j��>w6Vw`"X++n_/^3a��[�i�ݜb���Y��?0�xS��t0�I[��u�����-m=84#����5=$`"�
�\|�J3��i�Fi��^w�p����;��r}�4r@�`QK���Wz�}�k�_q��o�}~�ty���wAOHnS�ϕ���.��\� �����v]h�(�\R��p��!�.�@��@,�����x�s;y�%�_�$&�T���ᚷ��e(�T��X�@8�f����tU��u���N'b��v�]��z���`y)߳}L�K۾�GXC����*8U�Co���������j�3G���5�$Dux"��D/��
�=����
�]nVem�Rjv��ߖ�O*x��1��"H��RZG
��XY%���G�|��(2�P%!8�[��ޘz����2*Ծ2{�)KňcG�>E�^��[��1�r1��g�P���Q���G��Bjpk~��GPJ���n;���q�?DZ��������j�êt(}*e�3��2 �=�r���:��M�meƦ;l�2�~N��8��H�ia�b�u'm(t���z�NHe��Q���I�tt�0��V�B�ERv~�T*�����on�At���6&�XZ�KR����,ot�|�������D6���x����/Aꚾ�w��9g�;⠦��a���t��	}�ۙ]Z��^��a�M�����'�9����q�^��l��bXU4F+�L�E:rpr�P��do|�9�!q�v�6�+>S��$�2���)��E����?������ ��,�����S6���]����"�ٮ*��>[	o����s��5���U�9\q�Ԡg�>��,�1�A@�����(�#��΂gٍ����M�s�Q�5�l�(h��x\l���������!��+����H�{��}��t�u���|}�]���F�Ym���s�ݥ�*^ߴ	@? ��,@��J�fj��0�Ӄ��d���8��qB-���ژ��g�C���W��	�����n{ �ɠ@%BX���7�a�6��1�g6f�O�]2�m��<�}�S����T����>��a;��G�����s��.�]s�a�$U֡E�WR#;�`�����7 ��li|�g�a�V�;Lm9Q�b�;�o�9-�cRUe��^ ����	/&"(�9m��8���=��[e��塼��򺨵��P�M�R��
�� /��C?}W�*�*�����IV�<�!�QSK�+���h�0ެ!��SF����p<�V�!h/R������iV��_/���f,��<�xj�
�Q$��E\���8g�s��VC1�D�l��Ct2�/-�_��P2�Y��[̈́�+�lO\���ڑl����-��Sj�â�ҡ7�;���U�?��Gш�����"��UPc=�,5���[�.����}m~ ,j.��`�@��]>Q��Պ�0�,��;��xb҄PB��"��b��u���~H�@��V��j�]q4&"�u|'*�OԋG��� ��AQl�J��\m���r�� �����,���l�qz��&Di���U�=k�4j����F������I:�mo��]�	_w"���gOc7���~]�T��ř?�M*�%�EfW�s@�p��	�[r�T����46���)c�B�d30~ Ո��z��ZĘ���=`kg�<������E>$KC�|6��޵��� ��**�Ю�6��m��<T���s1�'�y��)//��
�I�N&����u[�;�����g��g!��Ɋ'T�h	G� id��,XL�Y�h��x��o�WΟ���![Μ.�����,��'��
�@ݧ.н�Cpن��{���Z[�Įd#���7ĉJ�kۡ�q��T�����E�WK^h��/T�<���;�;��Z��q�(V���a9*��H����V��[� ���<]V���p��l��|���&̂�.��9l?o�VbT��Yb<:E�)����o�8=��'0�̯&g�@`��؄��n��e�ubۦ���C�{x'���E�֮���T�Ɖ�3�eLn��R��b�zU�j#FF�U�� K�l�`�@�ȥ��Vgk��<J�ٶ��֑p㡕��UZ�^Ϗkx�#y'�k��j����:���c�f����l��/%.t��{��r!�i�N�/������0Q���Z��bԖ�Y.�>�A��QWαr���;ۑW[W)��{���-��������X�aYB��R0�X���c���o�\��J��n�iӿ_�S9�aԠ��?s �{�)��UH���U��w~���rH�2͂p�q��!�t�B-�6B ؊�lYq�>X1q=�N���?�7|��2��(V���C@EE�hR7?��Qk��L��N��;Í��W�9N0(7��lE���
q�ۘ�ڗ���K�|2��G2���3��uE��Ƙ�	�t�*`J��r�,��yUk����[�X�,5h��hSt����r�D�bC����ԏA�~�c�7��IY ɜ�L?񹞒��g5�6��>*��� �M�K�cmߎ߲��ƙ�� �=���({�R8>į�h��k%:[�����W\�P�5U)^�m�kpT2��,���FO�L�jOq@��W�~����Sǿ�����?F�D�_�y,qޒ,Ƚf ����9�����Ǆ��
tɬs�C,��$���1I-���[h9���e?'���b���ʂˬ�����"�q��f<���9tR��-�БJ��лH��t&�(\E�c��3�ҹ'4m�`%����g�l`v�xh��4/"��E�B&����W��&y\�j_��oK���V=�q��,����lTArO^�@õɃLr-�6"z���);1p4\�������c�)�}%��0w��~!���r9�A�Ip�*�.%+��{U��s(�@4\;z�i@��{4U�w@{�ޔd�7���}m0���X��XUDkp��&�/XP�NR��n��ţ��ye;���6$uT�#A٫��#}ep\��)�5\���c���T�]LF�mlT>c��>��f��h	H���Bݭo�SE_Z�*�d�'��L&���0��<´a��+��2���Τ�Y��i�['"B���Vו��=�
iiz&%X��؄����Ҥ�Ct��ÑDo��Cq܊l�Yy��<9k��k����De�� ��ߥض�e���Q(mǠ�V�a5�j3����ũ�<��M�v���؉�}Z��[���Ha��ڽ�ӑ�#FiT�4�q�GE�������@�̈́��>������9��"3h�p�Ɲ�0Y*[/����#$,Zk���L������E�)SV�F�W��`���0��]���E����0����1�n��Ѻ�::�st)Ϥ��9YSūN�%��2~��r'7����`�J���z�q���F>��J�t�s�G���Q؛�$��5^�����0�����]_@ב�Nt��8���f�p=$��E�8��ȗ�2
'/Q��}��$��P�����C������M�J�{Jrw�RV�p��-ќ�Z�@3e�s��S����-9�a�rY=K�.X1��[���C�1m��U���a<�]�Zs�Yb�v��Sc�`���V��)x�wJ���~�"9T���M]�������J�d�ͳ�b��Ǔ�N]Tn^�V�e�4�J�����{-��[	�6���w�8�ӧ˛;�!C�T�f��!��:[�"lZ'�q�UB9����,9��iҎ��|qoe���kG6�'a�_�Z�a����qp�a.��s=��
��I��	H��[��%����O����L/qXc[�W�hc
6d����b?u=k3mv+J�*�&/��'�ƌ����5.6�#��Ll�Kn�KHv�&(�+������*@p�VN
���~\ZN�"�$}@RC�W��Ӫ�B��qT�{���Vb2c. =�W^�,&�^8��q�#t�!c���#��i[��O���|��oTe%�,L�ih��d��ͤ����1c����(j���MI�aTh�ym�g��#��� o�oM+�X-1���~�;�{��y���#�[���2}=����c|�v�X����9J��ض�� uQ9��\�(��b���ܔ|+~��x���r(#Ʃ�%wW��H|V���Tkk�,��=��|��F[�!S��6\�ipx�� `�^��'�i�r�_��π���۷�w,uGG_�{RMxFJC[乾4/))G�$���m8��r����xR��D�(e�VD:$P�Q�匳XN�r6uHYfT7EW��/��;����}�"��(~6�=���],`f��緙�|=".r'p��ѡ �z����5T/��M�iYk�M����l�9�p�7b1���n�0�{�UB��\�<�u�;����B"Vf�h�͎H\n<����y�O��߼�/� y&�X��j_c7�K�23�'��8Y�~�4D�dJ��2`�[S�dpX琟^��(�K�����w�������MB�N��B&�l@ �ϛ��Bڗ����[�2D���u�붾�<dn�sm�Ġ���m0Gȍ4�(ڝ�Z5\�X��̸��yYT��5�Py}�È:ޜ��E7��<�����O,�p�A�W�v"��ź_$*^�';�t�r}�tሎ}��UbY}R6W(��6�L7�գR�l#5�ڪIbجKT�a�m�����Ҕ�ꈟ����Á/�&W��Ё!k?U�3Z���
��&�R�{ur�C�̊w����h�𵬙*����3C�N���IsF
�l��Q��N��D� J~{î�a��tN�-3���@�a'�l��^�u� ��x|CCj�) jj��^���j�nRK���D��t���U�����II��)(�	��)By,&2�{�FQ�}���#\�t9���`��3�6�B(C+{�~��[��a�#��z���+-�[o�4.i��ڈ�Nպ���=��wC|�^��֐|��b`
�������Щ�3=��Y�O�e���Q�D_��c��3��2�����U�D2���V���w�d7���Z�2{�ȥ`��葊mV��l�+�d����O���Ey�\����lr8�O��u-dљ�ґI8���0E�b`�ZǙ�j	B��u�Ƕj!z���㈬y�+Z�Ɲ����pcc�^�?�𼦫���2\kŌ�8�B�w�¢-X4���!븈B��e�>�n�h��F�?�\���l�#����W�^ZB"H��Z�d���3�q�^:ɹ�u=�3�1�Z�/�r�$Ő�G�3���N�2[����S�}pc@&���+ڿ�gZ�-#hn+�i������^-C"���G��Nz�:�Tg7=a�����8�9���F(�a�9r�#�����䍺=VJ#�Pq�R����nJ�W��e}ǖ5>�q��F�rxİ����
O�e~b��m׌��:�j����;�g)��� ��D��5���9PwtK6���}�6���L�vm=���͇c����>L6[���s��o�z$��#�N
�a�"����Inc��zH�wT�]Ph3�k#�{��/	֭��p2��� �KJ#�V:��y^�u�a����4� }l-Q�9y�����5w�2��(C<g0f�3�������
�oZ V��MD�2+x�c��t�Ur1~_Зj�i�Y��B躁��b�����U��c�xl�P��C�.~6����)��&�&�����EC#�4� ��S�0��,S`�в� �O�D�m�˰�7��J�)����5�	\l�#��l_���_��*O�**��5Iۀ��k�{h�O�v�':���M'B|/���F�[lC(Q�*���TQ,ꈅ?wA�2Y}{�xĠd�;i��5� <ހr��C����>K�L1��vL��/%��3L�w2�tWKN�'ԑ��N�Ҍ)��~8/�������F;��>v�D��x0�V���yb�� �n��Dx_�sd��Mr�Ί%)�o퟾5�-S���ʮwX:y�bTV;`��>�1�\҂xՎ����ek��s H�X�Ĕ�1�bo�f`�<0l��D�u��-��������	<��?�EZ� Fy���Ģ�{A�8��8�O��>uB[�`A�w�7���K���]��̾Sō���@��!����
�r�5��|�Q�N��G��÷�v��ux6Z��n|t>,� �?��	�W�@��Im���F����l�b	�b��kS�ڿʥ���[P�\���̿	Y�S��˔2�7V��ܠc\j�2��>��<G�[5|Z<�AŌ��C�B~��x�m��8�	�r�/�KNr��.2N�݋�[�����ň�p�ܲx�0�Y��θ
������<E��ι��>�΋�o+�(w�J�be ��X-(���"dz҉%��0�-�Z���0�����٪1��X�!}�ȸ"%��h�6�㞭f��W;����N�{j:UC�X�<�e ;z��4_+�ƞXR�O1"\<�_��ZM�P&)�OҸ�a��c-ӫ�qU���S匱��6:��z��,��z B�������b1���Q㵊2ep���NM�l����(���Ӕ�!����8�J�E-�-in �^���N�Q������dE��=d��R{	C�n��)J����6ؙ��@�P�M�^�`�C�aAP.�7v+��f-�����K��f���!�~�@���,'A�J���y��$#*���b\���:񂊤~ߝ6$�J�\x�ʁ��%���"(�[��&�)�l�!m!����j�n�#h��<��ۅؼ;>�a1}��ب���'A2 �*rH"S�	��|:�MY�4�%��Ʌ�ԙ,����	V���&DZs&�ꅭ�F>�:���r�f�d��A��dT삦E����g��0�Z��I��R�I���L���+��M�Θ��a[�0���Uhǎ��կ�.�s=�������B�3�["�D#�F��Td�/��7��d�V2�Y�L��wa�
����lG�����C+�R��/j�T���KjF?��7�1.�2LD]�|:��e	}�Ϟ�?r��C��pF8��M��솣zQ�py�c�v���.h6fk&�d����M}�+�Ib��q����)\O�_=;w�f���G7h����	N�w�6�����#W}�teC܆P��n"_ϳ�b~8J�ǃ;����}YA���R�Or0i��l�'��<J�d�xz� 6��b���#�R87n�������"U�ST ��|�/�2��E��_�{#.���vW2��E��۰�w�x[�E-0"!�9�	��L6�dA�k�&��cs[��;�VT(��ُ�K��B�"��?^4?�خ�����ʌ�q��a4�(�� �á�柏D�#��S���~m+���#3�s�tŲ�w��������'!�+hH8X�֜��$��X]S��1@;�N9��Bq*޸��.G�>e�PW���b����E�����@ٲ���K�L�i"Ki�C���U�It���W�r���j/���t �g�[oQ����D�ͩy<uD�?��;���צ��`́P��'`k'ý�|�C�iYΤ��P[@�P��^9W��/c1��,E��7B���K�P�6�,�3�Br�*^�LD��y��Tتi�[�U��X���-dR�D��F����13j��R����:�JZ���Ż�J�7qm�4��kr�yqi4��ZF|�7@_�<��y&G��m��M��|i�,y1z��t0�X��3�H���U_jk��@4d,�����Ū:()i��%a���i�G���l��2ܲ-�I����mA
bL�-ީjڬN�����ݾ��T*za1��e$}=V�H�c��0��p�e��69�4V�@#u��1<��ɦ�V5��Obg?���P���$[�/sa8i���Z��1t\�Oig���A���6ޏ�4%R}�"��Xa-�� ���+�:�׭��=���ė�����7��=7�1��Rv�y����
�X���-!9��tGfWC\�#Į�}:��q�P{m�.��D�b����pJ�Z�]�J�����q%�P��� ��bs��5�����`og��b�7@�C|�����������% ��ͥ��,!J�B����'A?Zb�G�!ɒ$=�]Z!p��e��=���xX�b��N�vT*��]��[/�0�k�6�6����5s�R��	Pqw�IS��������A�V��8byEcp�
h��U�Aw&��}-��8�~�������$a�Sd�'-���¨י�*m�V/�����-t�ty �uG�4a�=��+��}�'7�F�S�I!�]h~�by-�5�dJ��C�Uo�-�I9���x�"$�ܸ:��������r�G?�]�^G�j5>���T%H'��*�_�q��ߩ�G��ޙ��ޱ�QV�aѯ&�~�B���m��	N�A���H��vϧ�P�;�YlI�v���b�zf��Fto�8�|s2&J1)'`Q�Dͭa�����="}�`H������~v�nE�E�[�:rF)�Sq����7𾦝L��ܽ�>�/>���c8)�0��Yw�wZ�N/*!��X���ZE��=�H�M�1q��"V��)%+�[tw��,{>|Il){K�
��(����V日��!�����%�xw���?�,�դyUԏAU	�YTJ��d:qxV���D+�����s��uf'�G��Py>�Z��� ^5DoMV��g�.��/;/
*�8��@�M�|3z��R��L��D"�_�l�������v��r�����l���>r�$��7��5r8е%��L�R{|��|�h�I���0VK��>ʹ�(��>t���(E%��=�
���2�2^��]f����ͮ_�gg�3�$2����{ K1����?3�
S~�>"�-���a���,�&R1�E7d6b=`�w�ɖ���"�0[��Q��6���0���Da9L�VƠ缥���������:A�q�S0��M�kx��bf_��3������9ϔ��b-n$`��P셤���v��U�	��4�LɝKFB���%�5&P���J�d�'�_�`q_�Ֆyeк�We�n�`#)�`��ɽ CK�� 7�����7�d�tgI|ϵ��Q~hoo�C�W�j�Y2��>���C�� �A�Y����!�n�I��R/K8�"C|톚�8Sq�Xj�XU��VU��D�����c�7#C���穈*��^�8���N,q�돒�{ғϚ��M��R��Z+Q��}��{#����v��
t��p7��i�,d�0jC UR�g��@�U!��ވ��]�W<<�����ų�eAF���Vm���m�~ܪ��݆����+E�!�ato�4�xSEdg�}��D���)h�ǘ�\�����c��b������^�����]6�� ���P�g9_��\��߾��i��4�U)y~|O��@�VJS�-� ��癖������i4,�[*X����հ	xln%M��8���{G��]��ʸ�z�������E�E0�X'87�6�u&�gJDIK@��S\0���th�Ǎ,�?�QK7�����q%��?R2�:��"D>��q�;�D�m^�=�:#SX��m�7�<N��i�?	㡧gh��is �i����j��gv����6Xs��� �[�7�*�F�	n��i���>aܫ��b���EjO��n��B����\���XG[O�y���`�����/>�K���������b��u������R�_\z���B�5��}�Ӓz�����^ґuO8,DvB+U�N�����v	.Xe��fa��^�x��l
J�b,Pi?�9�o� K������`U=H՝��"S�W��d�%��',<�u���c\���k	6�h�͸O��ШV|v\�{d�X�$�{d4�<YÝ��~�)�PqH�Td��� fV%�uiÝ��s���o¶2�P>�J(vѪ�[���=��z�fg=�9�yt�� lऻ׿%ҍ}ɮ������,'���pi�����������x�5��{;s`�׵���!���M��0]��x���:1@DxN�&���8	F����ϧ9Z��P����y9F0KH8<��	�ȈH8<bs�>��"	J�q��,���M[�W��"4����꫙aؾ�j�0��q��k ���ʇ��}�l3a)��ksF�)0���qw=�l]���}z��eA������ ���ֹ1>����{7z��d�[��w���7IE8���o|�W�N7j��=o�;?���Y;4�&�����̘2�EN%F�iC8��a�T��͎<v�4�铰�c��d7a�!�P������?+ȋO�;;((]��_5�%��)��DdfհS�~bd��1�mB<��㊩F����?W����Pp���R��t�QG'�٨eK�HR$��W�[�s�$�0��g �uf*B��C�	=�Q>�4o�K�OL{&�� ���Uw�MGR~?�[���m�Kv�H"Ju枌����9U:d��>`��$]n--��"��I/R\�`��������UB��c/�"�pa������Q��͕ �B����'��\*�5uϏ�F���{�*�Xw����w:��/��Ш�)w����	�(����Ϊ`�fa{4���!��T����$���H�`Z��J�9	ⵍ6f6A��������fg���-iU/�ē�#��6[�W���\P�&9��2�m;s�ώ,?�%�q�&�gD0-�\���F��.�ߧ�\̚a9���/]-��Y�X���6R��=�/�Z�h�!ݣ�-N�5ɶs�"�� ����H�J�v��>*<U��>��F����p�檠.\O�^bP���[�7k��"��α�� 4:�'�MZ���.�N�#�u��n ����W����`��+�f��4��?_nO@?�U���b%��FxA)$���x8�;q�K:�����()X*v�W��:�6��#�0�R�p�����j	;#��4=ܙ��n�ؖ����-t)�	�/�u��m�a2zx�]LAX�%{Aۖ�k��r�i�Ws��Ov��V63*C�]d"���{��m0��K����<%���`���O���7�%�I�6GGԮDIX �OK�ġ�Jw�ը=T��-���]� "��6x}A�{��wY��t#x1���"w����E�ZP��6��q��!Kd_�7,�Q]�i2 mW�
�%U��'Ϊ��R~~�������/�ŀ��瑋�()�.�����qO��z^[�Xħ)}h깝+$�[��?)�h|ސ�}d8�T�5@K�M�`�'�/OuG֐��J9U��0���)�9�O�-[�B�.g�������R��Q}�n�&��Z�a��n!��_�=��+��C�����ii�Bg��y)�^�;i��*���RϦ����e��$3��Qܐ~H܀�J6������m����-���з�E)be�02i�r�L���av�&�Or���r�d� �:���r��WP�M�9�;�,9y8O���k=�$R������p�+�(�p/3�ŸWu>'L�o��Z���\�O&��<Rȿ�L�6�R؞��و��M��������L�W0�Jy�}�!�Y��֋�L8��(�`�=�c�gC态�GW���~�X(�dIj�Y8.�ы�S�n*{%�XS��3��Y���.mfuхNBL��Y�S�)$�n"�Q�a�i�h�#b��h�D��ŷ���~�v�k�^ƥ0��]�����o���<��
���$+(���\X��᳌�g�g�Gh� ���<�����Ғ3[y&��"��Zj���U��遞���U�x� /y[��J�|Ŧ��s�}R�2��2D�!��ʴm{�|�C�� �B�$m����FI���q�+�����4(���y�2�K���΍�y����R�{�k=8`|gZ�r2�)�����C�m���V����y_�6���mnS�'SW`8<}x���0وg�	ә�^�;�Ig�1_]1��dc�u���m���8K�������|�0:�d*�c|���q=��L�5	�MYq�0��8�T�V��-��O�7ϳ���4��zZV�� ��6�I*�R�9x��ь<S���Ԧ�n�]���WG���G� �5���,��E�/�g�ܖG"\Y(.f�"�����#��[��:j���ד�W9=��lkA������J��?hfrϒ�-�Ϣ}��3�����k3pb��]�;['��F�Υ�)�$�8�����X�~_k�)��� ���MMB�q���F)R��SP�ht��V���W��rtK����R
��\�se��q��zQ邥�5u�D�6TMxb�|Y��sk����w�=yKt�*{2j.��΀Ȧpk�j@��i\�x�?~u�g��o�`�[�˃'b�)�dӘ^��n�g%�#����BL����X"p^�YS�h������ ���S'�a7�\��R>7�B�	~�Ft�kV��^��%�2��\y"���d6va�zȌ��B-��&��w���9������K��D�Zy�N���� �q-���2܁��'Gx�4�xN�?�Y(� ;����xi���?���+��z*5�'g�lmS���C����˵�$�W[���&�O1=����赃����I�EN�@_7^Pm~��
�'l�y�	q�gO���n��������/��x�¨��~�.;鸞����!Bq����!#��&�U//n�#T}Z��_�iJ)�;��'��S��K��O~�9��Dv�&��\`����S����*�V���̺tɜ#�ޡ,�1l�����l�`ͣg��[�g��T�F� �����_}�s�o�#����+�R�H���i����ʹ�t���v�0��v�"���QwM7��V<%R�# ��n{�9��Y�g����VT$�X���r�よD/�|+=gۡ�Vf�>}��T"�>To-�����!na�Ya=�$�.�踲�a#'�m����h8�����D�B&L�Bk���4v�2C��C_;�Q�t뫁��9�ה���&�Vhg=��.���p��K��涊�Ix(9_�6�&���p��o.M�k������6��.u��Px?�S���ߛ�S�������$�J���G��'F~����Kj�� �S���}ך��m�-�d��=Zk+�Mh�j�%����j��vX��r�Tk���-`��
�>Q1��TP�j`So��N��*�_	I ��۾�N^���$��i���*UJvx�h�m����/Q�sK�2O�,���z�D�S���ީ���j�U�>��^���)�&&3�+�5V�B����G�? Z�Z�Z�@f�"׀�볏�LM"�F����XʎGRY���'�H�im�zO:�'���v��b�13�" ��J$�J�s�tG�R�n�߽��$��t흱�*�ր�$����ӵ⃸x�C��0+��>���t���Q��l ���bT�e�f�!�
���=��WP��1��3J�q`��v6�x۽�{��
������'� �^�2��c��H`./%���ʄ	b������{�̑S�:K
�f����/��_��[$���P�0(�~�H]ނ�D7��v�BE�tI$_�ZvM�����[X��Kz8��byA�)�N��@s_��L�Բq�F���{?�MY5��^�:TK�@si���gz����!���;���쓝Ȑ��u:�a^� Va���eM!��ҕ����WY~�Eh�cV�Ȓ�����r"y����h�%�3�R�Rn}��`>�Yt恐�,ڵ��8�zj��RQ�ūc�>�b�e�7�]�q��$��a'>�^Y7�F���)�������i�5w��A�aR��HߎyoC��`��}�4f�KtEUL�S�݈���E��o���M��F�UT��I~cF���<Qo��+���!���������W8J��Q)�Q�8�f��UJj��Ƶ=��$L��uD���S��u���8�Sl�i�%f���?:[b�QĪG�MN�=Iέ0�#�������ma��5ą�)?���0��6Ґ�(HUy<�F�c��4��Ku�ۈ5u)��Ȕt��FlC���I�B:g���O��}6a��RƆ��:��S_�>�9�����瀻�Rz��
�er�<��o$��AW"��ò�gz���+��x�b��D7�"��Á�[��r�d�=�c�6ug��a�M�`�\@�AҌu1�1�V�s���f���0��H�_���֍}%.,L���Lה4�J����k��'�4�M�	l;�"<vj%rp�x� ��d�2%����Ap��m�{x�G�3� ���_&�����q�n�g '�����,����c�՞�oJq1ϙ��������r��[�-Y؟��_��,��FJ(Y$�ڛ_]��b���3�]��x�!�hJ `@#�Q~'h�$s�r��A�AY̪WJ��]c^��X��O`!l�u��1'_� ~9EG�����ͱ��P�1��4�v���1K�]��%��`��跧��FI��BK��
���S֋:&7�XJ�d؀?��[��P���T�}/��F�)[d�\=]�����e�u���8�|����̙3}��l�9f/��C]G(���v���5�v� ���y��*v�t&�ͽ4J��k�N�>�ӊ���#��8Q��U�� ��&�BV�{��w�5����g�������@��Xq��ŀ�p��J���'��du#�^����D��~Of5JU�DX�q6a;:@a��^��`�S��n�/�-��)��Rr��eDG�خ����sTu���FyB���<��R��ȺEn�f>��� �`�dU���*���S�2���ϕ�����O�:��?�G�P�r=����G$���WJm��0tYĴ��6V�uG��;b�,��}���]�W�?4'c��yR#t�d��K�-��xj;������gC^5=���5��3���޻���>�~\d*g��!�c��� 7�0̧EaX�k��p�`c�M���3'=Gձ_�;m�/�=�J������S΄�"�i�X?4W n�����<�'�+L���*���b�1З_��Yݱ`)�W�~g�B�ꜥ��M^�k�K����Z�l���$1����b� f���8#e�`�{�
�"�(�`'Jl��*�И�c��I��-�I�`�{�zBѬi)�'(�j��&F[͏�:���4 ����@!w��3�S��ĦJ��/�)@��NAԄ���}�~4#l�L�g?|�E�̒%�E����W���m�ԚJ���`2^h{Sq����m}��UƏP�a�0�j�J�cI*�8����[��9���r�pb�]�~>����M�	�:�,X*�#,�p�G~խ�?�RV �����a��f�cf�ھz�;2Zd#�gX�0N�e�����y�U>0ِ\��Q�=��ڕ�o�^�v���:�Hls,7LA�c��RRL�z4��e*�w��ȋ�������ʙ��/5B=��vf=!*��B@�$k��'��`^�s�l���*H2�d�)��]���<�;b��?t1ZltD Џ����}T��j��wg�s�:;��6;Ι��`�1��(/(m��Ī����U^7jum��eEO[�7������űI]��d�&���e"����|����鑆�m��&�FN���x.s���ъ�տHT{�E��na�
{�4Iĭ:UK��)�3�d��'��>Z�|?=<�F-+	w�.��-e*wQJb�>�\s�B*�7e��bBxU�a����:�I&@Rtzz���ރѨ��$ٍD�`�� y���,$��b��9<�g3��v-�c�y�kß���t�{�����ol���n������b���	��3ցH�몷�ތ��w� ��������l�C:@M��ca�p���U�'�W`��J5Tף�89��^��f]�C�!��ࣟfO��T�/܈��F�bL]��z�wt�c�=�-�Ku��յ)崶�S%�c7nvYB<����v���)����u)O�2Er�����*ޒdn
d���3����jA'i�Vs��Umւ?���풼��ΰ +pᵌ�dx�M�,��q��q\@ʘ���!��97V�G��L�C���ܢ4��n��خ�f�qf�u�s��PT��>e�P����<�Z�1�;!��2\��^�/���c��[��J �F�	��"Ue��"=�P'�ý�ݐRE��'_���ه'J�Hj�T���&�o	��������ZH��PU�I�'�6hUkY�/�)���A�C�)F��
d��YHR��j*A����\��ϯj��mUt��@�A�Z:O����n��/����࿉T;��5A{6.Lϐ��-9h��#�q��ң�L<�~U!Ӣ�#H��T���9�_������y�&KF�e�h2Zx�<g��~����W�j5�z�#��a�/����8�:dС����eO'dJ�j�(�Ob��(8��S�A��:�{�qx�I��e+�8�h!s0�K�L��I*��5���K~�����Vlr�n1}�4um8��@ㄷ�������n:�s_�ѡ�����G��1���������F$y^N�`{z�d�<�Q}��O½+ғ�b���"6�ML�O_>��g�f�s�.�-���I�GxF8�aH�2TRr�1s@	E�#u0@A">�s|K�=��a��}瓨Z��յX�g��[&@B����+��&��v�998#�O�t�Ӆ��ά���&c�O���~�O��dP�1�4����ҿ�?Q<Pi�!3ma̸*>���@����>��o�y�?��t\&�[�<;��'L6�@�}���B:��;T�?O0&ȫ��Tpkw�q)�:��|��&n�����ݞZ��]��� ]?f{��x\N�Ƨ��W-���f�a�30>ee�8e��-#+�ҕ�Ӛ�z�����l��6rN%�� g7Ƞz���L\GB�&��V}B�o?Ԏ]l��LPLʌ���C�	�]�Šp!诎��̯�y�	���\�2���w�N<��[s��,r��?ƌ���g��������-s|�ͽ�����x_��$��o��IA>tdL?hi�~ ;����j��������,�2��4��GݢVwI���SWK���넍�h�����fC)�=�5���U�V�}������Ś�د5y djT��E��H�(Ӧf'{��F���M|{������>s2D�%�U�p�\Y��P#�֫����/(�Ɂ7�O<L5񕞥�ߋ:�E�<�����:k�%�KY�2���� v�B��gI˨�ƚW�z��_��H돪5����E�ً��GWO=oLM"�&D��74R$�H��U;̷���~aK"u��Y�_[�P��)���h	e�G4?_��|H���4H ;:x�p�v���sY!�l�حT%<J��Mr���u�!9�X˭�����`y���(�C�܃MƼR]W4�ށ�����ñ�7���/Y�v����{�Պ�14�{�d,��.�՚���a�EĤ��B�[ 0̇A����Y���o]j�8�O���Ȑ!*��!uյ��n"XG�y	w87x���(��!
�\7^Ö�"��ŝ͛�0��f��q,fҋA����SDë��40;�h�]��B'��wؔ��(W�}w����'�5e��&Q�4�a
�ز@�}CZ2���>$m�ƛԢ|g��G+d�%�����ҥY�+t��;f��q������k���Rq���Yj�yՂ6���Ŧ��7�/���O��*]W���_]4���E��
���r/�u�/�0��/��"������)�]�7��J���s���u��챹��5S(#iyv����6�&H��,wT������n .�nr/vkbZ�L0o�S�]Xƞ\���N2^���X�ىRZt@��j,��feʏS��&J>`�O}5r���&ۇ:Qg"é�a�mb�;߅<DAJ�v�S����m�N]
�15�6���}�B���P�W�$����h*�{��vrV�q;}"	~M ����FQ9����7�J�^��C>��J��Pμ��" �lN#7J�<�E7��h%%�BNs�EJ7���<���9ֶ�es!_�g������^�jY���� -� �i�R���$9ԑ�W$½�`l�������>���I��D��gōr&v�LNY�Ũ�JT�CT�Cr�Y'�w�:/ ���j���A�/95��P(�aW��TbJߩ�B�����nq�%E4��Ҍ8,&		�XRC(�N��o���#�Ж�^a�(2Y�P����5\�n����]?����Bm|`����0|?P���*Q��}����m�x�P�g1���d �{C�-a��R�5LA�;{.4���V��N�u	ld����1eD��l��U'ix�0L�N}�9� "�x�t��a��>��]r�SҪ� (���A��1�d\FRj*�`deSaI�-w�~�a��E�JA��o�;�Z{~)=��i�~�j�{�iTA��Fy���9��P��YΕ�s�W`�d�d,��'��7\���k�9�)����Nɞc�ή鱋�B�)��S��p��:۞v�
lRH�#��Bn��"���ɕSvA�O�I�/$Ҧ��2{�v��8s&a7���{�Qo�/�Iɡ�oΜ9�͈T�F�Ɂ�����|)�;��ؙ:�����)�+�+*
�����+�u�:�wT�	���9x͠�t߹��hUV?����m\"�U
.ׯ�T!/��[�e��h"715�gDבMS�aD89��� ]8��?�D[E�`��u�-H���p���2�z�mO��y´�G�8�	����ɺ�h���60@��H�.�i/�%j7��>V��%f�'J�L4
��<Sc_Z�Ú)��Jɲ�j���id��&���o�����i�Iu���>\P��B��\)��\z��B�.��D�r����h�7�1D��4���+9ճ���#�R�'�8'��ˌ_��= .t�Ծ�XDFt����žG��bj�	6d�Qw�8z�+�&G��/(�ӶJ�h�[�mfǙ�Z1��5��冂N��j��a#0�k�Y�<vRb�̩Z�_w��ZIGG��w�-Nߏe~|2`���p^�yM�we+�$
���/���h�Wa�G(E�"�8�c�Cw�'�KϾɄ�ka�b~�sh�/*�f��7�&d|�Sa��TO�ϵҒ��eՊ�������8�g������ ӹ`i��I~8�q��;��Q_�OL�<���q��	�O�G���pk=���$�Z���ǼѶ��5����8��|}ZY��]��h���q�>N\���L$P�o����B��65�Ѹ�BUwN=s��f�_;IZsQ�*2�l�$Oں{f�0K��`#R��MaN��:�;�Z���7�W1T_�]	o�^�*��c�ߢכJ
�n5��K��^a��EZ �P��=y+�%s��,$��ɘ���y	9%�G�D�n�"@��)YK_��G9���~��~N�5 �����^�@�=EX��D��N�*.��	�96�7��B�������Ps�n�g"�Q���T���2�
��ʏO����B�|� �n�T�>�^�(%%�*�l��L��o�l���
e�d�]I�kTd��|�>iL�r�j��u|W�}��J	�+�*9-:�!�9��'�:�)�If���WZ|
���x�3�+�B-�m"~�ȀRw�xXZ�
�]@��#�4�]������6H�^=�Z�鲥���R<��?�[B�)]D�Ho,x���\��ԝ���.F��S���������*���y�sp/�:�M�@����r��:ùC�`�V�P%�`N�^tR���b*���ȥ&�\:KR��ڇ.�^Xk?w�A�GL��ۚOxJ�� �ѫ[�Ps�w�;f�0ud�d գ�@�)J�P�.Jl�G5'����B߰��0VCo���^���ޙ����N`���H�x��';�z�X��>��ur�$c}��jrD�^c>\�Lc��kD��i[���(��v'-	)(S�n�	���C�?��Llz��ݼ���Z_���y�pL۾!�������7�b	G��������.��v򋸔`��j�gꋜ�	T8�/�|!Y���$p±@ǜ�y#eH�Z5�w������_�_,G���?���N-��A�b�����Í�����CO�D��#�Ϸ�#L�)^X8��y��Ϫ��@K�ܟH�����c����w�g��xKk�N�ȱdg�Z���c��f�)Ck��H�(XMN�B+�Z�Q�13��=w���G�O`��]�QWj04���PSx���v�,g�
%��Xn�	�R�a���̄nIՂU��;@* �Eڅ����!�3)%�=�d0�w,}� ���7��D6��V�G[Ol��L�©/D[�d(����ѵ��,8�Z��M�kW�+��0͇`(ћaV_����� �'����06��G��R�>�_�N�>g�c��n�yU3c�ԗܧ@q0����{���C��tKD<����m��Y��ܟգ���T����!;�2�@z� �m��N���D�9�U>�F��d����[��{���zO���������F�p�@:�<2{�q�Doq�+,����7�t!&t��A5�����3��؂�oY9�GW�,�F(��f��������L�!�	��q��a��?6ʄJ�4FN�9W�k����x�!XLyE=�]�	�t���s@>7Qx�B���p~#�耎U�\�_"L�yﺟ��f7[{M�8�̑zIK_�5�G'�)������p�8C�o����H84�����)�ؙ�����x
8 X�E�K��H�}�h� �ׇ�]��9�6o�>n!��]	�ٝ|��E��^������XE?5��h'����|"�lZ*�vV�$�&yG-;(3���p.n�зXS=���v����|ri�7�@#Da�2`��}=����u����ғp�����d�U$1�u�k*ꔖ"�����X��Ti�6N�1�|�$�$6��#�Y�3$�Q�s��~����O�����ۆ��P��cW2�y��{R$�����ZQn���H(���%��}2,�{�^��zXI�f���w҉�s1W�eĘw�_w�h�y��?%����F�2����~�6���b}.S��U� Ԣ�~O D)�ַ�r�i��=���XQ����JG(�QK_�2�pʓJ j��G'M������_�Lv�vMBO�F<����J��9Zڢ!�C+�N#�"�c���k=mI�r\�)�v��M`���
�F�%2Z�5�Y�\!R�u9A�$i�=����v1���ڿ"B�/^�t���y�n��}��ĐZh���P��j�|rK��]"[����C�8i㊮3!^0�G����	�}�u@�����R�;�e��['��Wjmkk��_���O�/eZ�b���?�C��C�3)D���sh��{b~9��0�*r�tt9+(4�|�?Ǟ{H�ݶm�~SC��.(_ɦ�qPF�z�%�>҃������KN$y%��EI���Lߣ��̪�,��t�u'��������R���9��w���Z�Ǫ�� �o!��2)�X䉀���������8�������Y�N# ��cՃ�����^=f�B9tO�>����mӤ� �Gj�ή>����؏�\�v�"����V�
Qi�¯_0� ���,������7���lMK���ˠ�m��͈U ��D���Xjngl�۷�[�s��z¡R��L��4
*�������*\�~�CnG��{_��vmⴌ�ས���K����u��V� ���4|�l�0U�`��ꎷ��7k���S��#q�����Ǻ5+�,b��?Y���6����k''ӏ�Ak���x���;le��|~�[���<-ʽϋgc���g���6�wŋHq��F,d����������	�醦ܣ��Y�#Cݒ�[��VhT5F�卟W⡌�+'�̲���b�:��`֥������7õa����ße%��X"=D�	��>��;��yf����Í�t ��]��&G��n��}g��:@7�旙����S�O�dYw�C9����Y@��rS{-�7s/$���lQ^!V������ِO$Q�uw��b�q�|h 1B�5�u:��x1ȫfP�p�oR�6�*���xn��:	�s�4�7DjH̺Xy���z�"�S�6T�I���V23�t�l�V�#ѕ�� a<�#ș�QOa���H�=h�?��ER0�=��Q;j�QF*�Y��P��$��$����;�-��Vގn_��}i5��D? �U�W�x��n7�������罊�����)��A�$Aɋۅ��-X��v�ld(���siS�xz�w:|�0"w�/Vp��A�����A��EO�����$�@b�,�"�� �%k/i4�ErF(]֠-�\4���)f�Q��8L�I",2��z�����3 !�@�;0�]�����}\-�A�!�gXMAl���@�k����Y�>z�b���"q9L�͚7r[��l���HF{�B@_�)~�މ]έ��jl=N��v��z�<��8J �P&�)��dñjP#:�g��w<9��E�/�Y��X*\9C�A�:�Ί�Y3p�Z�՛�0���{+o2n�[�cy!� ��(��R�k�d�� ���_y k,�'{Ow�������+Y6��N�i��I�#��Q��F/$���^!.ok�%$.}'!�3�Ě�o��CN���&�w_.r�tjp����O'�e����z��^K�M�x�@��}"F:�u��BZ.WU�[�8敯�n�*H�Bo=	K6��Ĺ�p�u,��e�=z&C�j�n�GE޷c"x �`�g���2��������/C��?�U�^i+���ZR�i���4�`���P��5�p��4�N߳2�XO�W��~����b\����H��~�u�ň9�<�,�1��.وj�	��粒������JY�d3���D�dF(��z�"[7���#�d`����ڶGV@v;w����bp�W�:r6�j�4#C:��F�F�n�~��9&�s���`��	
!�-KUjqA4�~��3�����&s�.�^!J���� �V�LTH��4yP��i^�`��a��V�����R�bC�*aL�]%�����c��م��V)ɒmƔ�F�g�=Z#�X9*tSW�]�Qj��=|�t�=ų+6�(`.}��7�Oƻ#�s�8#6;�%�lmf��ȭ$� �>����/Fv�p�u\-0� �(8l�<���0O��8���].2�a�sQ�S`��J������{��_��
>���,��Z�??�0M}�P��
�HX�Qf��w:~~'�����I��\DZ��~�E
<�u���6m>�8KG�2�ʸ\ˠK��2���j=�U���g��m��7P0����O+�=������X����~�'��'���~֪ޛ�+|c0�-�7��rӛ]E���)$����;��7:�-&b�8��G�������R3c�@i#C�u=��m�i����0Y��t��?|�lH�ǕVW�7H���>	~4��Wi�؝M�u�&���ƻ`�ꕆ�ؾ�DF�dp����X"7��ϑ���O�g�ᔭ҂V��$��'�^PA��!k���d����F��>w�D��!���'1mD�Lm�V`^�6��c��,	�+[)�!���ت�5�=A �Y�&'���)0�{�߉��t�Q�Q@�����# K��Ѭ�t��#ɷ��O�cQ�|䡾�aJ�u���$DKh�� �o�=#�cg&��m�4��0�~{D�{���'��b.�ON��lb�!��78���~�,VH��Y���~�h� ��9���
f��~yuڸ�Y��{DN����a��_�޺��\+�N]dg8�Iۂ�]rq�#�����n���]Pіu7��<��Sy�n�碑�nP��i��U��^�}�LY�Lvm^#���ѣ%?�d1.�ˁ�T��g�I��p���|�6�#�3��K~K�tlæ���B�;��])'T%���ǡ6�Sb�[B����oX1T��1�������a;�M��!�1$�*�Q�R�MD���QX�Oڍ..YԀ�\+�.��R,�
�[���me����u{z`�$���e��t���}���j�Kr�s 
�EИ�o�*�������N���_nC�����wZ>�7k�h�<���D����OPs�x�7k&c�j��t��N����jL�H���n${6����|=cYcS>���M�3����G�C�_���OqV��0�������G������r����.��p(z��)�=���*��K�_~�(}�TX5�����:����m3�#��>
��l��O�� W�mM��+�B^��%���a�ͤ
Z8,|x��ɹy���[���숃�L���UhT���a�m����.)����}~�Y��&�c��`��ў���I�b��~ʪG*�����zk���X�;I�]��(��,>=~T���/uFI{�����~�1�E:��Jߘ�5���
�*ާ�$�n�؈�/���jC�2�p~>�
�M���c~ׄJh�9�� ?r�h�B�<���M�̫�Zj�~�	K;:�;c�oi{]�{L��9h%��m��$ �����3���ϩ�^Gկ�,u�m�j�*X��)I�7�J�"�cdB��GͶAo������W��"8l�>9���������cwo�5�C�����;KM���D������b��<.8���'��N��+�<Ee�
6�Lem<sA�S��t�|�ːo�)��V�C����2�]����%�7i-�I�w��(]�Q�u������Z��n��<�o���T�útL��y��,p�ʤ|߮f8H	Kjf�^��?��_O�[��c��1�z���&Hi�~�9~z, j�o!F�Qc]�W�69:j9�����䵄N�8��9k�z}���e��G��r��ףF�YE���Ѐ�tʀ��M�,Z���ח��/wM�e!R��?st�w֋Cy��C?ҕ�C��dR�"�l������Y���텔�G�Eɻ�b��N?>��FZ2�N�ST���htJ��9N�5���s�eMXb�{bؚ,xQa$v�h�O�[��: &zD8����{�������W@���me��� �v;��p���e��65q}*��5o~-)�3Lt�b�y����������u�>�-�0۳p��� �Ô]�2M����3ڋsƠ��{9ȉ#e\�����/����A�l����(�g��s ��:Ly��GУ'��eA��73Kc�Q�^D%�\ALc�_]��Ղ�l������r��	_�%��N�	bj2�x������lDm,�u��C�����j1*�d�"����.���'o�=]��×؞r�l1|�|j��%ƨ��R���X������?��a�Le�V,���2����y/�ˮ�ZK+���|�
���(@'+��j���ʞ@I�ozk�?��V� ���)���;�`�X�J,1�,����N^�b��w�c��]�Tk��d]5�(�^�n��WV}�N�r�Vr{E�P�<y�'�T��W�������y]��e5��BZ8���d:��������:$��?:���kJ�K1�_�(w[}Y�}��-#+׿�g
-3T�vģ�7��+���c2$�oS������BX���H��Hw�1�Y��>�^�%f����ۉ��9����4���2e�s�'�ްU3�
�y(G��s������b�^���YdP-/�3����N�ÁZb����~F�Rʹ�:���%�C�|W>I�a��0��o�ԕ�j�L�rN�6'�C��ԏ9���
�����k�L|�����X"nR��)'}�Z��f�Wj�ո�41y�~��1�U������B�����?��*���ʍ���<�7�ڻ⟣�G��?Rי3����U�.�$��!��R��S�
o�^m��z,�Qz��fn���&���SC�F1�GX�E_R�Y:������jU|�.%NK]�j�I:��2}Kx�0�k�3�~*~�_�x5��F�Q�H%�����;]k$�g1�������;@�͔QV�h!��Y�"8'�j�:��4�D�\`�C'����a��+G�u��ɾ�Mԝa�q};��v�`�����1�9U�qsl�	@��3d@c���ʇ����W��)�f,�i��?x��&����'���|#��9��eC���H���������m�d���7wբ�c�^-+��.
��Vr-�G��4E�x�n7ء40'�#�CL�n��_�������:Q��q�}�$��}e3�[n��^�,V2���̦o}3�&�~Zꨵ�@_�~R����Rz�Y�N��G�)0^�� O��+ل�A��Q�h&9{��14�7�k�(�n���+j�6�V���_��ٓ�MT�]��/�<�s��
���	u�y	�Q���
Z�6���w~ad�n��I���]#BD9�bM��L)`+��MVq&���y�=�L�����´no�9�yzaN�`�0 ���
?N�W���E�t��Փ}���J�Ő�ykd��N[��ep�9�M;h`���_6��9x��|��������8df�U�.��	�+"��Z�v>yH?��z�п��������#cv�[�O�pDH���s]�m1�k��Oi�/H�D	5�UQ���+�U�N瀐������u�d6 �3��ϣa�+ĕ�+���bK3�f�ת~��X���j=����^N�'�����}1�I�R���c��J_��\��&�:g%�k��\q��Æv�q�.e��6��(_-��C��c$*���Q:��w� N��S6?
���V��ߡ����`Rh�1�z�`��'s}�e�,��r����s�r"s;,��P6�f2�^?��d9H����5�AŲ�^�͡�4ӕ��T��]8NQ�ٱ3^�&���ԩ�"&�C-v[�KZ��j7���>�g[�%�)��3Р�,a�ޘ٢�n �m�2�vg	�B��qp����'�[��7z�<z�q�S x�	�$�Ͻ��s�~�������������|�{Η�vR*����������8oz�WE��/7h�?91TA��C�P��/��WQn1�^��3�~� |��n&r���WbtY<��,�K�p�����l��1@&f IT���tX�Gx��;λF�\�ܨNǡZy��
�"K�L.(�5�;F24�2�O3�p!8�}Ⱥ���n#�=:<�~j|IMyd���^� ;ojK�c4�
����Ǵ�q�N@�L����c}3���m]�������s&aZ�}3���i����7�XjJ,��L�	��=���Z�{���ώ�P�va��I"��eV�%���2�vf��uA_�A]�Y�rԎ���MLREYv�[N���M�S�Q��w�_���T��������xN�5��x%���@�3�~n@���C��<��<�;�=tآ�צ��_N���=ml)��"�t���ű�j�J��2	[�R��`�yH<�s�u.�����ZQ�10<�8�(�ľZ���nPT���B�Cu-�����#F�^~��%���� 92ۢ�� �����]j��;���7G�7��z����ו^b)h�\�A:�!����N�O-xt���::��~���L
��/�~������BVs�1ڢ)j��zFe@v"��[&[�����A v&�
�D�>T��R�.��EB�#Gs��藞�%�k�������o�o�����q*��,�G	��Q��V5��FO��@��cJ��6��z��}��1E-�/"緙��.j�Ɇ``c1{��|��=tH���ˣ<��q
�,z*W���$�"$��gQe'#+O��-	���w���1�2Ȍ�|�:�;t�]gU2����"tIV`3���M��L��"�g噏����*p���.o� r�mMSȴ�H�Z��4���x����6f�ő#R�P�۰�)Fq����!d�>0��VNY�i�)K�z���ff�ֺg���`Ӈvi�4$�Ϗ� Z����ZK��Q>_w���G��8�ef�I���[Z�Z���#�%u�Xb���Z�O���ms���>(I6X��2��$F)oL��sK࿽,�CE�ꟶ�%����Ê���ܽ�&s)�^���P*�`��0��I�T���;�Ƚ꽐˦��uy��[(�������e�Yd�Fp+�0t��|�����)V�����{�L"��F�X�c��6}l� �*�P#Y'�՟	��-�o&��w6�8�Z�6 M���/}����;+@�k�/"�Û+m�����!</�﷥p!N.^K�t9fsFJ�8�G��[�MU�큔������u���#Ur÷����S�B����IdeO�s�@憹��>�5��	�ɻ��(�ܬ۷��K�=����ZIh$���V'Q�]t��7�c��L��F�eC�b�O��|��'E=c�<!�X��EDu��mA��s܉�'m�Y��M�8��;��8w�жeNcoi�2����\F��H���>Q�y�B{?[�=5���&��s�v1�tK�m ��WR�P���ڹ�Y�,>�?(�4��y!��5Qټ,?���&�1���A��(`��������!��/������ ��$_:�7٥�Z�{�LӀ/�p�m����`:������=Cפ�GO���Dfy�gJf��"���x<�u!��i*dm� ��*�{5%�ޅ��	X�z�b�	�3O莣4O
��1�s�@sD��lSh��f0�	n�`�?଺���h���RO��5�"d�<\�}����m��gN2�M'S��.U�h% d���-ǵCnUQQ=��M�5NMx�毈�X�5�Y�+S��y�a@{X�D�.��"S��7���MK:�jZ��U	P�z :�V����r`fоM�k�3��}`9���pf���|'	��	:�$��h��EF�=�4;����&�YG�*�<kBXi�k���b�\�����ۤ/�V�hfk�R�o;�⇈�TXv��O;N�5�mcRg@鍑;<ۿ���+��;�!����qO��΋v�_����>�@ծE��MoL�@��Ɍ�[*����9o:�O�O���B��t�`�h��Fߏ�H� ~��-�v��[�b�"��ӆ`���'I��Fw���3�`9�Mh�m�9��1lM)���W� ��*������U���q�^�[QYfw'�J3���Bќs+$���CĒAVLA��U�Cp���Y/�FJw?R�/ �p�O�"[�����>�`5�[6��|�`ϕ����	 �s�PP~�b���gLwX��G�bW1Xf4rԈ�0��c��8cu8�RJ(V��qh7����!X�Z�ӟ��.|<dI���Ǘ�eIk��ΔC�$+L��`ѻ�n��Z"�E�q�Z)��O-�x��Ih�Ƨ��zqc��������~T�=: 	�z@�f�%XD���h��m�������x+��5b� �S���shN��P])��k�hyψ}�l�~h��ap���f�s��!21�����>~�y�C9'wi�T�'8�1��Ռ���4�0��v�-"uE7�|pܨ����~�������7z\�j��N�v[ť���Z�����.S�婝A}���;�r�e'�;��U����m�S,Y�����Vvz��2�F���^�lf">� '~�6@��N��X�>�)�4|�`p|�ۮ�K��ƼP�}���Q�s ;}�A�SV��12'2�{�5���w�����t/ӳs;�5(V��bq6<�Ù�υo`^6~z%�]���ijK�� &;��\18��/(���T����9�t�*-\4{�T�}�V��aT�@r�צM�h�����o�5��$|����5Ռ0Q��R����(�R�c��v��B\�rf9#�Z�q��zt��*הZ�ǚ�2u.hAz4���sp4t�'΃�����K$߉ȃ\$(�)���|����iXT@�+<���62��_%w��	a$~�¥�#�)LSGg�
�p;��-���Y�0`5�O�Z&[Gq���ᑿ�O�4$ձpR��`)tZ$��ZN�TE<�)r���m��(��b����*�0V?ʨ���i7ZH�<s!R+��[f�G$�p��g�����1��q�����>VE[�X��!��6 �ߝ���|���+�S �y��1j����ekY�._���2#�(�$��.{ ��+�.tgꝐ�'.�o�EE6�mLR�A�i9րa��$!i�$v���{�y�W}�.7%�i�߽���������]�t5��8�m��Vˠp����oD�	��^�_��y����%�'h+�zށ�`gMh
05���H�pR�:e�k�L���~8�уM!�DC.m��R�8f��4Nޥ��9
	���sq�e�K1��X8���(��3ݪ�~������'�k�'�X�j���q�e�0�>3	dOJ:F?XK<.�I\߳���t`� qQ��V�4;=��[$��c+4���p��>G~����lŐmТ܁����'?l}V��@�<B�W6S���;�[�4g��#$��*9v!����r
�!�(�¬��U�@� ��.h���d�D�!�n��B�L�p�X�D|�/�l�kT���|􀮴RzT^ȝ����Y�x�K5����yA�}SF��ϻ��1D�`�> eK�Ky��Hڟ8��^Ģ�4k9;�[��ΕKu^|w7!�͘��^�sШ����J�{�ڧ�Z��@���0\����&b32LDV�����J�K
��7���y�@0��~���.2t�j7$�~Tnҗ"f."0��	��k��n�!�H3�%P�Í�d��Kj>��C�(�e�c�E3ԯǸ�;f��<%ƈ_��N�!�D{�XZ���bs�W޴��V:9��u1[0�!?(�ooh��f����.>cX�&�x"�,��}#�+XBkH��zs*H#�0�b���=�@l�+6�4y_�vN�W��'��#^�,i���CϪη�*);�~r�7%�ƣ�۠���Dq.[��P���a�%���N��׏�K�N����ZJZ����W��X%��_�b$N9s��>�]	�bV�A��*Q5������,�]+�6��u��\�Lր<���PF�\��%\5F�=�KO��=9��\�υѹ>�Un��Pw�Oab�<EeR�i������ Ȭ�Y;d>`����u��=�A���d�Y���KR���2�P�Lq0��,ڬ%d��lQ�p5NZ8RE�"��ҽi����/�8����{V�r��1�ӽ��7X�l�+�5��5/7�&���M�B�R1)�g&�$�8�L���~u,l-zS!�Kg���1ѕϭг���?�oDD�������H��R����jNKt�B 3u�h_�y);ҭʱ���٠�pa���u����g�rbȰ�P�߾乙�ηx|�A� ގj��iϱ:����byy���?��*�;�nOl?�c̱&����Sk'����P2��Y�9�h�s����$P���R�k��ym0 "0�~l�t9�m�����ƣ~u�4W�ҘU�ư�o�et����D���`1����<����9���B�b^5(L�R���19�\	T���)f@�7�!C:n��M|HL3��J	��N��D���!	�wk�"�+e�Q�@��e�~���yFo%�G;!n1n=K����=���"&���ȓ_�%��8,(�jJĸ@$�َt�����j̓S�]�«D�i]~�g1ฦs�L����~�s:>!E�	*���:��@�R��;�~����/�8�#A� 	�$y�:�V*���g���������]�i�-<-����d���-�]wzj]Z�[��Ȱm��0��(�<H��z�+��E�e�Q� 7��u��c ݒ��z����vi�H�� jq^W�Ӻn���n�Xs? C��K0}��T@�:��uwGf���U��ũ��;z�^a�>v�&#��P`)U��
5����8�}�l���Yу�_�s�;\�G�|�Ң%nR"%�TOq��QYWPnKZ������>"��n�@��&��g�;��ź��S�M�����79���4p}qB��	C�'�b���?�źlo��Y����΍P?`Ma����Z &�����k��8'Hh�|5��&ǡ�A��s�ό����"��}FX��,�:i܋d�\�\874 ��&٬� d�W�+��*{rޭw���*e:��ʄL�"�4QJA��m�uX[0��ؒ^�3�
&�i����s��,_|y������SVb�������̘*�K,C�A��;�d�6Ӟ ���n0�tq,���֑�'�f����v+ݎto���oF����8/�<rCi`R�ֶHH_����<���@��\���#�w�tkjp�o�F<T�~��.:v[�����sy%T�J0�),��ءփFUf��V����f*��jѠ:@|B������L�^�v�ٴc)o�'OY7�@�)P�ô	 �`6!���r��׎'v^?�|>񠓂��z��'�wԟ���ʣqJG�O%�K{g4 ?5���8rۭ���(�sA�W-�@'�µz��H��\��,kN���ݺ.��KشQQ�5�%�c�\c?Y�44��1��@d_ڂ�x�{�+�d�Ԯ%��Bl۠����+*7����޶��m�iK�$��\R��{�rbE�ZS�#�M�m�b]�>����e�<�9'(@zb�y"=�HH?u��pL�-��R��"��ߦ�o���lGm��jx`�|W�T��zNt�Y�	�V�xh��hXOi���b�Ȏ�^I�:�K}�k�w��t���.V�KB�dx�Y�9�!�&渊���l��o�p	C�g�dqiG�BOR��	�D�Ϊ}��jq�&5Py&��Cz��z��l'&,I[5�������pF� ��!v��#Q1����t�u�_���h9��v�'�l�v��ݐN+���1��b�[���K7lr��t�������Z�K�H(ғ2��/�/�4�y�F�B�� ��D�Px5Qf�����.����J��iU��}br v�G�K
󙨫*�fu�������w�M�@��ʿB���W��9l�T�s�%�(
; ��ȍP�>GS3�=hV�|/��+���֮��$A(!XS����uEN�*U�=I�������qq"����˦i���M}&����ꙮ���B\����v��Sف�]��S���'L��V��CA��M�xh3?Wm&�mc|xY�(G�;Z�'��q��	1���gGm�yI?;&�%�vd�����q�W�;��V�U�\�A
�\�?��$��H�Q�.�^.Ω�%1iI�1��I�PRS51��i@�8�ʍ�0�9`L���������=�-s�>2�Gڟe.<�[+ד�eI}]PwNĢ��Mx[)#����է�׽S.����-�� 3����k��Ҹ�"̔� �y�I�y�e=��.0���(�ئPy�F?3����6{������r���Un�p+�V��w�q���W���8�"m�>�u�/k?���"��(�?2�;ÊUPԎ
V:���h�ӎ^]�̧v��W�W<�gܛ�C��Q�73�K1����[�4�{T�)���<�kB�Q��/U����eڿ_��:�iYܷ��ŵ�0K�BD/?P)/���V~y�Ԣ��j�Yr��o�������B
x'��z_�d9�5q����js��'�w:]	d^b@�`���:mIڎQ��� -HÆJ���Z�1�V�T��z�PS>$��d�k��km�+�#`ޢn9�-$^J��T�}���Z97b=�p��x�*oC�&|��!]��_���]��/��f�R��/ �
�#�L���$�%'�f�ц�p���q8�bT��'#z�\�0
�Y&V����
�U��b���ҟ�����}���=�E�d�2�]ؖ�� r��j̧ވ��祿�#K�cH�i�����e���H�X,K�t��t�T�5ր��!����g/.0���_��m�d�fUB�_�1�!ZaĽFA/�
�����ƨ��_O�Q�d�T�	i${�����w@�Y���]DcI]��E_���*$//v�%�prR*`�����4tW	쩾�Ţ�P�.J�LzA�ҷ���cس�_ua���}:m�>
^��-��1�H��m��3Bƺ�>>G�˄*��H�FNVTi��zr�cf�i&�Z:�$-
5�b�zɿbie�h��J��A<�$�ns��^�nVb�"+�W%�@r��%|��P�|I�'�u1&��W\�=�2aAGZ�jo稽Z8n��c�N7#�Zh^P����\H�\��D�'�YKDh��Uw�VnYˇ*�;��(q6"v8���Y��s�$n���J����b�k'B]�u %�4���3eEI.0�AN4X�Yr��7-�v��e�nf�w*�ᑺ>�Y�28s���.�֒���Ko��=9�6�g����Kڵ�	�d����2�:�>)�=J��&i�\���l��i�<y�1帞^j�H�o���f����Zz�z��@
Ͷy��w��o�y�p�k���ٽ�)�� ����P��[�z�й��6u�k[ut�T=�:�x���]��ʡ��������?�5(���b�N�����_o�^����3�#pP�Gb������	��FZ���,��%�ݘw+7i8K�r�A��Vؽ��R'HS]��[/��ȵ��al����SV��[�\}y	��)��&���	���0�X��32�KI"�T��*�)9�T�?z	��ϦIy�z���,l�lV~`T`��26B1�I<�V�F���ݝw�������ķg.��D�"p�����-���;θ����B��y��#q����bԱ�	{'q��d�+@�V7�3�m�GS�+�,��-��d�Nُ��ĥ,ᄔ��}��3�3���?��t�5]g��r�Gm=��6��5�<~�*d�Z_�W����s@M'?�F��qVV����oP#�!��L�{k��7��-L\�|0C�P��.E���3�9y��x;M#r�)׶-k\"il����
��ThTӇ��lL�i�P�o�I�v%C���:֯���:9�eS�7�X/�@��\�8�B�y�}'>��!�DGE(2�Cֶ�E�UퟣU�ho-w��H�Lh)��0c�5[r9�P7���d���"*�qx�BrѠ�jN���8g�S\��_DL�'�]k���#�.��!Kk��!�L	��1t�߾QV\��|]����w	��͒ɏ��=�P>\����'�`�j@�4�1'Ч�Mg�w�=������R]U�$���7��&8�cYi�r��-/�B�|e��G
9x��1%k��E�u����6������4��8 cԂ�¦����i��	5��ԉ��(	=&
y^���&�/OFL����lr����pI0{J[��	�O;aWG��x���@��V��k�]d���h�u��)\��m?�� "�m���a#gS�:/�Ϸ4�T$׃�{P��c%qU�H��g_��|d-���ZLh�qg�J������O�Z�@*��K�;����/�?��6�){Lz�����>f�� i��S�YRހ�M�^���]�xe�����I|��/@b���耯ZƱÄ�b�����B��n�γְO�"O�5y��M$@��>%_���I�n����u�+W5�k��ٴ�
Ѝ��g9�o�9�������N���k�����H���)�ߊ/D�&X
�� ن7}"����bQ4� �S�\��wI*���"��`����I���"o7��:�r���1���q��uE�F�(Ԓ��������{h#�m=HS��aTq�(K����cQU��`*e�J#�.+�)����
����a 8�hu�s�!�ylALρ�Q�c��윎M�G�VBu!w��R��r7�4G��)7b�!e�R���S�002^���-�2'/qt7d���1)���m�����@M�4��0*��T�o[�&{)&a���V������SG�HX;��0��)����Z�ܐX�EJI���`dA3q3]��^E������aR��j	��ygТ�KL��O�^�N�p�?ؖ��ן���ۋd�H��;� R��A�]�m�y�= !��s�\�y�1��3t���_���\�R�����ئ��)�2(���T�o�Ic��L��F�1����ʭ摤K�A�����Ϳ�h1�#��z�u�|���\�ǈ�|២{��=픨75:���EQu&梤��kȋ���Pi��#��vt�х��B<|#�=�~r�q3q����͉�����ݧ���B�t���e������r �J���@�ϵ
%x�ϲK��� (���[�ӻ��'�G���;�(Gf/�؇��1��?�����R���)�(l��T��� ��|���y���"�Q���4����;�BF7qzi�w����Zq
��`�\�/����
�z�8���\�;9�ٕ��ڬe���jn-�OT�Y�!��K�����x�,9��G�v�C�G�&��fM�uOy�μ���q]�bjS%���<|�
��/-��*���8`c�{�7�>�<;>�T>�/bz��Q�i���i!|���)���pgh;
8)��<�¿	B`�U�,ݯ�^k�0�(�)�i<�)����˩��/R�"��� ���7��p���p�5(Ƕ��;�}c,��_��h%�&���0��T��<DŢ�;�e12�*�I��4��`=@&���]��*нȮ,�Յ����j!��}"���.��6��	X.l���Jq"�(��}S�yI,�P�1*!�M
���#�ͺl	�4��;4'k+�TL6���7�*ƃc�@u9�� `p�P�Ă���hҼ$�fC4qyrDs�d,��n`����~�q�D?;����0��<`�<�h�L�%غ��h���Y���<�T �w�̓*g��鉦��ȯ��|9��R�O��Ғ��57毵��S��ZJ>(������l��簉���2�vP>�K���ZH6�܁?�Z�{�Dg�˒o��uF�A����#q2�I�p��T��Gg�-��о���Z�m���W�$�2Y��Dk(��;\���]6�?�uU̐S�/�܍d=��۵���y'v�����];$����{zW���lT��u�W�/�e�Fm�{<#<�TΟ�;�	d��������|��˟���q��>��}C��N����u��3��; :��Wc|=yX8 0��ֺL��7ld0^p�����ڙ���ey8�"p.x�{A#��L%�����F	 �7�@*�nkUm��E)�)�~��x�ë�ǐ�����d x�w�q�sc&"υ}��qؘ��)��/�ā���j�7�٤�-!G Hr�S�ug.�e���T���{l�*7<p����_	sm	��=�|EBv"�&v����w��0l^=�tXL���Y9L�8���e�4�4~~#�H��yƬ�T36�s_�^��)�M���[z1�� ̩4�>Tp��
���]5`յ�8D���'}�H��"DM�d�#�_�)�PXX���"��l� �Eɀ�7(����8w����/b��=�*��p�c�Z�*̌l��߾�b��]� (]U��_OC* U=1�</�aOw�s�ˀҾd�M��hn��2�d9�1��V��C����v���p���R#����1�f��P�W���n+U�H��y�X����7�1��F:F���@Av����q)�=fu;af���PI�R����J�Z�@�q��"�=s]W��T#��9�"��E�1��[hs��' V��`��d�ixh2�3r@!����ʡU^9��"A��F-�e�,ڠ~{�x@~��	�
^�u�A������W�~p���&��t��DU�9��A"dg��� �c��AU6��*32̰�(�xRi�O�Jr}?����Ʋ�C�n�eF�ίgLIRP�~��:Gxh�dÉk�b�e��\��M�u�%2T��u��ę�������c�������BC�(�xU��+��|�M���U�?�)�d��Z,����x�h�zW�6y�N��D�I�V�
�����\�o)5�z���śL�����w9�Y��y��C!m�_�#M�s$ۯ�8ӌ�b��c��-a̙�p��n���������nc/�t�*��1�u��-3����Z��{
�K���vۊwa+̄�ե0F3MvHD�$�퇩
suS�[��m���j.������`0���G�<�o	S��T�8�^f2"��J�5nFޫi�+!��E�D��Ȯk�CV(���B��,1"�n8�]܄��N�HkO�&~e'Й\5K�A��Dɜ�n^��cJW���J@�bo[�Σq����i(W�IH8
@<K����;/�5̦�;9f���Ʋ���]��6)H@�{�S�{�#[JPٌϔ,{[�u���jÚ9M(�j�9V��:����:���@��l�=���42�>2D��I^40�eJ\S�<l�h�<��.���_��P���V����/vj��/������[���F.N�j/�QA�XT����Gy�!�l����i�	�Z����3z�D��;W͐n~���@�3s��(5PHg�xz��YA�طm ��L�ͱd2�,#�m�	[,�8p�3�"�����2쎹`�΃��a�A�%I��0���b�n�:�	f�SUw�5	�`�غ�Gm�1�g�f�8�[BU���WW6�FW�",A��6����Z.ū�%Q4��#���D�����હ��������r���� -���ț�Ix!c�S]L�d��c�[�܇�i��h�2���BcC ::7"�H�|jW���nw�%�z�,��G�@�Iʸ�H<'q��� $�����j 	�I�� eb`��@+�j��Z����Q/�Υ+'�eS(Dh�Qt�9�xM��뒫dF� �����ɔ��hKA��|$�B/xhn�Ԏ��ǁj�s����j�m2���ä���\�n*���|�E�َv�pn�x����F�0F�1���kq�n�STm���kLC�[e<e`2ht�f�UH�LL�t��� M;-�_���	�P��0ӛ�<�N��4��,\W�����jBe8y6��8��ڣ
#���ǌ�a�W�$��ݲ_�q�	$V������o��H���9�>�oY��_��B\:k���K8��x�=�ן��(8f�Bo�3b�k��֦4���\B��2���5��w��rt�[�ݕ����o�r���D*W�f��l�����k�7�E������&4����P:a� ?����h(���sC�뚮VM�����	ۅip"},e�)�����TE�(���
��7˖�_7������K5h�#���^�9=��CIPӐ�r�S���[���	GSuK�8�i�/N�*��0 �~V�Mi;�纫qd��{UIoʊ������c�����+�9���}2>��6C����uA����r���-�WX��q�Ȝ�u)��}���?]�����e5/�@��-V�������	�+k���:7P$��ş�tV6l��Vqj�}��z�e�S}�����n~��N��-�vP��xk��������w�� ��q⢟�Ni\SO�g���8<�)xq$A��p���eO��
lT�C���W�l�I�3��T���eY�$^me�B�|�W�&}�kw~���e�}��	�M7ȧ��?�*�� �c��$R�y��[rg�%o�� ���t(�vq�Ux�LJ>#�Q �cQü�Q�K��(�~��m��٭�[f,֯�3	��*�`$�pEF����]+����Ҫ���ȶ��Z��JR�F
��W���J�G�4C�^���S�x>�V������2jװ�d�I�=P�W���]�Ex�o?��X:�<�H�Yn52K��Gp�E!����
�~
��Z*��1�101V;�U�, �R���Dv 	AM�!�NO���q���z��i� (��Sf�Q��#@}"ܪ�S�Y�Φ�a[���j]��b\�z���6�;��ư�tg~k-�ޖ���?�t�rGq �3����W�s,D?D�	Wv�
�������hŅ�5�N��c����\,��)A�xA,�d�<p^X�E �������GY��L��	��Z��	��w�[�'���w��3SY��ۛ���������e���w�0O0]����r�Y,���X^PfSڝ�)`ZW�/3�1��ÙO	���͔ҍw�j�7�;��}faY����;&�(F��4%�툵V���Pik����?%6:��A�MNh�s��2<�*������V�/Έk�W*���K9��\3�Y���lR'4���^�QC6�v3�I���l���]r���H�]m��#��S�>wr�Lo�K|T�C�8vq:%�������l'|0s��z��	��Vu �r�%�or�?����;�{�_'ɻ!M�OX�ke(U��C��A<͉/f����$5�"�����:��a�㛡+��(��+zV-��^ �MY����u�Q@Qj9;�׬��VV`?�b�0�����O�R���\��]L��VE�qg@ݐ(e��O��.��=Đ�'�� �]PJi�<1�@(�uߟ�Y�^�<d�jxvrZ�D�@N�5�抸h��o�����3"�/�Cĸb�ك`ė��n�4()��5߽!=��AzOy[�������R�7�u�=�7?9�-l����1�_���4����-��4i�~�~�i}0�� %D�,�kYN��8�Zo��c��|
�Ŝ��9��D��V���"������yC6[B�ۺ�� �������6�FB5���"��c`�5����˅�#ht����x��^_��a��zj�����J����Fq�V�l"}��҃�~cWFF��,?�����x�ѳj>� $5�F�ű&Cz�[����ސh �č��W�� N������j��uN0V�՘�㟬�/%�ٞ �~��^>��)s[�S�T����Q�09�tiv*E�3�j�,O�|����#��ǼY����@H����ֺ�1Y�/�J�b�
��
쥽���I�qX*��[�D*�js2�?��ՙEc$��V�%�n��	�#��x1�d�ϛ��/vV�J�ژ7�����78b.��6�,��Ԑ���꣗��*�Q��7���b@Â��`�>�*Afñ��Ƀ��h@M���m�Q.�LS����Ԗ�lՆ��/%uT{�����<�Qh\^� J�mu��^k����۷�����#�������E9L�Ua}�/P����u���8v}�� �f��]�y�� ��Z�_GVo�`	�IO3P}?���.{2�>8�F�Mq�S��ƂgKU�,0�pYA��kx�:�{Ec���U��Rxh�+'��H%$d_��cк*���;���B)HܑR���)���}7-�5l�o��`{v�����a��������X��ߪ��u�o�����H��h}=k6�9z#��W����N�P�d�55���Oju�21��Mڕ�,I>��F9GXp������|�+ =ؙ�����]ʥ��5�^���8���b�C��P�ƪ\n��\|9���aS'�d�P$@�_�tdȎ���6Єa�N�P��ѡ�*,��ɛm�c�m6�x���0������ʱ7Ke]3�4$p���R�D �|[_ʘ�N���X�r���z�y��ь_=~�|��{г�ݡ�x�!�e=�S|�%&,�9��]�n���w�.�$���	Oz��?�ѐ�`����t����x�����I)��s�֨�����^%�DAO�,Bl>�9nx�[�oqե�ӗ�Hq�U�]H{;��p[��l�!0@���cf�5�\o��k6����W�%��j�B	|x�3�U$���<�p{q�o�����>���٫|��r�R����m��b�)�m7a�w�Z��$���q3�	�ѵö
����@�}�%R'��&q	����J���&i���`/�D���|3L��Y�<��T��f�b�ʲ�{�g:���5�bǚ>Kb)��fgj6F��?IpY��aJ��������Rb�rH��Q_�SZ��u_�=�z:%�b7_\�x�Au�մyp��w��[�Wl��z�tO.E���D�^on���ɔ��Ō���f��p���_J+VU/8�x��!�r���Z�%�����$q��%��$0�ݍ�č�~��@�H��S�~�>E6������c1F�~�'�{�r�h�{>I��ǡ��r��kRP qY��
��p���e/>���g�ߨWcR����qzP���Z��?���@�y��4��5�����_�^������c:���d�)���ih2��)Xf7�M����ㇾ����_���V�9�A1�����dgOc�n�A���y���M�J�@�o\t�
�Q�l8#���3F�ۂON�8d�5g�@��
�X�:y��>^�}��'��Y�pVK?���\0��`�o�nh��Z�|5�V��O`<��2;�1*]D!�#�b6vJ�q4C���߇5���k�6�bm��	eNG�C��.��55�k�zubǒ�DH�Ϋ��>jR8��Q*��b�zJl6�׵m�H,7����qj���+��A��[r"�ժkK��ƀ`
O��2X�{i����3O��C���������i���{��#�_n�Ip�yh��o�P}P�4'�КUU�E���k���I�M����7w%ud:�9p;D��X�=Ѭr�$P3�&��s�J��SQe�cx�V��O�>�����/m��+���R��Ն��29L�p��"b�A�]���
�`Ib�R��{6�N�Q�_�	\��N�)���V�[h���]\*V�ܺ&F�;��k�o]��	+�Єf�i�Q���2���LP�{�0u�=�.�A|�a$�)`I��H�:@�kX�oSLQ��u��n��q���?7��t�D3i	?�r�T�E��DlII�\a��	?׃�8�)g�{�?Rrl&��7V��ޔ���7��ˁ�6�݇�4���G�ڑ�K=�K�{�d���_��O��`���l�N~%�LC���e��}����Dy���n�؇ Z��g�6]�
���
K��Y��jbTD
%�h[��~�So��׮{��q�����[���6�EB\\�A�K�,?��OW�gT���@$�����A1���8������@�FA8����i훂[�C1�/�Ic6]�����5�ӷ�+4��;>.2ǧw<	�Sl��HL�'77�*�	w:^N��u��E�q��ŷ����j��ז�	�/�Z�>C���6�6�\�S�1���z�t�Z�҄��3az��}Z��П�4[gc�G�[Dr�LD9���QZ�{7�/���������������6��h���T��
:	�D�c.UuѰP�]�j��� >�_����̀�ߧG9�O껠?B�=5$lC���(����zJֆ]=��L�3֍�a^v������e=(�:T�*�) ��a�]�P74*]V���g��p�#)�\�k2�v����}¶W����v�S�EA���A�B������ѵ92�8��m�%	Ju�����Z���*qs������j3]���WT��8�����¨�	w:Kw��D*��d�1As��������'�sj%| ��O=zӅ��q�-�=�c!�����R�^��/li�;���?�g�d&/��~���T�N�#=��X����[O��{�<(�X��$��%_M3~�)g�_9a:�Y��C".4S���˂J_l���@*Bo�O6���l��0a���<�s�JE��ʷ�8�;cF���VnxZ�p
���rq}q��-1ւ�9E-PT����Cb^����$!������L�[�J�ZS�
��+/��MC��M:d}��s��x�O�Gr�#�����4ྤ�+�3v���0ΰ�d@<��yf!�F��n����4&����EyoR2�L(a�D���:�j��cM�P�9�#��DET�t�Z���n�&��H�iWD�5�he�hN�[|��@c�]���r��,�c&�O
ط�?<�גȤ��t���as��<G�N؀!m)+�O�Nk,-�����on����:5Q^c�B
T��@I���7WI���6��0�}�\�K���en�2~��	��!'b�U՜%�'�I�*�!ӲĬ�{k���s�Z�;��B�ꇑ#���[�kW��ا��C�;��Ǚ�Mqc]j1;�^�`�)�E���I�5�{z��� z�8�%�۞���{C��$���H�f��t`@)��c�|�@�l^������@ˎCb:	�qz�R�%JQ��өp��^����e�=i�)sV[�[&�C���b��v�tB�����L߷ˊ1#����}?1�HMa(�_^`W�0J�ʛPktH��bo�'�^.q��#��n�:x�o�ܬ��j�:~M)Z��ڷ�~�>/�顂���(��\EN�=�����P��C9����.�RFN�`��ɘ�U1��;sa�C#�=��oH����7y���>e}ø����U�pO�G֦�1Q�+i=W�pZv~�=S��$go���5~����h	�e�E���v�T4}��$Y/�|��{Æ���N�J�sS�?�Y�)���պ+�6q���/%W_D�{B��� �t��+��E50ؕ @�}��zEׅ6 ����.���}[m�ƅ�/��唂_>�[�@N%����6Ͼ����I�ao��}˘F�w�ZC���\"��5�DP
��څ��J0M�o���r$�K���m�{���7�	�g�إ`ˈ��? ��SS��[��9��@L�q��rXdg�C�? ����<�K(o����mQ�5�������1�i[�?y0�x3�+�Pӟ���"��.Q�{i?`��ŵ8Z���F��ƋK���3a/)�X/s�Z�O	�3`�-�Í��i^�S�r��ʹ��u*����iQ,�-�эM�J��w��W�z�c�P��aG�:�Nn_MUЏ�R��՞-��{�Z�δdg=�G��ig?_�&7�Dp��s�0����M�oѱ�od
[sT�.�K�j�����h��7{@�*�;��^6�+?r���;�
�7�76C�_Y��Hw�KP��p���j3�"k�L�qLVCܛW�z����X
��ݹn�32��@�� Fy���iz֨��7�Ä��"��'��U÷��~����C3"�p�_�>5��Dt�6	�Z/�)����}G��z��wJ���L�:<���3��T�ZI�Z씷$�E7S�0���yX�?��� h��s�3A�[?���@��s`Їæ��qI���V|Q{����m$=�A����f�T_K�
5��U�
@�{UH4D�.;Yp"R}��<��s���prW�5S)rs�݄���q�I�'�n���-6$S�B˵av�ԙS����-;5KW���@�qS �< �ɢ#K�#C&Nd:Z5^k}�i�$N��D�{TǇ�!�1�$>y��UQͪ�-��*��s��Q�ןLMҒ��%�	���=$��=@�y���#����H8�J���Y��շ��6>��֦]2����-G�H@�x4x#%ix-����'�}�B8���~��9A��e%����W�n/7�ӗ~T4���<m�/PI>���:$�Zb��-be��e`�b/3j�A[�\{�	�k��]�J��,�6or�C��oQ؞z��Z]n�x���XC��5ٞƔ�Q��8H-+���.@c��')R+P6��>�S������oǶ_�hq��nOc���O��S6������p�Tm��Zx��Z������rx��k�]Qcz@������ϫ�R#�/d�Y}��S���#��\���Ⱦ�õx���./��5��7�L4����S\��glORV@Wr+�$�^���'��Ր��G^n@�'q�)�e���l���z�N	{��ҲE����������ƾ�Qzt�@�C���i]I�S8��؁�4B�c3���^�,d��L!ajp�I'#����M0BGj��Qs5���z,���3���Ֆ��~ ��%zv\(��5��V�
c�1�|�2YKa��;8#n��0��[o(0Z���2�/��vu��S�-���*�e�40��ۨ��Ed5B�sA`=�i�O!�4f�-_�ʒ���I,����Y��ӹ&��5��	Pe�T�F&�:�P��w3��V�c��tk���=?}����r�=9�rL�<�����bӔ�� ���@3��k�9_{�����)e✣�ߤ7�%t|Q�����<�^�Y�>�Z.G�&${�
�mǙ�Ħ%���&g��1��ݳ���aߗM{�k�T:�˵������DV���~@N�'P��,���T*�6�3�d:'f�y5��@"��ps`���ح13���j���`�+��	
?1�,k��	�%� gG<}�T�BXF��pB�m�*�;��n��R��m�c�+q��u���"^R��sr*A?p��{9����2��!�(�x؁�6>i�~_>����
 
�J����<���҂{'�GN����?���Z,��19� �),V]�V�\��]{a׶��%�"�킼\�N�2��i���#o��{p�&�;�Z�`��
���" r/A'�*������]|����Q��g�>������v~��=���:�������������3Yp=TJA��'���20	YRY�!��u {�4���V���v�K���H3�h(��(��m�%0�F�P��c*�4�{�5G^ͨ	ձ��F!���v��ȉ7w�&�J}���D|V��]�Q�(�zHA�5�B�F�M��!J�_���|M������Nh�-Ū��AH�	�O[s�A>D�'�&p:	,�)�m?���l>��W���GL�I���R�}E��#.-�_Z���T�2�%+-���l��GW3y�<	oMv_*9h�'t��,���D�ꍋ�2��t�J^��UK���n�-�)��f�V�k�3��S" �u�Z����8>N��Mz�o��Ϧ�~Z!�3Qt�,�$��"���}{�J����r=H�r��X�nA&Bx�fzX��g��[׳K�=���Qg�x�ߪqz⇲�ݘOHw���Ip��lԧ�x�!; I����v���[�]Tj�<��4�B[���M�Њ��ڜ0�y�V�̝��QN+���}��a���.=	�n��8dK�;R�&�.����i	�<��Ig�E��ms�'�"�=7�����
���:3G2�n��q'n	qo�`� -��L��a�ڞO��ّ(CөnIMYn.nw�&Dґ��Z���g)2���uo<t��	��e !U�8��:B��O�O	��s�t��ͻ4�搂W��j���b���w�h`@?�{��L��}�
�,�tC+��;��b����$�щ�?�&L�7��
L1eg��xw��S����]=�ӏ��i?�5~�ɡU�O���7eo��s�j�S�FW�-o��s�l�Q��B+�#(�PSXoz�3*���!#�I�r���=�]���d���~a�RSh���0��u|U��(���`A��Kmy�����6,>򽜋{I��j�c�W�h_G��w����bYsw�P���k�R�+5v�`h
 ��+=i�,�� ��C�f�}�BXd��*`��t�� ��/I�����x875�n���fc(ƻ��$s��,~����FW�j�ZP�lE���_ٮ�H`��6����d)t"lk��7D���q�±�i ��s���h��T{>,)��,�崢�<(|.&e�
�����v�W����ÿ��j@��όT��r�C��ކ~H�i��(�]q�p�.�@_g��W �9c͵#&o[8��B�#&�w����o�s.{��f1c����h6��Fx���ʹ+Wrm�n�f I�JP$�kz��7��)c��� ���y縒 �\�c ��e�m��S�2�;�o��]����G��4h��c�m-V�+ɻX7r zR�B$�ӣ�����:o��EnW�,�)�� <mU1Z��i�Z�m�H���:�E������wm6T	�]�yKc�ǆ�ެq����K�ޟ�@Q�L$�����k|&g#I�}_����3���oLa��!�dϢ&o�eÍ)�e�B�fN�,d��Xpo�y���)"���k����c1؝zuV�	8�Q�h��Ŀ�~��]�T�'����m+ƗdE��D<�~�T��ڔ7B�l$6rF���e�W���#��L��_O�Hv�G}Q�KV,t�D~�/�He��bR#���7D_{��m�Ƕ:AԢ��J鎻ԸZ��'�Xc8�7%v1��F��{��c/��_���pN�k���g])����8���`�N�sO�i��*��M>ѥ�:���M�)%��펬�
�/7�M�?� ǽC�n:u��J_���£Z�d$���:�D�7��EH=�ft�O,�\u.ga���)O�HotMl	��_[��E��|0�?�#�ۭ�%�'M�{�N����e����3��%�o�5&��e����6a�`V�e�4H4�+���p��B�0�]��]�_���=�:G��K��;��̟�ٟ~Ү �$bh�`j[�-V�P�t�����~��~����`�~��}OTZ2��_���)��/��8�_�mL�NF�K^����S�z��rsz�ѬZ�{���7G����E>M;���(0ш[��Z�P�Z��0�-��T�~���V�,���%�"Fb��)����jmm�����W�l�ZI�-���$p\#P���;��5��ѝs��0���I�g#�O��nx�^_�߁��7�_��Mk=�(.�ʼ�ě��Ns���$d�����?��T�����[����x;�P�B�@�ת�A7	R^b��htɢ XF���V̷z3:m��V�=�y�@�FN��V�����1�G�,(LkÃ/`����(ea�∼ t�!D��6������S[�������Q�-���m=
mN���딗1HV�m t�˂�x���������`x���P1'���=�D��.E���3��h}>
[���n�>�����+D�^�~��=�*��r��,i(��C2����9�����I�=Cw�-��vDC�л�����l�~{*���+3�_ h��)�@���P���b]}����'��-�"!�tn�C�h)�%�v��1��]v1Pq^L�ϑ�M,��!�ޙ⌣�0Q�Z����\�9��b�����շ_�h�u�J�?c�q���%���p���Ȁ�4�]Kg���wS�����x��)6�_I��D1;����?����2@�u��B�l2��F�^���u��*�H���R�U�C�'<s���N��0?�@M�n�}=�jW�qFU[��p�?�<����Rȩ�8lu
j^q�{�3��f��e��W����&���\U�SBu�Y�$;絼��ȵ#�k-ͅ�ud֌��A@�р+Ma���\I!��FU��Tr�)И��M�a�
�⣕������&H���M(n�g�;�w]!�x��r�N��)�������-��y��|��Go[<R�X���{쐲P�y�.5�S(��U�5z��sb�K8&�K�b��"��}���I%�3�n��N�����]�b�(�)[R �Z�Y��2K�XJŹ��g�d�T/;���kV{PXcn�G/(L�G�Ll)�����GV�%��M.j���\����I�z��[qk��+!��s٥E}�t�2����t���1�D�Fr���N�_>�!����,6�=�8n�����5�,�8���0�+y8��F��~��,%����ۉB��֔�(�3�-x,�.���Y��A��z��)�!+Z��)�I3����������B=�TϪ�}U�31�VwE��hnA�Y�{v�Z�Q�D����A��j�2����O?�����<DP���W�^l�Ky#)`t�����kB�ʘ���_�x�j�D7�&Xm��{�Ȧ =�.vo�c�l�c��_w���*D�����	C�-���Fsڊ	�Ɖx�k��E:G~^����킨�`�Z98�0a5Ę��K����Գ^��D.��cr��"=����#�𝶍}fL@E�W�47z�dp�V�?fg���'0r;Au�=�ݺ�T$��~WV
����4���Z(��1KN�2�jYx����s�0d�UV;u�/1L����4����_bl'@�xӗJ��nfb�*}���r���Bi�*߰jR��:��5��U���µL�r���z�g��ƁQ�ɛ�r�H;��iR�P��MR�l�_s�s�'9��i��O�����4R���/��j�j�*-�f;>�;0�)Teqɖ0W��6a7�D� ?� ��@�0���4���}RO&�t۪�ɇ�4�>�~�q���@�P6�q$;6�G�l���Z��wW��N���B�~���[j���D�_"K_�Gh�~%�a���l�Ԝ��#Z�ᾯ�[VH�֊;lE�Tt�}��<��, �������Aj+]gd�I<%+V��)�> ���գ�iL ��]��3��pа��M�!*���jO�A�xǔ��ďZ�D�Jh�����e�)�q{��O
����XD��LC�~�`�|��vd���x��P���(��Х:�^�i��ګ�"f �-�-��dm��Ôn\�'5��>���O#�ro�k�����1�9�EJ+ީB�[P�am�In����v��ƛ�%�9��
#D|	��d��W	}ƨ�����{��K�;O�J�g�k@�*����\5����������k_\��g
������;M�� �E$�͍( Qk��4��K�{�>��8wK���F2|��(S�C�QgS�� ��&��Euҍ#��LN,��ٻ�ySs.�2�h�/�K�����z�è�v��z��4k�q����廣�pU�>,݆&p�ƿ��b	�Uґ�Ԕ�C ��д����ҀG�"�T��tL2E][�mE�*di�Z
`P�遝��������x�E6{Z%+���P�]��̤/����~��v�MW��}�zb�\�v8L5ٵμ���A��Y���-��m�K�d�m�C�3�*��:�5"[����%�����������h���p�^�X�.Y�f�Va[�:�~��
�enR.���!�~�U�c���MT��{��X���	:�����8�x�I@n?�Q�a�N��tT��ne��,(jf�Mڨ0X<�Bt\���_q6�����+P2� 1���WU �yT~ꕹD0-�=u�L�N��������R$��Ȉ�Ō�z���	eU���v 3T��n����|cB�����[q�����8˙`U�:��zx������/�^c҂6*X�����X���&�K��3w4�WJ.o�y& !�N���
��VݡL�����Lz଩ ����'�
�_m�E"��v�V�^v�������d�Z7�m�(����$�I ��������.��/�����(9ں{�.�`��{��Yb� ������p����l��	B��_�]J����Qtx��8�ç�r���HF$?Ég$�ӑ~�Sg�.j*�kX=�O���f/��i���$R	ӦTQ2�E��S�B�)뀃3�><LB�%�9�����O��F�E:��]Onm�ԹEo�h�{�� �:$5��*1Y�K��v�n�]�G�.��N�P/:��H��C�UHɴY�y��wF�t�j)�� R��!f$x�+՟���?��a�G���κ�o���J����g�g݆���H�]�w/'�xVS�-�v�1��+EH����X���kN�/�(4w�D���[~����y�Fw��T���Y��%���L��)J�ZB�Q��%�,G���������x�`9Ү�Bxud2�����?aR�/	=V���{,:��p�L�
�Ě�����zp~��_!�ɵ�a�-��B����az��;��&
�p���ֻ�'�u���/�z�	��(��B�(��$�Ok��k��B�/Vа_	�N(���]����Z���f�0I����3����~+���iᤔ�	C'�4�M6���ُK ���=WwZ���! D�]R.dӏ����]�*�|�H㪭���w���k�0(&��tl�|������َK'V�?�3��;мsX���XT^4e�q��@�f�s��-^"�Oy�m�Ne���A��#Uz �ۺ=ޠ��A2��B{��o故��F��V2aڮƓ��>�'�F�Ȟ�l�,���{��h�Ż`����GC��mQ�3O���vJ��;.s����Z	��@��J�L9Pql.p�"0�Cm�2�tyNr�Lȱ����C�QH�@��  �ϒ��+$�<9	��MBV��=�*��0	��&+�C��
�廎`[H�k��4ps+��=������S�7Z߀V��Q!a�9ժ,��� t:c.uΗ���Y��'P0�R;�U�B_R;���3[�Դ$%�J�}Vů�m�q���Q�}Z��g�s���Q�2�WMv�O�	�?�o���a������	i _�s�c:���E2oԮ*YW�� ��*Q��^���GՔU�+ᵩ��:o�yob���g���^F�������+rYX���*Hbߔ)`I�-N��{cx��*^��B��2�i�+X�u�!.�6�����xm�l�Ⴝ�iP4��"
�0��b�ܯY܁�J!�0??�Eu�OEW~۴�P�5U��u��Όs�ue���{fg�a)B��wX�|�py���Z��s�����W�@�Mĸ����N�/�BA`d{���$����@���Bb���a�/3dC����j8����z:�}��G���~�ɒm�uSK����x�A�,�����J��&�9�i�R���)����mBݞ�Y{����;�␍�<h�q�5�#d�6�A�Iȓ�}4�s���\n��
[T�%�� q��Y�5�󆃡I�3��<����L@*|B?�לn3��<�˜�a�������1��;~'9�k�|!�Jo�[���է�Bs�` �gOs�����V[���I1�&���K��f���u1m�<���  2:���|��i@�Y7���!!�H#u4NӸ\��}�'���k�y�᥈j�凙�}�
D=-L(��>�����lWo�f��|��2��@�{>���*��e��
�"���Қ�b���Z6X;yD褲���}h'r4��"��#ϺHg�+:��j����T4u�e#��elN"k:F$�K�c�����j�pn�����q�78�����s�.4(�4A�V��}*����8�S2TR��VnnE���!T���O2�:���_���iJkʭ�%�Dp��,�-l�Zy��/���k������,�T��8�q0El��:<������P�-mך��RW?�D��֙,��$�O�{ۡ��5�	Q�\�M~�p[ѭm�1��"-�s������ԑ���$ʔz��܀u�7?;�CR�!Ԓ47|�>/��3���Nk<��#�֩��&�����>߅D�`@�Ɵ]�H��rq��յ�}2:��; ��hX ���}��6����c
�o��
Pג#`ea2&/�����֞�W���Q���(C�8��Q9� U��ז��f�2̡��fG=i)��L���?�.�F�1�����Ud�w���i?�9R��L��O���ۄm������GWe^��:
�R���g��m;��Lx5w������L)�-)�����$��ѐ�����0n�T�Vm4^)yga���?M��hw��&��o�؜��*
���U�0�Ɣ� �o�6Ӵa2<4�~���x �=�[-���"�u:�v묓�E������M����Rey���s~�i3�/�tc�:C����6̭�6d�6JvrrJ�ړ���M~~��:�ֵ���jE�SC������p��rm���x��a!1l�w��4�~��ƴ�g������*M9Tc�\�H�T����x^��*�+$�ɔ�Ҡz=ߵ#�or��^�v�4����a�ՇZ�7$9�iw�Xk��=m���
˸�6�y�\����V��G�H܊P�|�����s��8������5$���_�� I1�����^Ɠ����V�)���bI�{VV�ז׸�Z/��)H��@U���ٽ�X���	f���7"u��SY�Hg�JDy	Bw�7�[4E!pu.}����e[3L�Y�o����F�k+�I�EC?BR��.��X����\�)�<�u���K�p42�m(���D������W���^��+�8���N8>��We������/wE��+]C�m.�a��ܽ�hL��C�_ܶ33t �,i�"�V���tN�������;S���$
hׅ|�;*R1�()��&����$Tr���ʳ�
a�R�Վ�u��xh7�`��M�aϗ�����JZW��2�����ѯ����EIn�T��<�%��-N��L�lD��y'���\Ɍ���D \�z;�����`�t���5�}�d;ǟ@��(�i�a��7�X?m�v
Ht��%�g��t_듷�|cJ�¾�xev�F���5��r�vs"�6�ᱽ��ŻM��Q�/m��Z�x��44D'^`�"i�0�s�3!�P��V�)!�*v�Z3ų_(f��Y~�{��G��
���$�O'e�˒65��9�0���%�B����1\�g��Щ�U�MA��퉲zs`�;s?��&)�0_�?9i�u�7V$l��P���K��"X4ݐ� �xu��^ԕ�'$�%@w�C����7&S���b;uA%E8���@r��u�	�J�s�@`6���{�� 8� 0y���9�-Z�E/7i,B�	
�tM��=n�V-��No;.����]{&lmKĔ����߬���o�$Ɛ�ߤ�3>o�_N�{a�y���z}�,��'w$'�-��9��]2���tp�����8K�������u����a�Q�:Z�3u]�pc�E	�h&i�}n���#%�Nwߴ��y����"h�1$&��N�璹/�R��=�}ZK0��d�Z2�pK�g;>�	�~��':��\�E:r���Em52�i9L#-�1���Y�ͩ�x$�S��2.;�1����9W�����+C�J��Q"��x]_� ��>o(��v������t��ہT���Ǌ�l?�f"�u:�N�>MQ���%��*��z%����E�YpI�>=;V�A�^�[���wW�L.R�-��#�:��Tn�t�۩�����EN��dG~����'�(�R�]WƇSZe�����j��"��̀�!U�Ǉ�bD�7P�����81��,E �8b	�{���4��ĭ�"������!�p��*�'n4��v�D���= �(�ƾߊGa4e��������}��#����v"�4��}h�d/��;[𡻽1���� �QBmjT^�/ E�.�e�Y�'3%1�콴�-6�b�A7"s@L�B}�>f��0���d��Q[���r�у���I�M�*mXw�fn�gS���(|�S(x&TO~�tc$4�.�St�8"߉�{���C�'݄��������R�	;7�eX)�,�R6�^kG��{�S�k.9�ߪ&L^RD�����/��ԞU��Sbe/@���r@��
�4�'�~��t/X�ҳ�a���N3�3� �t^������I�q���B~��g�큶5�r�
�j�g|�;Y)�O����~��w�}+C��;#�ɍ�ue������x�c�ąh�gcw[�9'R�ZފFŎ�VV��X	E^uT���(����lg�U��oʛ�`�'݀r�>k��hi�q�^�S��}hݬaùة��A�b�8(�T���+_GY	�ҫ��=�9(�m��0MO`Q�ɿ��1_E��7g��!����L�WP��0e��@���R�z�!���,P8E�ߜ�����ZA�Nŧm�/��:��M1V ��h�(`�ݖe��� H�ޛi'ݬDS���3��|�U]��9|��J��d�P���E�0�]δ%�Y���� � �0������栐�I�cݫ�@�%�4b�7�>�"	�s3���
�zHd��.pܴoQ��)!'ݲ��u���'���Z"��&[�����8s��r%��������`�����8ڍ	��{�)P@��54'�r�V<���Y�A3�WE��q���_�O��f�p0'/HR!7$�z��27�"�­��e`��e�"����Je/z���趲�wIW�&���R�㧕�/�&m�<�+��9�G�֮�$V�F�a�b����l��]?�� ���i�!Tb��� ���k������:�M��?��e�~"(��	 �Ƀ��ěcN|ϋ-��	�Ǔ/96���|I�[����O�7m��@
�k ��VsXt��~ga�P���r^e#�6�f�L-G!�����Wn��@��Ǝ�P��'ZƜ`�pv�����h����&<��!v���Ы���Bw��+boX��Y�8Q�fՍ���/o�@�id���jF�8:� ��_9�W��4�v���S�6fU�d��Z��U��{w��:GG�;|(2����"�#?�;b�(�y��������l�~/#m�W��&k���|�3 Qr�lCJ�Zǒ ��7��M�sPX[X��<��Y誖\&|g��;�#������\5"��<9$5�C�&/R�K|H����)�'�oA�P�?�ͪv�a4z��̏C|��O$Y����ow2�"���ҍ���%�y�&6�������2c��Eu�6I��e��R��������Bd,��E3�����umOPс�We[AH�=��t�LQF?�G}����䩧TS���?�P�w�;�����tU9�\�TL{��l� ��qͫq{S��-����9�Os}p� $Gw.ᡃ���=���"���8Y@\�������B��6K���c�h��+u�ͺ
�7t@C~ ��2��!4kTDz�O06��{�Q�V�<�b#�",_`.�&֤�@��?����cǙȲ@�Jt�{����5�h�{\����8�2n�v�[щFXdB����'5����� ��~�KZ|g��{�ڝ�5���zFI�Pj������ͧ�OG�*��,�Y�L�������3�n��쬵i�@�$��l�X��Uo������7˹`��n*����it�����es�QMz#
�}��{-4>�dfF���Y�&��q�`ʵ�_;y�7�*8�*A����
#���ˡQ��..,$�A*2'e�L��p2�J& �;L�5�{�9���,P�F�����Kr�_5<et�&2E�o�)��:��pq�fo�y�Dzw�):D��Fhx���X�P���BU�	xc� ӓ)���SP[ �c���H:xQ��o��"vn��d�k+�'���R�.�5����M�� ��r"��-��l&�˦cf�����&��7�tz8�N�9�(\��B���dV���F@�,���ʭ}!��H������X���Q�A�̡��E�_��G:��O�p�C4�Ϗ�-E�Q�:Z��2l�r�S�2�/�K�ȩ��\b���V��ޘf��b��U+��v=DOh{M�/Ndu_�@��-hm�g%�MΕE�X��)CI������N+3�O�Y�g ;B�h�`I�+
��12Cˠ\Ȣ(��-|n�ڄ�א�I	7ӥ�dA�]=R��[��w�q��i���4����H��-�Π��1��6����Lm�Lxak�΍�5NK��m���m�gI@�xl��O�&�M�d�M�p�#�l\��+����? �'��Q�TpfǢt!�uI�27��_+�*[U$���b�,����9z)Y2��ӈ����;S��m!��iKxu�T6Y�)�)16~�qk�,"V<��s��rc~�����>\_
G��i����W*R�f.���RZ��������g��K@+6�Յ����d4d��
�g?���3�� ���%.]͑��2��~j��*��)�պ�ꐈw>��5+�����W����;:Gخ��7���)��?�����j�{�ҹ�25���򷩝�ؑ�-52����L�#���r
Fٙn� ��ِ6FF;'ZV��7焴�Q�%�B�ߒ��t�4�BEA��xVtF$�>�$^К��~�[���L�Ў�H�i���e4���j�Η��|\��X���5��J�p����B0���˲�a�A��j����UգD�.ʞ���v���+sY�k�\�J �,�u7�=�̿�1��X�pzZ�g,�'׉M����K�7�t̺!�K~���x	���{q����P�~��|�y=bg�������{�q�ıĎ�4u���݀�s�׽�f��a�3�����R�łޭJ1{r���'���ܣiF���:R�Ʉ9����A��UG�ư�l��:g�+�.�9���0h�Z�T���w˔�G��\���������ɡq`�~��ù
��y�OJ�}Q��\�,���(� ��A��R�Z�A���ET����{��v9��W`+�2:�j�i�)`��	8JX��Y��Ǣ.��%v\%�����?/{�KI�3s�V?����[���Ozt/���/����OVpR��ާ��dN
�ꩥ+�Mn��YKE��y�g���'z.�:4B�upt��K��ƹ����$��g�ؘ(G-�b]uqn��u-��F�Lb�8�}�,~�nr2����,��K�s��Jբ�5�'��ɐx��n���q{Q��Ƭ�(����߶a����U�Y������� !CUo  ��n�/��.6C����e�dI�����h�Қn_���~#R��^K���{'ä�<��c�2C���v��$��I�ru���i�r*�R1@�?,.to4�J)3�k�5���H�ŋ\��ܜň�}Ѣ-��o�{b��^b�ح{�F8��ba7d��:�ٕ�<b��h����3z������ �__��V��]�RG�{�o��q5
щv��K�a�җ�c�jiL+I�u���M���������-A�'I5:��$��O�ϓ .�o�\$cΜ�����8{���Ăb���t'UU���vCU�$�?:Z������Y���3�$KݒSM� 4�7Rt��6�򙡱����z�'�!�ޒ�;!��zj������Q��x�V�,��)��V�9}�~����8s/�����#�~��
��4\�t��\z�<�rQ�-�a��#�r�wl�T������v�o�W�<�=]�4����<��}!�TC��2I���?�'w&��6ڗc������A�#LTZ�UV>e�5���H{<�%�U��1A����[�N.��`p7Py��:���j�Kk�բ�=��uS�4��|A����x���<�)��*�N�9�(��#b�����Z1�Nt��'��0g*Y3��r�7���Y]b��WX�@��Q�*]3��=UD�hz���4�I�l�����nO=��2��u2���Cc�$'B/�����%�T����o�h|4���f��`��%d�M���}Ո@�Y�A|����!:	a�HHV(GmR���Ij�ca������ke�#��=�b}[���#���H��� ���,ɹ�Z�ZU��	�:�=9lR*�eo?q�T�45u�4��q�1��f�8?!`���Mw�'���SvL@dM���#�v$�=�]��� #&+K�L]����\�nӨ~��35ϒv�B�j�x�̥���y|���H{Vk��9	����i��t�Sp��*�^'Ҁ���%��\�vA�z^o P@)�+;*�}ά� �ȁ>ZoR�*~(�!$)�le�|��b�x˒���@\m��
����_
���R�Lm���_A�:�<�w��r�	V%�B���R���y�<�p���6�R3�DfɼX��!:��4���&[��3��t�=�gAG;W�`�6��b�Ӛ��C��.6���-
���H8�%�Ɔ� L��y{<Y�kB��}���n�����F�[CBTɟ�}��E�V6�J�eRl�:�7�X�N�u��J��-�_�N��w�F\�H�qN���fe:�A�<��"���Z�*��hn��4��!�O��j6i|�tyF����:�&��w3�A�=,J֏U�S|��#�����*��F�`�x��m�a�uQ�����8����e�I� w�����>�#ZTH�G��,b@wg��?*ݚD��ԑ��@<���6&�^�UJ��q��a����� ��~=5��8�v�c�������}��A�v��ANO7��� ăڴћ<��+I
L��7�-��`�#�o�I#4�
 ?�/��i�\�C~�x;�n��}�>���4���ų�W���`�
jx��z^�n�u�
{%��_���~G-�t��x�� 9�H< c���0���|��ѤZPx�۔��$Cr ��+��ݥ�n��w��΄^JD����i�`��Y�%u�bH�N������]{��=omZ��Q�}��7�T��
�#���*J"��"._�խ6��y4
��n�J]�{й�^H�$���ȯ¤8�¦W��R0�k��)��SM�X��W�N���n�(�Z��� �Ɓ�6G({N��
znT)O �=�dr���h��i��[�9�"Ƨ��?,���k>�@�*R��2�e�������8(��:�:�]� ߦ��ݘ"o�L�)���x�]�N�����P�O#�|�����z����q��!.s����Q�/k;�5t��M�����*��X���((+?Ğ���N�V�}+��0���Ogy�ߕ:��������ym���׳����EKf\ρ�����<���`��l�lk�έ�#/Z.k��HM���}����s"�E��E�������}m@pJ���4Qz�7zv��,rWC��y1��I�����\�y�1d����(J_&�&��3N��ض�VgxnX��3�7��u6}����>��.�֌0��,v��(j$��3�a����/�����
,����׫k�x�[s���p=��[�PƪP����y3�G�'h 0Awe���Y������A�8�����2�"��l�˫]�S�+���d�hN�Lq&�u�6Q.�����E�f+M[SyzVN�ڰ��v8���q�u�h��JXI�����U{�V�R�22�L��`D�5T%�rO1��c�X�D\F#LY<��e� B�ZCv��>�Y+P[s��Ч,�=0 �ll���77`�R���2JyT��5����K}�������f5��~؄�A���.��l�@�&��`�/{�&���4� ���7�3��g<C9���
X�Fv^f7S�Ö֖�y�Vz����I	&�����)@$����$������gZޕC9c��C��v��3�j58���B��
�-���d����*�w5J��4M1X<)q��L�h�Lb���<�I�{�=0�t	�zhq����ZBǮ�	�b�XD��I9��E�Di���u�T�`�������@��C���v���^G�RD��=B/Z��}5����B��S3��W�W���>a�}��6Ҫ��Al.�R���-rC�35��}l@�s�L� 6+�������g��8���a\J��r?�$��7���4���dxS'���isRm� �{F#$ۖ�� ��:���UJ�����Uq$j>�8�d�1��������IW�3�j��ڹL̪[��%�� 6���L�u��a��[;��e9�.�;}U!��Y�"4ɟ�q�&>�O��UY����{?�x�Xi26�Z5��Jۻ�z���Q��.��ڊͦVdu�r4���ݏ2�h�,�R(*���V��V�1g�&�����"�j���f[j@=ݣ�,��ܥ��f|�U4�����Wm���"�-�7�lւh�M@���sEmu8kJ"<(�(泹�9m<��''S}��[}⌰5y��j(k*$��HH�� ���I!���d;&U����<%Y��w_�lI��lB�$�s�@d�C��Z�7­Y���c�#L�'�&�^��&K<u]�Y?L�'|T΋e��!���5��>)jc���:�A��as�r�FȢ�s�;!��a���"
��QuqA>�m�j�p�2�T`ȳdx�'wn���P����p��2^7��shҽD��KÂ\(�,Q����.�#۞s;g����ľ���*_g�g�B"C�N��Y�w�B���"o��{wq��/�>#N �\6�����mף[}_x�M�1-`�[�A���%��E#�<{���y?����ܖ��!��oN�Dݍ��ؘA��@EؙBG����a�omm��v)1���py��ЃIٸ<��p��YF��<"C(��ҹMj�]��b�y�Ik*�Y�f����8=銲�RɁA߽�}W���Pđ�!-B�_��s]�D�k���
}/�^Hiy��8��.3���h�]��*,�&��7�
��Ѫ�3dPf�o����l�2	[���{�6��A�R���lHN�`�Z���d�<~�f:��R���h޼�"Mʑn�������O�+q�����>�|���RusPc����k�0E{v{p3�LD���E�8:�B����!�_0�1��ٕͨ-�},�\��
_<!	4,�:cv������1-���t�gs�j���Y��eDI6ȡ`�g����ш���:�pk�� aN�^3T��W�P�����3*[[���$So㿃Zw�ʚl5aʝ��L�]��ݨ��tk4���pn�� �n x�����\,Ϩ����xZv�ܼ)�ذLv��60B����x��bc�%SqS	�O��B�n4 ����;#9�N��CS�ڢǢz[�3�A�`���9����
���'P��	�����h���<B ;���)��b��ze�4���&�.C��܏h�L��v��z��U������eSD���=O�_��]���!��t�"ٜ�%�@�8
ך��&y��y���v5���Uh���'ϯL�\��7��sr�܎2��^�=@��>��s.>x7�b5#�RxP5&��z_��4ET0�����3�"~GmXT�rc^���^�����1��9��ĪjNI��+RWPOu#��P���;�K���fho��$�Mݛ4Vu(�a�a�x�:�"K���c��^��G�6���;�6bc�B�Ga%L*�|�	��q�L�SMU�W.�G��rSW�#��jL�`(��<�pM�2l�	ª>@x���4�2�Y�B9t��dd�"� 	B�Uo�p�	v_�v"iӓ���w(�˿�$�A�\&�U�1:�q�И�>�Nz��,�6�:�Y�;k��I�
�C���X���
�Kx��4�c�_��J�dU���.���+~������l�+�� �� �x�T�&p\M%��)M���M��`��7�5^X~�R��d��ś���V��d;]>tj��֕�Ѝ�u~�������Ȟk��X. ����J���F�����TU(C���E���e�[�▯
U\x�/"��'��?��}��O�=?��� O/�좏pWŒJ�{�ǡ0��JR�q�����xb-q�Ow�ύ�[�7_O��D����+Ȋ�� �I"5�M��6�r���U�V^�b|�a�F�'20C,&��Bf���M2���	 c�?�����H��BM��B|��A����kP�k��XwU�[w���V(X��|�ZR��CH����h��!�S���&��[��6Ia�9�!� ⿗GZ�6��M���-��5�(O�n�{�e�K�ՄFK�ԋ�ы�����f8�R�T!6#�J4b��M��N�*�%�9͇��m_6Bo5!� TPE���_;��\�d;�� W~se�2�u%��ĥ`x�+��n+^[�\�V�
��!��=@l;�H���t��_Լ6���Sg�H�N��e^�&{s��i`k�9����M6-$�$��U��E�UR��7�s�Ʌt�����j��L;�/<i�1�Pk�&۫q�	�����Q�e�{��8qh��}칿ʿ�j�3MC��#�"P&��>�V��Ҕ��gY�I�:��<(�w�P�]p�a�u�x�H1�q����V�V�@���:z!�U���Z��KG�<�S����l�*�������/�!ojGXZ0{��Yll��o̹yBsT����3 K5��<\�
�C�ܧ�D�\:�(���XʗMҠԤ�RX#n]��O���!Hܭ�e7$�f�gjS���ޤd6f;o�5�b�x��9����^5fܳ��w)���Y�K�|S�`n���ja�j���t�0m��>Duk"h�6[�{�QJɢ,�sT���W����D��p�oC�����������#��1��̦�)�K,�@9�lc{�}���F��F�ߩ%��MٹWI|��z�*|��u\��\-����;��I�My_����a
u$Q�#(/F>a������y�az�v
��`�fӈDH��z��>����B�V<to���!�D0�[H�O�"m���:�R�x@���<=�h"Z�� :��3��(�G��+]�O�@jx����~��Ɵ�P�է:�#�r+o�PW�0�l�E�ޢ�IN��w|��-�'�Zs�U�l����*�id(H /����Ӵ��i9�����e^!t�ޙ��&W�B�܌�.ܠ�L,xK4x���JؐE��� xGN�|���;�h_�x���Q�@���S��w=���������V�
h�tULNG_|=�(�IX%�Af@��L.`��>ygGE��H��THpө�����ϒ��̫�Th�s�>!�szK�Rg{L6>���j������8��"������������BAn�3��8tX}h��z�1`ތ*�&����x�^�M�-}:��P���f.U@�A��u~g%:~�Un���U�����q+����]rC)������Q�oH6�7��,��X�u�_���l���KYR�����T����p�~�s�0��+ �n\Cլ3�ny'SY��vO�h+}��̤ �!UA|Qw�4�|�6��V����m"s��([�#EA3���n�]�[T_0������'"�;&#����������Wԯ1�]�s���@VQ�dz��x��l0g��2���}H+W��
�D-�WJ`���Z%�E#�7���b����5�b�@��ր�����r(����NJ��7	$oa��ia�;�
�E<T��E����6�4ɯ�Mh���;'�ԐJ���n�պR)��p���������q�,d�[7�oJ�P�l_���� z,K��Q=�i%ZE�ұ�������q+jq��Ik�Ot�ͪ�N��6-f�D^��/� }���E��e�'ϳ+8y�p�ϻJVD� ��Q�&+i�����jӺUI_��M_F�E�<��~)e'=>��;i���+�C��G�h���-���d R?��	$ճ�*���:q�Sb�}}��B�����h�l�8���~����ʖI�
�-ܾ�|F͡�u�F���!���J�w��]
%&���z�3�Vp�8�3\�0�aJ-f
���Ce���N��L/ܨ&�%�H2kX�q����������Sm(p?.��c{bil����'<�oh#�HKՌd��ka����߄v[��r��쐒�D#8�VS�C�5�+e�8a�Ѭۉ?;j.�r̓_�jsc'Di�m�A�G���U��K�Qj�G�̜�E����_�uV��Kvr%�t�h��%��(������ ��o���,�`�b���Iw��ϖ^#u�N�>5��$�"�঳�|A��
���y:��]awY#x{k�v�?��bj����c�������Ԃ�Hz�ق���C ,g6�H�:'��+����ԋ�~w�,�aw�5\�.�n��_��~n1�/ lG�����'<E0\� ǟ�4����=Y/�R�+�%x�V�9y���k��oG�*
 ��"DG�m=ny� b�x}�X�r�r�b�u;Y\McYɪ9�$y[˅��W�1��n�br�z��RC��}I+�u�C�<;���¬��:��qXX	� 
�(m�W�]�(����gh�[N�p)I�F��{A���L3�ٳ��۸�[h�����ה�~.�j ��5��c�
ʹ��h_?��	����Ɋ�d�A����Z�u�ľ�
 ��{ �i0�I@��c���|��ϥ;䗮*w}��\���6���
�B��B�\6\(-Q�82-i���y|�@�����>G!y�܀ە
��侟H�WD%M�V��VP�/Od�&6HJ���_�C4��0@
gp&���p��Uu�_��Ʈ��$ �X�IѾ�E�ue���"�(*,��w�-�T�_T��̱�ԍ���g��W��.��>~�e�h�� ������������~�*|+��Qm�{�WaG)�G�NAL�7,�R�����}ә�q�m�I�؃;z���6a*�'��
���?�����Q�V<Z���jc���p�囂�N5�Tz\:�����v�\+�P����t�ӑ�[�b/��`�U���is�u�1,[^y;QdV�J��U]uj��7ʼ��v4��.��4�[�,K�:��*���&Au�\�(ħ,�jx��b�W] ��_��R��Z����>uH��P�����^���j]��R��{�����{�>�h�L���c�}�Ġ$�[�(�6�⌋�p�?[�L�RR��@d�m�����Q5Y|�����׾og"rf�t�ԗ`v�H�X�n�v����&�K7b��:l)l��s�Z�,L��x��wEU��,m��"Ѥ�N��F������[�u+��W��AHYU
��"ۿف�u�qh���Y_�=)��4SM��^��6��G�j���lDX�����ꄱv��T��z
�zw`�d����2��q★�^u���E���mŖ֚KaPF�*��\�����cc�`�(L�k2��?��m��k��-�&�l�f���/���&�~M5��Mt�m��14��� W�a<O���@�P��nQ�_���`^�nZpj�@�ůD2{/����uDZ��֝N�Wg�_�Vm+5���`8�fa�"�p~�䘀ǝ%�HD^-���	ӻxդ�_	k����ň(����(�!C�<Og�W�=O�fU%\U豲ܗ!s�C��T��(��=Q�ޙ��\��_yF�!~����e����]h����r�D�wX����﹩��"� �2������^�ڋ�N+j�P\�3���g��;�ژ]�"���>�m�Zݿo�gP�|D����eo�;}�7�7���H���@�	%g
��>�,����	�;WK��C�EP�e)�'�5�uh'K�]e�[1p4��o5�}rd�yGA�p����"T��c��m�u�S;���d�=���]�_�g�D3�?�5�ʬ�@�D��h�:ND���}�?�9�m�$ɽX���[6��hARn �qdOE�W�y ��LU�҇�L%ڔLm0L�hy@���W�{�j$ؖ�5@u'�/l��_���~y��%�n��ձ3�UV簆�^"M%ywX��d��ߟYv����Q�G�B�,F���9 ׯ��H?4��n����|Ӭ��^(g��4E0��K����@X�dկ�"|�^vW�M��7�\
��,e=P?}�1u���d(��5�_���KY���u�	Lo�������:��1�Ic�_^�G����oO��̃B�6��
(�5��<ThS%��z�u6�ˌ���!������;h�gd�r�� x*#SOM�K�
��`�r��dԗ{ا��	���+T=|��Q����$��%�p*Soe�QhBp����&d)T��N��[Dp�F�^���8O�q����$����ௗo݌�[�%��k�� ���%*V�R��"w��|��Q����>�a�j|EsD{�F�n<����E�v���n��1%#��L�_uO��g�B���n��%�ʟPmu���mҭ^Q�����,�~ͅ!�&�,�5d���av���iA�4�sT�.E���d��Ɇ�y�7���l���Ӱ6���D&i|�}�A)p���1c���^r��+V�AvU��̉��������.$pA�i�x�;Y8�������p�dgp��>R�
���@���N��D�V<5��_ZS�4���=�L��Ƭ�F�E�����Ip�} :����M~�\�0�q�'?��&"ϸ�Tߐ�	���|�45ɣ��,E{K����3��}RlR2#�墰H�	f������A�"�b�g��Vt��?����ӝN��W��j��s�5_�� c5�E=aU`�3��U�;
�y���b�^�
	m����y�V�
�7)�f�єL���'/�E2�聃���M]��Σ�> !����[ͱ�}Γ�.�@� Ș���<�	X\z����V�$�Rڬֹ3���wA���(B������ґ�ic��"��;�Gі�PM`?߰�Ќ����2���\Ҳ^�2c����D�d��?�hrl�$#���O#�/��͍Jd:5��޸��Vxg�u����t{�ی�R3�@�t�2�5-#�(��a��b
C~x�֭3".X���B1�����l�Qr4n�Tt хۼ�fРߚ�V���;O��
�[䗦a�.m	j���k	yC��8o��	��+�ʔ�~��TWV?�� �f�{�}O����'vHZ(`��s�� �s��q�����Y� ��i�Ϣ^v;��:I+�y��d��!2���_�ه�%�iO��0��/3���\&��}8�P�oM��ŉ'Z�)&G�d~����Yݗz�q@���%=��\��j?a2��{�R�����.V�*t��{�'X�y'N��
�7],o�G8Ъ���]���¹�KDh-���Y�p����\#���L��-��ڿ�ǳ��'P�B4P�\*����Q��B�CZX�c=晚iʱ�زսT�1։KiP�G~SP;`^�~�dw �G��d��N�4���[>xD�-[;ѭ����
�#���[��Ti�'�Y�����MJ.���t�̮��Q^�}D�}�`�*���S�-I�w���Z}������!i��@��Hw��	���-�1��)��&Q�֢�.���� ʥ�(^XѵȻ��9��F�߷���g��g��A%�� /��9��a״�5�Ѽ)iq�A ��Q����+3�.�h%��L�&��(�Y&��`�< R����h�hk�}
t(*�����8�%�������#�Mٚ���;
�����J�n"��!�셈��;*l�:�;��sޯ`�,�Qǐ5�<��CFF�ill~-�(e�H�E�)����S����j���q\�}�k;ф�ߡ���Sߗ"�9����\����\/��g��o�^?��Ȑ�]��R�A�&�Ӕ�oZ�)��,iI�{��\�B��a��a����z�!]x���t��L�EM�bě�o���M[b�n3��]�����B��y�Y�ʦ9"��M"6C�����%����}WL��qZ�\�<��_c�3�{=�Mb��� v���cx�e��WP��'��*P{B�=
Xz碹|����C*��A�䑲6d�K�v+!��x�ݮ��uy�����ϟ��D�
ZDho���/���[-��"���8$�q�9v���\���$����B�	B�ޣZp���HD?Q1��B`�?>_{W���sZ�yѼ�D.f�����H-�Sp#�S�aRJ�����I��Oeg�~�����.S��9�j*aP��8W��1�[���ê'^\ysCjF}�h�����i��2�A�i�)�낲`�;Z��ٳ�7Ҕ3��꫐(��e�ך����k|��í�]Ί(��ʆw�V/|<�Kĭ�騩�S�u�*WA��)��*�;�iD����P>y�,U(_�)�V�-���%xS���v�4�
���{�F�S�<�H=�����Jo�����DW��w�t�hߓ\�r�pn�읛�Mh���Bq�ٖ�8��ʓr�6"��b�P׍�U�Օ0H�?c�4�BYl���>�~���+�#,�ң��tm��$VYŀXU�m;��^ݠ�O�^uB�	� ,#�=��T#��y?��+x[����!z�\�Q�pIĉ�A�3��8B��ڭ�=}�z������8�8�'����b}EVW"d���m�rtL��m����oF�����\#�h��cG�xr�����Ѡٜ�Ό�~+�N�$�FY�0�v쀳B��lZg�$�l�A���%��IN�L	>yiM����8� }�6rܟ�3�SO�{�1욝�9��0�h�^�N�uXLiA�:�	�&u��2k��4�M��R�=�gu6p�pY�;�F�/h?��)��M��t���n��D��RT�����=qAG�9K�+-���:�-~A�Y҂h����e�G�1�^Z�.�T#<��`�j��٥����mx�GX8	e�#6њ%Z�����:�O��^�0�u���JB�X�ẉ�R�uDF����\�+~�">P�neSAd�̔p�e�\������p!�B�?G$2�S܆�<�d�YF_=)���F�Y��\��.��u�U�q{��DY	;{�P� *����.f!<���V�>MLb�ʵR���`�5{�3_ϯL�������U���<�j���$}XV�C�:����^�8��kE���}{�Z��a�x#[7�g�I���+Ҥ9_��WKB��5'(��Z���x��
�I��I�s��&L�&"[��ɰKѵ9�5q_4U)]!�,��f,��8��|؄n7G	�y��>��B��%_���0�b�ô][&��׷n���#R�ғ6�v��Al8�dYg߶&��ku	�G�:���ՑA���Vʳ�i�qX�J���F 	w�;U�67.��@�ъ�׫�����Hy){M���TZI�7'W�XM�L*�:q� �i(&���%�{9�'
\
��1��_�f\W���$�8K؎��w1B����	���H��2~��� $0��@�v���H�١hVD������˻�b��j�`�3
�ƃ<:١v,�;��))Q�y��z_V^"ε�ǴϪ;�۩O�󋧅�4���c��w����EE�J(3�%��0}R �S!���jB�<���ڋ߰����q�Â�Q���<�S����W)�q.#rl��3��ц���%�ÈbJT?�h��W��Q4C�"��^�/Pp�2�X�\]N7�_�o���AN�I���m9�u,����mix"��C)���K�/"b<�9޼�H,/K
�A4٬��_�ZyQ�NJR-�� �Ƿ����Ƕ/0�q����`vɞ�e�-�� �G�����3@UG��3s���kAb��֏
�A�y\�2�0�{�պ��H��#�m�b�S��G.��U�Y�6&E��/�k�~��ِ�\��?���A$S�--���QB�%�^�?K{'��NN�9�"�"�f^&�5cW�E�!˧�u�=aH�U��Q�@�o���"?��}5�L���C	d�ľ�}nԲ�rpPa����۞h�o��0(R+�ktX�Dxl�>Ne���T�X��:�,��{����]��@�5䉔���z�/vÜ�����i}��KX�=�u�Ē��,������M�Ҫ��k�b=��rDV$��N)p?TN���`�1�+�Gr���1E�a�+/���#Cz�<�-�,F?��K��y��y��S���L|�h�!čP� 'SHb��[�5��c�7��K�B��V���ch��>v��:��X:z��W�?un�BcY�I���=���k���s�t����|h�H�Y�z�������׺eCz4����w �ȗ��w�-MqH�a�V�/��B�
_���?2	n�k���p����5g��(3P���@�H��sY:q��f���ƴ��Q^V�~����Y@|��޻ �\sI��KL{�
_�g�k���<4�.˯����{��V
�A�;��QE�_#���xU���/���Q�n�3���b�[R|.��Ѥ���=���<_'R/+��ш6��Kٮ��ڹc4�<,/�J3X{���0 ��CXA�I���!G�zT��l���l�fv(�d�|\ӿ�n��w�oG��DkpE�鳠�� ������\�3H�"P���E�P�>��0�j��!��4���$k65 �y�w��}zR\�cN��+���	p@(	��jjtE�:Zϯg9�x�γqp��#�۟˄�a��� �壵��D�vxBmBd�Dw���<"�Ԁ�KU��o�]7�zT�vG�z�+?����FS~��Z��B &Ҡo�f�1�i�>6(%��c��D�cQ���p�\��^]a9���P���.U��MG��Q�Z|�� u��έ��U�:|Y��x����~8�*�}r���Zm�e��Ҁ��h}_dZ��u�ѰÊ�V�~�S�l;+}h���5��G{#��~S3Dyҙ���d�R�h8��ڔtV��zO�8�`�����Yf�0��'?Q�I�`G����A*z���I�Lۣ�o+8�w���=,�Ww�� "'����e���f'�u�A�6�ۑ��=�@�1����^U:�b5ן�-N��)����j��wk��'�)�r:�\O��w(w�_���F]+�]k=�T-�/b��zՈ["���]��S������R�a������q�>7uv���3�^gP	�&�Z������ީ<�.�|*��Y���̐Ey�!U��]+t�Ŗw]����;?GtoX�U��5�傏��鴿�����!$RCS�:�8��Y��}Y��1�{�:��7�~�N�_1)m!�h��a�&���8U�Fj�%�c��$ g��������GR��zx��ʫ�е��8�ӘLn���>:q�.*��Rv���� ���ߴtmw� �+0�;��`"���X	����ЛN*�`��ՠ����Q#<s�V���m0��{��g���^��ĝm�*��	)�)�'�����U=,ȣ1r��E�
�A�?e�� �r�����u���d��@2���x��ʺK�6������K�����KL2���V��N!�)a���ŧgZ��s���e��GRU��������<�.�1k�@a{wY�m��3hFUH[�U���
4ۮ�tN᪱񍐎�A"a��N�ܒ���3�ʴDc6q� �^��"���تDA	35rN��>W�>]�8�W�~�����`��E�o^�ṋ�V�����l��a��bh����C����c,�L�I��ojp���%$�E�RFt��Ċ!a�����đy|�6���:��"���&+3.�dXI����&�V`5)jI�"�� ���g������)�49@e��Ӭ-;�~?K<�8�gB&���oD_ v$��ĳ���%
������_�}�ҍ��E��5�/�nE2k���|?M��!~�J��yCI{�Y��B���p�7�!�㳷i�w�q}�r}�.��Vn�V<a�+u�9Nz߇\ƍ�(�B>'�_�R�Ֆp�D���L 2�+ ������t��2��X�������F�7j��U�5+^�w$�FP���l��2C"����IqY��K� h8�j��C��>�F�,.�kc� u��;�g�ZC��;�x/up2����@CD�T�x�&�m8����AF���&���*��s0V���O�c`�U���h ϟ�%3a��I�����řy�A��ͮg�9K��j���\��t�w���AUGf�������Z�"~xK:�6B_N�f<��e~'I�7��l̕
1�Q��^�;{3����G��/����l��Ӿ´5g�*'(w�|(7��S�ݑH�ѹ4^W �Tg�����, �5���G�v�GuI50J�Z�r8:/��r��6�BBt$���|
�[�4��כv?_um*�K�bg� S�2��	ף�F'9\*a|,�P�p
 ��σ����[J�2�9���3l�g��th���՗��0sh	���H87�G���_�#�)z�g��HY��A�]@���q�u��h\Y�f��S�c�O�+��쀙�dӀ~��3�_�f?i3��4S�uLe
���w}����-��� y�%�H���<Obx$��C6���?^��!����f�a��w���8�Q���g�Q����jBh�G_�aH@�`x�5.5�힬�Bp�X+�����E������+�t�l㼊����Z��O�C_��T]�i�����1}w^��M��C���l����O��^�)�;?����Fa�Vd�QF���HxS7��"��B{�'CB�Ϟ5LJJ����\�_:�H��9�����1��SA�ؖ�ѯ>8�����?�x���)��V$b��g�U%5�b���Z��I�E$x�G�m��8������<���^x��s�����Zm��ֱ���$j�~� �6/�jB�,�0�{E�y�������>�3Z^�����������h�^}/M��}�-��"���q��h-��6Ƀq^�3Hs#��@�pSAP0u\��W�~E��̱�_�f���vN���Ct2��fx�{��ñ��X+S!>��ɣ%9l�����N٪/n*F��J��9�Dt�úoӚ��� �# @�C���ì`'��}�M=�IZ7LP���R�$�+Ǽ�0@�ewd�雝ɯ�b��5��ݍC��k$��0�qCO�{�<���r׾��frP�(zR��J�X�p���v���
�$��^�y�sy��~	*J2j�rctc�,�9�v/���qL�J6�����&k+����vT �E,_a΅���B��x�(�|��,�c�U�b-�Ǭ�F��ma����x���TI�#[.M;����H��_T�jA��>��U5��i���6)7��[/3�(����p�c���3��!4�iɍh.�J*_�/zlD
��..��\ɹ���E��E�n���xhp�������A�azm9�db��Y�č+�$���S��(��˚x�!�Ķ2��V�ڄŘ'����5����wZ�(� ~��-�����WG�x�C����<�zT+}sɯ|=ִ���]�Tq�{���ޝ��������	+c��-ū>'�A>�/Q�o���QӃ^�l�����v+�j���g$Y�C8v+,����N�N)f���~M�`e�$������r��$L�%>hcr�tyn�t��R0��z���� 
�%��N�����Ch� �����X�W8�*n�s �x �)�"���8FO/��\+"��*�^�%��Q��.8|� �C�<E55�W����oA��0��U��^N��m���E�_������sg*n *ѝ���{O���nmD��B�l�鲜n	��>$UBs����^��Ԛ�K��Q���Վ/�:Asy"�SJEh`D�a�����K����Ì����D�<����bY$�ۏ��~�f��f�F���o#�-4Ԧ���(4�.��|�&$��R`���
ݕ{;��}b��׀��*+᭰���@n9�� ��ǡ�L8b��&
�gZx,���^b���I��o/��5��|*�k~���L:�]#�s)Zl��|t"UG�~F���� ܉��Q���^��~�}o��2]ҏ�4[6���P�&�u+�G�݀���[��1I�W_x;�D��$��4�M�����d����D�K�M<���Vz#�Y�mi:�[��@&�&�6���L�>x弆��}U�6x-,��D@$ڥK5*�nW�X�,,�w�]5�Y���̘�����[
{�85v��/~��� � 9Y �q�u0\:��7��R��"'�cp:'�y�6H����kz�k�{��a�`����V�X��\�z�N��� }�؝G6yg��R�7��f�C$r�-Mt��~1�VX�b_=������I�0lSX�Kε���@�����ˊ-�u��Yz#W' @X��r���Py��'E�v��
LE��ز�3ף��#���K�m�"�0e�:Q��g���E�!c�1����T�~�� ����m���r� ��k���gsU��sO�19�?�Vn��~��B?ߒ��m�|�c/�5��x�4���|������SL�+h}`�zDZ��T{73� E.E=� �zz�i��T�O�dǈTlLg�F����"��턲�p�MR�ԉ{�S�}��#� W��������}a��ɐ4>M+ϫ�a�L�S�S-IK��\���]۲rp�Ϳ��`1���Ɖ��$��?D��+lAd�oy��/|8,l���y��z�N�����ã%D��q�q�W�M�� &j0���(	�s5e������
�B�� �7Lx����M�{���
�R`�0]vNp���g?�+us�� NtE�)�'I����d����Wl4?"�J�.�L�=�R�m�-��"�뫋��~�~�����9����մ���}�Sa#�:8d���wn#N<�/�(d��2���D��0���&_�(٨_W{"�z�-�����51R5���M��A��b��S+��xU@Z0�	�|�z�q�x�=-�Ds��)�Z��"�꺠�[��m�+$�dWn\(�̃�;a\�ӽ�h��{��{�t"�Y�g⤁9y��L�2���iN��'roK<u��tc�;V{kMz���%�i	���ٻ�=YC��b�쨾qtx�%7J�ތZ�`y�M��lI��`��n9�.>fY��
S'۸�D?�_2XC���q������Y\ٯ�qՈ�t		˔
��a�!�����%�����< �k�LÏ�gU�#fC�;�G�ݶg�,C�P��(.�W�;�/�B��f�:;U5tq�r(��<���|؇��,od��hT�.Ԏ{x��峮���`�N|1}��G�� � ��s�����'�4ܙw,�X����d�JWM��3�;s�gQG��#R'�>	�[����ŗeRn�����|�k��%-�Ж	r�SG{����qA�pҹ���`�x��c���#Z�p��Indl+]��[%+�Z3�(�XE����kԦX�:;T��t�������5!�����M�㥻ԃ�@��qU�Q���I���8�S(�дFӀ:������_��`�珺���O_��GB:�!G�z"d��s@�@o,h�{5(;��fQ�Gك�pN��f})*։�8��V��apN�c�:����Ѕ���{�r=�:{T
�4��[�dCJ�U����{��L��i�g��B�
����$�#m�Ά�f_������&�&i�~���_�xg�w�²d�2F]���%��MGˋb�6���fe�It����_Rd>�Dc{�I#\�BQ�*��������|�%�%g��(V_`ڽ V��(k��_x"p9�00��qU��47�bͱ�*{���(׶�aC��DV*��$����0N�������{�`mK���q���fR���3'UlBᤅӃ1���_^�^����-�yL՝���>�-�-b��gDu�;�5mi��=������Ah2�X��9����W�vz�#z��Po&�N$�e�m���9_�:O�;�T; l��'4I��L����(�+ mL��b�tW���(���au����mc��N�g�8�Q�����	&~|_y�=��o�W�K�4�4���9������J�z� 8����c,����.>�a��	����=����(�߻����FKG��H�(��zOO��-�1�9��T���)	��ڈ�LD}��ų��

��#=�Pé�E����P`��<��Ko"+%^���M��kY GQ�9�v�seC�1�C}��%�-P�jm'L$z>.	iL����BE�8�t�8\���;��KO;�a�U惓b~���@�e��@F�>�b�L�n�����B�ȧ .2��M������<v��r�v�T�2MHnF���B��+��$Ñ����X�������n���hp�u\I�U/�뾊�#&�gr!%��t}��oJ\a��1��*�P�'C����.~����UhJ�g>7kފ1V��d��Y���z��J��w@i��$����;ۮC���;/�����g�͋���Lp���~�o{s�	��ς�tb7\e��O��sK_����������tLHx�E&`��ݫ5FC��$HP_�"�rfN*y�7�/D~������N�}~��^�����\�T �%��rVl�#�I�p��LQ�V�4��W�R�\��9��C�Q��m���pW�T�PR���B� �EFc�������[p�4^��#G"�8F�����m����Y%o���8��z��\߷�:8�>�,ZY��\�/<����U�y�+�<Ӧ�إ$�T��ˠ��EkJ�"°ԍ�y5��ޛK��fF�7$w��&��<�_�T^��B�@�Oɐ��%��f=q��*,���q�V���[vۻT�~��Y�jHȺv�
:��I0�^�D�BC V�Zx� £s����5�_�q�)�����fga������Q��8O)�� N,&�?�`6�*�7G���[�m'C�T��'����@�V[��R��/	짝��4�"�K�������X}�N����;��6��Sa|��d�ۓ�w���{�H���D�ޙc7��P���l�gT�!З
�o-�"��oFxT�[FP�U/ ��=������ű	L�E.����t0��5��{��rP��Ѯ	�Yc�lS��u+͎�op�*J���xD�~{�r��v���G��䡁�X�G���p!�!�R�bZ���mǟ�� 9�-$�ж���=	�;}�?Pz��9��5�J��Q�EN� C�ʙ�S��_6b���W�o��j���@�v0$�&������Tc�5]Ԓ=�	�԰u�jf���x��1)I�
x�&�r����"Z���F�l���z��߀��㩢Af(�V�ta�d��	�6tD��"CJ���Å���FF]�90�E�	�@�1w d?���>�Ȕ�w&$Ad���6�,���ݘ��8�ի��_��~]W?
�'��b�W���)"�e a���6g��E�y:���j�)�s�Ց1����aV�#8~�:��2֣�$Y��eɹ��
��IN��ȘJ��gjҩD-
���.�#��7�� u@|�p���Cףa[��62y��{��|C��X
j*��&H7f�����pG(��]�XY�J٫�%x��gy�E�i���b��#����f(�s�~�j��a�W��N�\���Rt���z�NE��ş��w�ԀwOU��x�N�xM��+��m ��9�T�l])ȍ��>��A�Rߗ��?_�U�H���"��t�9��i8h!}��2�������%��iY13cG�^@Zͼry�J:܋���&���F�����uˮ��?EV� ������ �Qw4�n{-2C�K����']ͥH?�EX�X��lr�h��Ӽ�!~9�?�r�hh���A?~^T�Y
���c����}.��E?t�_4蒩u�ٖ.�1��8ِ-�'��x���ɞ!�_���v]i�L"�p����M��e��RF�0�̦�	�n�� �P:ꮤ�yZ���!�9>��\�����Ÿ�����Z�/������yQ�x��+���3���8{8���<��Sk���nn���T'.��������9�����H��)U{x�uZ��T�Q:7ͺH)�Y�;�|C�lř���F)�=[#���܋��/���8���Lb�v�s/ꙭ�(�I֊��g�W�L�S���s�k�в�
�*�[�5dq�o<P�R��=�g?�J �5.`ӳ$!$e��^�4�؛�+w�3%T����>�+���3+�h�7�kP�𼛞(��N&��^7�oKA/)L�I��ck)�y��,v�U�t����[l���4�
�鉻((p�$�lr8�A��SO��I�ȞU�4�q!Q�]�0Аz?/H��`ƭ�ƍ�?`�*��G;�\f�1%����zAI%G�#�n��u�iq�s��� �?��opṉ���a{�0�ɍ%8����Q�jh/���g�*���s]�WT����� ��.���K� ��3���S���跆t�c�A��6#3���{q�6���[E�(I�\�-�G�$��~E<�$���u�9�~�3�\���b��i����A���G��`�$��ufٝ�&1<�^5�ǆAx�F����i�"kkW?��%�B��Q�*v$-���abT
c؃�K��CY���m!��s�����	r��U���rO������Z�����Oh���H�}y�z�<��uE�Fd�sc��F�:�饨ef�QzaI��1���ܻUH��F��5�Y?�HjVٽX���87O�œ�V��z�<����,��{�������bdw��3#�x��2�B���v� �V�����N�oy_Oi6�R��H#��i�ӲP$~v�q�w�KK���8ѻ�=K+L���K0�_�����hS�
���;����Wz!ci�N�o������K4ɩn��T����@r�'DD�0(*�[�O�4��R�VM1��!K�Պ�}lĻ��V�"D�zȝ�7�F�\�?&�OE�\L8�8��e�����d��8���z�bY5��� ��/y�X�#��'��eߤNC,����>�0�B5m����&�+�I���\6�s�N&n����i�o��C�"�Q-#����|Dk��"ٞk݊�ɘ���dN�z*PKdf�����Ȯ���kK�7���&(Rf�)����@�'_x�Ń��u����r�+��G�2\�:e��_�h60U�X/�5=���nYg[Tv����F��Ms
�"k� s�j��d���ZM�^EPO���v�l<���ɴz��-��pdM.�ٯg���ܦ��:�ӣ&B���R{��d�j{>R$�\2����|#yuoimEd>�������C������]�������f�JV�L��AJZ\f����e���;/B�Z#�;�Ⱦw�ۊ��ʔ2�cfKh~P�\A�l�2�A'f;6��29%s�歕dE���Dm"*�����c;�Isv�+��:�頛��=8�E�l���Ň�)	��̨G����UsA�m[��`j� n���Z1~���9
/^�WlK��<��W��ea�D�mC|���X ~�z���G2S�����^=#�Y�f$�:t�c�cޥ���P��mg��<@�4c|@�+�eD4좊�P
�ڊ�˶1����$�~,^^Ʉ�%�_�&`k=U`u�ߙb����nj'1�5�k5qW�3����o��Y����g�A ��z�R�q�!���q���LJ���0��qz&�g��}�	�Z0�k�&��y4�J���-�VDO���(��oN������Z�=�XU���v������V��9��~��?`<k���k�� ��L"+wƭ*D*�`�m����*a���&X�l�?��6�ʚ7â��$`��|#s8�@�r|t�21��BA�Mw���ﳐ�1�Z���W��m�� ���գ�5)nM�3�?��yr��������^Ѱ}y�՞�0_*4��+�C���'�I����ݚ���+Ń\9��!p决�:�܎Rs���x��r�{B�I�{s4젬�6.��T¬���|WRx}��82�S�<�^�x��CBۘa�^���_<º:�T�w�*3�;c\$�W��`>���5D�^*��wP���=l�~�<F�%�R�:댧g�1��O�cgF�,��Vs�,�-l_6Ea�;�McC��D��F�a����.��vQq�mS����̙��jpi��m�ϴ���a2��ޥ�$+؆Oz�Zq����7�N_��C}��K8��Y�s�\�=���T�$r�C�:��`ْQ�7a��?F�Vwх��� �\G�� ��E�T��/�}�n�7j�JU���W��ؤ�]k&��o۳��fZ�3��*�%�*�j
@1�ِ�R�<-�����@�X�#��ks
�'��Yș�����s��lp���3���&��M"U��<(&Js�������4���yAݝw��㭈с`Z�H�9�ؙ����~vC,����kΏ���g��/��v�'�̶)�}�Q�֟��g�L���jL�f
�ۥ�2r��t��zξ��2챌/[�KiJ��@id�0O�J�3>H"��S!�i�CHx��Nq3 F��$.��6j�LGn��M�@؃�Ev��!�Ր �~Eu���R��9���n�$��T?���VϏ���j�eW����=�&y�یJ�	�e�+��K� �5�8�������ii&�ٖw4��o<���}Nb���5�t>�l�X k��'�Eu�װ��z����YP��DG'f���G�YC������-/́hŪ�U�1/rA}�qE4Lf�O��{���ߌK�T��t��V���~1�����8i�v�I��ՙ��Zl����X̕�z���x/��r:ӄ����J %��fc�Y��|}\�Zg�]����L�d��r\駵
CV�5cþ�/$`j�P�!����
�C
��UU��)0��*�ǌ/B<ٔh�D�H䗨?�a��c��ذ�Զ$�H{� �s�s���a��ʖh73���2_uЋ��de#=�ΕKzhH�
�D$�y[>���0������	��
W {��%Y���ϑ�/+�P�i\z�9��q�۷�Ak}��`����z�����ş��y*;\o�YL��j<Xv7�y�B��2�$�«n��n6�_U�xQй���x:�W�8HM"Ҕ��k׈��2=�}q��s�w�.����j%��L�D��g�ր/��1�Y��B���L���9�"`�����7��]���;�na�3�V8�{.9�r�<`��C�"�3oN�j\��o����W��2ƅs�����މɊJ2I�E�4o���/?�f����l>z��PՉ��`�0�W4�B��B)p�p�Ǿ��n�ל|2d17p?*��PPAr`?�����_�;��IQ�����Ȳ
������s}7sZ���Qo���*���O�(s���=��o���ܫ��@\�-l,�hn���Z]:���bw*oj���=�H�Z�ʒ��Hv����(��N�[ST�L��"���bQ�W:[.�c�I�%=Xh�X1���[2��$S���� �`B7yf$Y�t���=�Av{;�H^�>�g����<7�����P��:�RB���/��瀞K�o���{y?�n��j8����q�{݄�L�7�@�nh�VU���~�d"�4G}�5��B�!q{в�gw_��s��4��`���)��ڗPJ�'}R�<���R4x�yoݩ��p=~\�5����������Ϻ�+�pR�om �a��*� �~��b8�m�='�!�c�D�E���#_z}�q�������겏�#�]��r���ČH��b;�Wݱ��3h|�	��{�(�kN}<�_���1���W�d�y H ޝ	ٵ�CAچ��&�C��Ħ����e�66m��#�Z�*~��5yGM��؞Xʒ��8��Xu��g�iLH���
<QL��t�GE��3�&��}D&���3�jf��T}��Mo�
,�h|�ݧ�G0���EG��q������)|����f{E��%�wַ�7�4�W���^�L c�եk��Cm��.8	&��Y���Q����S԰��2�~��7�dH�׈����:擢_2!��i�6F�,W��3�����5�rT��&gO�Tl,}����������\�pe���b�a���`��$��
��0���.!��$���+����_�'�)o�uI�SL˃���1�X޴�E�ͧ�SX3劆�!�ҡ������tZo�~blbʑ�F��^��Ȧ��,\�NiHw�N��aF1}�d�j
Z�IY�����Ɣ�)�X�E?��3��9w
��������E�8�F9�2�̫tu��x�+Ēl�<(g;�⍴xF��RX��L<�)yR����>�s����A����x�Urwf�\��G�����J��z�����"i4K"���I�e::f}!t7����-):1óH�U�j�����cI��%)���\�e������bQ>�j3UAf=*	�Ё�7w|��)�c�f��L6�� �f���ݴ�y����q�O��
��-ˍ��Z���@�XL��7�2��\��SZ�*NR��i#�:Zu͖����߅�$!�"�@���S��G��'e�:é�ls�kP�\�����{tE>�t^U3�N��]����lo2;�4VZL���g)�2/�����^M�4r�L�ɋ��TʊP:F1�	r�Yۍ�I�����b�o�0W��D�~׻�cd6�?2�%>���>��
�R��]����F���;��X�(����&{z<d�C�E�_�6�Ĝ^�����	�ys!��HBd�@�rt6�,����0k�x�t��|���>:/���z:�^���PӤ��7�Q��U����=��ߑ����qO�`�&��o�X�Tf���$���K���G�m)*^��f�E���p�0y\j0�o��v��SF� ��/-6�^"�����;�K&J��,0�IQ5B�ϻ'*�$�M�7_����&2��u���yIKZ9�]/���I�q~S�;E뫥Nsu�����T�M;�2Az#��}��2e�ۯ>J	����Fr��<��G�ø�T]�sa����YL��}����-�[�+�Jؓ��"s���j/-uN@��4���sA}�Z��#��3��0��_�ߐ-~��E�����G��7p@��:�������Y�4��L��`��q�PԽ�W��<��i �y?E�ե$ ��|�L:��vn�3��yv��}^�>��Yj�ͧ�>ثX>�g�z~��<e�oʿʒq�&u������|8/7���d��t!v��0���
�� �U�^gB��
f��$7���ٝ��>��P�7�uIW�'�z_�x������	���з�[�}����F���m��Ή�&��¿H�@�3�z����#�s/r�t� �U��������n���}\���x�=�D�t;)�]O9�Aa��Lׂ!����T�G��
��C�ɗ�y����В'R�ꮨ�Y,���*�@��.�"����a�$��ڎ�Q��+�_�l&�F�A1��[�wmW.>���a����3S��%���g��>���OJA�L�cp;wq�J��^�����Tw_��;Pct�����6�(9��_C?=��:�4t,�VK�q��T�����n�i�H��з���.�E5�p����r�`�	�K�Ey$0g2@:���r�� {=c���M*���bw9�?z�8���T\��	kW���=AG�C��7����g�����Х�T���N�a�{O��3��:�qX�]*���˾�=���{�"`�g����^�˹~����p�r��}��ݓ��W�??���<TdP��N�qh���FEӳ�[5u� .�<ꅽ�s�[���k������a(>+�t����j��r˫����k��'6׼��oB�.y�Xf���<U`�� �PY�� 7�Zb�Biu����[~�W�|�o.-0�-Ƀg4_�6o/��lh	��~�K�LJ�[�7��R1~���#�>?O�lmwC�Qɤ�*���~(�EoHJ�o�M��x��'�&Qg�q!�6SK��s}���71@�T��b/u[�)�C�j)2*������;��E6D�1����UX�8fa�����T���g�w$c̗)]�Շ(��mSUE��9���K��_:��0Owk��o f$��(��W]�D[�_�8p_�镓�'�����3,Z��$�iǇ
k�Υ4|��3|9�ji�����	�a��!^��6��I�:�XeIb����0��"l�VK���c�J�C��=�./%��S�]��Mt���C���Qn���	zc!�O����|!
o��YRo�H��]�Lt�$��=7^M:^Vq��<�l������{Pki��r�A�۹dD)�[N>š�qR]�Z}������8�d%�Č:®�3@+���J�{�	��\~UԂA\Գ-��R4l:���s7�\�$���Lk�&�9�8&�uE���wH��5<�!�QV�ʬphMl�Y���5���f��L钓�ɛ!fI�-�9� ���a��1C9������<JrI%�L�ïw��(��2㼯�^��[rߎs��x���͞1����N3����~�|C�#��w�A0�.+��6�.E�,f�~����Hԉ�s~!�`��O�l(΀����* �W�C҉�sx�_�f��o���KW��O��&�ui�P����a��$84���<S���r�N	��B5��S�0d>�.�Mg���}�9���jB�XT1l	�/��ч͌E�	g��{W�g���� }ϸ�&�{zA��Nq(v�~�xu��r^��j}�{ڹ�D��%T�+��t��"��Ȥd���`�[X]HAr^Zg�H�r9r��{h5\4ev�~1�~2��	SA�Ϗ�д�>��|�bQйٍ�g�~7�q+��O����uC����hGG��@�;<�4_���ne�g�H���q��cB�&�n��H��d�u'[G�J���u��&|L����p@$+]�d0���$ʲꤙ��Z?����
�b�xxl�?�`_kYڷAqYB��*F���j ^y-L	�?�˹��!Jt��"[<G\ȯ�ٛ'@*�Sv�#Z��E^&��p�$ؒ %v��j� a�;9<��?�Jл�:����e;ԾJ4O�r.p��[a��5�݂���_;�n���s����%h-�p�3u �b�yRݙ��Ѿ/��3j���.�<�����jT���|�H�XA�сbkd�J��W��\�m-��}6��g�v9o'�M���[2b����K�-9�ӡ:i�D�� ��fL}.�+���]�g����u���axs#rF��
�$|�Ou�5ţ��4YUfk�L�
Af:h�PQ��yVTN!�K���MY@�!��u=�~����ζaD�J�ME����F@��3���MQ��c�8s|F����W��9�17bHK�a�FP[\u�J�Gl�"�:�6<69B��^5 '��tw�5���A*��@�ckX�$�̆��Z\��=J$w�kD9�0�.�$��ā�~׬x�~����I;� dp��I�p�{�f�\j�H0N&J��e����,0YH6D�Vz�$]k=��py���k��!hu���[$z��ᣍ�����+Q��m�F4I�I�*p�l���(�����=��5�R��䳣5�E����p�O[fÐ]qF8;������<w|E`B��Z�Pw�j.�����0QX��h|E<"�Aв��KA����p��PX{dp�
<yc��Wm�"��/�������{������RfyN�ɤ�	��`�D��fQ�ɛ����U�5Ĥ���k78PӗT~��� ��ƽ)ܺ��.�[3w؆$���R�m���Y	�hE�Tѿ�� ��ߎ�K�o�����k����הڞ�-��LK���yn�`�3b|�ֻ�	������.�e��c�f��<!�W<a�:UFP�Qi������2��(���o��͇]�|.8��V�.���V���o�7�|��gT: ,�,���3�d.R;���a�)����q��7��8X�%�M'�HP��@.�_�J ��+��_b7�g�庢��E��E�%_p�'�����T[�ϡ�Vŏ�!�L������Uu|f��eV�����r�퐅�&S�����]*����p��*_�8D9�:��LAk��K<DgYR�7R�=�uw���I�Q�4�2g�t��D���e��/�.	W�%����LmJl�{^���x�0g���^�]=��豟M_I�I? �V�>���<���K>(�̿ˊr��+��PSe�+�̧�~�&��!��®��e�@���xӁ��1 �Hqf������!T�#*��6��1���??��__Q�6��6έ�-��o(ɽy4��[����D�t�&��*��V� ��+���Q���<��j��<*�q�ztv��h� o�o�j�sP+K�>�iN�E��D������Q����kZ�*�3ݒ���G�ȅ�pl�1�ct��p��������ށ|��P�����u�Vf�UXȔ�^yjb\Z8v��_v���vBA�MƆ��/o|���Y$Y
�#������D���]�«d��ܰg4���B&,�q��ߜ���������(ȹ�zpV�4��V�H�29,="�|㐐B�C��x��>����O�ce� �R�y9Mch�B^��*L�Y��)��̼djMۃ�O�X��Rw�Hy�}�Mk���C:�h�I{}�3ZX���8��i�ȼj>?�����j�Q�#���F�쀹� G��GP`���u�-�{Ni]�ټ��Z��3����5J6�����VN��jߑQ<|��ஃ%ސ�)�5CX@Z�!�OK�,�@��϶�c�B�Ga �4qS�-M��8lUʭ��ܿ]�A�n��]U�;^�ug�3����?�=+ۖ��Xi����o��EB���#�2�����ů4�;:짍��V��̍�˕���� ���r��>��ri�	UoR��-Ƥ9���n�q���;>�d��>ABԩC���+�L��h00vEa�����Q��Bd��Z�����,��"��j�$�BH�	��`��o���&���q74�}��lN�l-�ӈ)k���9���g �Ƌ�ю��Å�x�0<:���T|ͥ�\�:�Ƴ%1�<���40�i�6r�<��������xK9��qX�&kJk����ڞB;ք��7:{�<�h�zV-���0a�R_B��9/q~$m��!F֥�w��\Lc���u�/��.��@�H@�t1��Y����sK���.�߹�0~,b~�|��2g�[-�Ba� 1�ݕ��πL�%�:b�k��/�Pف���
CPD����y�=��0c��ɕ48BZ j���sN�_J[�0����^�Y"�-)n�s�FlHk���";u\�	k�艍S7\ƛ��$����o�Y:������#�lדM���;��E�Հ��q�FA�LT8�Z�4�^�b��&J5� 5�uڊ,�D�!��p�����FM�Sk$~ʵ�sD6�˗�OS��ew�F����A�+����h��Ky����$���P�C��nw�N���9�K��W��ϡ�Ԅ�tt��G��n�K���B��E$�;@r̶�����{��m�C�M���x^v�SR0�gm�s�$!'���[%z�d�t\Uߠ�l#�dV��k���P�,�P8<�9�i���r�����@n���')o��d�@n�r(bDJ��n����s����
��.XiG�z��ɹ��A���4�_a^���S̷b<�w�N���|�l�)h�W~�E�Z��v="ޥ�U=å��%�@��R��;��Z��y�e@͛h�	��,��î�{>,�|��=CX��[p1�<�/���͏RP���~�J�1s�%�M��jMN ��O�7���6�&��%�ˤ]p�6�-���x
j^K���gwa�,��Y^H�s�V��!�A�ŴN�RN"�m��V�d�9�[��I
�LP ̄?s�>ˈ�~wǅ;�	�$�Lyn	���0�Ts�̯�o��Q�Iz�ga36I+�"=G���v��LO�WB ,{�sG�0W�|Ʉ�!����V;؂����V��R�I�1����h�Qx��,�:>;|���6Ee�~��:yT�����;x�C_�@K�8�ho�����B��D�2���� fX��;��1 ����(��/|n<t̚��}5�PJ}���X���-�]Na��:8 lw��!c�s��P�#T��U�������/�@{�􇸍)�8�ޮaiS��t��bo	K�-�׹��]p��u�;�Ha��UV�Y�g�a��.�Oސ_����%��iR��fvN^����?��J��V�������M��I���I�������w�C+b��H<M�V��֒�\���q��3�Oo�/czե��9|ܛ�Nz?�q���ʤ�^7�|<y��D��T�@1�{�X���-�����J��/`v���sH@� �?mD2�u���H板mR��Ռ˻�����V>��ZԳ���e�:�Ɏ7Pi%;�3:�5�9���pb��C�����I�k��2*X����� h��sɐ������TQX;���������)l4��c���2���cd����+*�{p�,�U�M��	�[q�U��<��[
��ɓ"����p�]P�3�����Jl#8��_۬��4��E=�(����40�@�`�^��rx��fQT-
|�'�m�t(ۏ)RXE]=t�CC�E��R;�Q�&l��fC��q�z�$/UG��Y���_�N�(MX�|&�$F�^%���Lg��|�'B�.��5h�7,k���ҟ[�ENxt�I|�7F�D9����;=!^�|7P�iE�&yT߈i����9����"
��5{�6��)&�;����t��m.���_�t�z����L��R��>{GQd��F�\�y�O_S9�ۛĊ_�b�͐��t��$�
�7�&.�$%��>��sيIUA�s݇'�I���#����@b?���?ċRDΖ@��WG����2*����Su�T�%����_��I��%ScJ#p�i�;��}�z/���mSG�x�פ���$7@��ms6��\N��w �}��U*g�T�6�u�Z���V�۬h��=�p�92_6���R��(�����?�A�^��Z��2gD��
9覹�d�U�`:���|Gd�ع�\����2iu��h�쓫5ͤ��l�59��:g�B� �S�%���Eض�cb48�`#�ʯ�e6X�Wb-f��ʇ�AHKDƧ}ř�S�. CxJ�[�
�k��"�0'I]�����81"�؂�4j�ifi�뫆zJ\�W?���>�dt��U�B���˜�O눥9���)�}Qq�Bv>nz�JN*-�F��$�[R1!p���b�ʑ閜!.�{�K���ּ���Չ�>�~d��%S�&���-�|1�<�~Ì�Ͼ�.��_~4t7�v��DC��� &~���a'��i=����)��A�诎3T����-�麯h��)\-讠���W�\�$��W�U�{�+��d@-Wܳ=��^�F��@@P#�9 �S#\�7��԰ѽ�=��2��MV��WԻ @��_x"PA��E:�Zsp��޷b�_s�ꏚF �R�Y���db��f̉����*�	^ v��wo;mx�Y2he�ث%�9N	{���ͧ�!�#��Si�K���d�P�,yat��ٰ����x�\�Gc_��\U�x��j�o��� �U��s3j��rCJ�3�p>>�5����[��ˮɵ��4��`a���uf�O��=�a��%=�ӗ�6@��� e��fc�D��C��(M�/dxQ`1�'
�lJVq(��Ht�.��$0����!k:���09��@ԁk��ȫR#�3=q^�RGt=��bsm��>-������R:&�۵��s$(��&�m�'@��b�5y0u������sW��S�4=k�.lx��ַr����.@�g;���	��+��+��@�EB/�Eb�X�^p0��e:[���𘒘���g؜*�a��$&W������9�hَ)
wU��֗It�"\әxzL�?���]Zޓ�i�=�Q���6#}n
v���?�ɋؘ���)m�|g��fݿ_���@B����E4F7	C��X�A��t����|�	�*i��J�>�����)����ԇ��6���̼7��b����V��с
(��2��-6Mg��y䬓���;���t�XK��G7�yÀޙ�+� mp2#Zܜ����;��f)&;�=\�����g�;�_r�+1\�j�p�D�'�4Z�g�}Ғ�*�)))������-n�|�"+�g��>Z䔍��t&f(2j6�l��J�~C���+Lk��JrF�B������m���(�(KnZQS2�a�۽���W���m'���5L��Ȭ��V��E���5�?��E����"�ÿ!�� /�u������c�\�?�`�ݟϻ�b�Cy�� �J�9^�ȥ�|��,gQ���/%�sM�5-���#�<�)�ERiX*�+�.O���CX61bXif�`����X�%��z0�wQ��B+ܓik���ņ^��b*��U�O( BE{���ݓ��Ho&C8�r���?O�2���D� �1<۹}�F��)�U����R�{K8G�;E��S����Vt�6�B��Z�]k��}2Z /ڗ�<��O��M�,^�5�d�6S�ba���&Z�6�nt����W�F�U�1y�|y����������ws	aMOt�����c%+[����WWV��W���fe���40iE�1$�}����`��K��s��s��ɵ��m�} /�h%_6ۖ�I0�)��ǐ�&Ӏ���̋r�'V�j�x@uX�BKE2�k��ߗ_\��3�u�y��䯡 ��z�z��S����5W�a��h�.�D�'ˋ����j�;5����Qd�$L��'�����S�p!�6�:��<�1}��,����R"������l�b��>���S����y���m��������F�Z-<uE�f�?�H�<'�qL��!�_u�ﵿ(S�4��.#f���6C_�_�m��b����(�C�^��W�,NY�1�PZ�Ӻ�q+�`_�nE�	�)���=d�(1�!^�@.�y�C;�0)ݭ�0��!��7�sy*�<y~���A|1���I���D�&b~i�*Oʛ�)e�Dk�H-$k��M9��`�AG
\����fk���Q_ߜ	2�n!b%�lt^��)�6�Z��~1��Aqa}BSt�KޱeU���CI]�lD��v漮��91���vNm��*c�mD�F�*Y�+#*1B�|s���v4l���F���&{�����"�S�n�Ī���R�V;��3��:��;,ɗ�;��0(?�7�����\pݫ�����a:��D���_������.���2�	p�&��X���~L��s�W�&�.�r�ʍ�S5�i�B���:��N~�7D�_I����_����\n8�+���R{I/!S�����$>&��0�t�����R�,�X0$층u���=E�n��|���/��"L>\j��P���At<ό@d�B�6EU<B�^I��|H�R(�6Hy{�����K+�����"�lD<4Er��J��R��R5u"�A�1@o-������Q9��xm�L��Aa`/���Hh��
��e ܟ���<���[k?2O�k��*���K[K`R��-r�L�M�� E:l�?�v��2Y���;�r|}4nl�x� ��y�.���V+3o?�s��}"G��f��hS�/8���26��](��Fśق�#tCe�j���E�g��_W���{�m2��G��O���%��,PY���ť��ie��Z!c(��;@���+���׽�A�� "��'��ɀd���S��hZV|��K"B5T�)A���{���Cv���*��K�5D@����ٸ������������ʇ��4�t��n4���pc>� m���%8wdH�R���/ǭ�-^�'�Ys���ֳ-�lC��z�]��{L3=���mDQ�$���]��k�o%�
]^�G�����1�c1s1J�i�M,��K���;6IPG��A0��%R���
�=\��5TN����|��!��9@�����ex{�|п5d5�1��&�O�I~h��y�[薶�y ˃�	�yY��|�e�I��п����`�Gv�$ʼ9`ѽ�ԃlv��ԍV�y����eȏjK����	M�X�uF���E.���Ӏ����]��pOU��SYҝ�Y�!��+�����n��>��-_pH2��ٞtE��L1�o��D���>"�7�G��^� �K�~���;S���L�C�����-����\=�{��O�Z{V����|}�b����#�^e��������W�gAy�^E�"������?�u�7�P�; ��3����X�:�B�p��x��c�3c:��:���>�m�d��83f�������p8%�{_E������/�nB��B.��@�3Y�&����������pD�)u������ ���}��;���� M@�9�����GxM�˝g�9�u�T�D9��o?��x�LN��\�;��"�Z�W�q�H�t��䌃SS僋.�~���+�����?X}tzv3}�w�s���J����*��Ft���1+2�gXP5- �y �O�6'v~c 7��n3�1�\l�`�o��b�Y5�b���B���d��eHa kƛ,籗$[}T��9�^�Soi�0o��`�OzM���#�d���a�E�X�����X}��}�2�i�Y2;C�'׎{���8[�«����]r��#�mX��n2w����`��ƜO��#�Y�����ٗ�-�!�:����j!������L�Q�1j*%���۳�cE��ec�xJmY���-&�s���~� ��m0Q-r��OvW���P^f���h��ҎLʛ�5�>Ƌ�[<�e�QEyܿ�Ig4k�c2Z [R\0�?L�B������u�?pk�6�_�j��ng��yR��2�]�<Ȓ�R��J4�Ć3��39+!��R����O{u	��(z9�6���Q�4��KȢ��z��&r�=o�6L<~%���ڂ��4�m�\�6�=2l@b���F�ۺ>��m�TOD�r={��ٷ�2� 	��/f����{s�&�b���ʌ@�����K�l2	����)�`��D�<|���Ͱ�JV�Zi\�"��q��q�^ {�>RY�߄���{!%`<{X�5�����,.뼚!�8�}(��~����g���ݤ��� Eݏ�N�J�[�&��9_lޤ�x��:0�^�ߌX	�/v �!!��h!-1]w�1����8�Dg��^�?'��:�C'�4ն?�=��S��J�K�FCG�f��2[�?h6kPT�D9�:��x��ο*b���(6jwK�g^U?�Ta�#îhy����[��?Q� �k� �k��x�>�r�L�x�Y�UɇJ#8��� ����Z/��Ԥ/�[:��O�|#)C���mO�p|�T)vK�u�2��+�wrC�L���FL���uu���h�F�Z�D���I�!G�0�y�x̤w��>&4W��g�^;�*�]!�X��`
���/̃��0�|�|�mw�Ƹ�� �>��ۘ��E�m\8�ZZ��"�1g�=�RA_�RH!0���G��f
��D�	�H�Q���6�R�Ƅ?2��'+�����?��p���!�p�I5�ȕB���ץ�,������պ�j��Ӊ[�ͧ��vU.0$;.��q2��R��wy^h�M2_a�TԾn����1ue1�L6o3p�,p7���z�^ӏ��	dM��#��>��n�P�� i�q|Źh�f]!{�}���hEs�����ľUKڞ������B>���P��e�����8?A���%�^�qF���%�0B����4��R�o3;@>DC��o<|Q�FJ����R�}Y�zSb=l��T^�I©rI�LV5�0W�i˙#�-��Zr�L�����RlF��>
�9�6��Z�"e{�ז�m���p%ɪ/rn�i��f޹�SNϐV�ᘙ���eD)��ڼ�>�<\��!�K$������8��i�"[�ȕ|�6ɮ�������ImN(���oϊ|��O���˝��>�E��s����RU\��Z��A�fo�S�B�e��xŎtS�����5�_�?��^�	�ye5ֱ2��U�y�'���kv�a���u�x��3�(��K}�|q���i��?�F2 J�d��Xg��z�l:�ֹ�q3���v�$�+p��~�	�p���/ޛU��'��u�Ŵ���q�/�EU����5���&�`��s*DUn��]�AKn|�i�iyL�ք~���c��<���h/��}�{#�]@"R�B�Y9��鐋��@G>�?h�`?�*/�U������Eҙ��.�����5�����נ���S�#�U���x'q�g?�Ԓ�u{��2�k5��f�g�_P��x�̍g�O��Bn0ϖ Ӳ����7$��҉��L�!�X�Dq�M�9�#����9��d��%��ܞ��t*�rF����	P��yXk�d�/�����r���LMHƟL<�e(��� �;����b��"��櫕䨶��M�{�����<�N��-�h%-kc���(VOh���9���LJ6�{.��.RT��~Q��V�!�����ǉ\:��}Ts���PKH�����g箮'�s1�X�g��߮�S0���)T1t5���!!zҎ�$r�Z?������]��v��s%!�&T���5����(!���t�����J�7\y��ʈbJ�	b*��3�C*�V����pdc��C��0�v#v�滜s8-H���=�������?D
�=ȿ��-QgBh�0�t�ْR���� �[���y���X"�0#��8@M'`�?G5׫R����n@���ip~�87_ ����0�|�{Kޛ�����ș-t�J�H�l���N�M���HJ g�w{}VO8���]3dF�gs5���Tn���xRC	W���H�޼��1��1ɯ�}2��3ZC߈'32o�,����s%1�a
�V����n��0�4Mқ :�`�_�D�N}ū�+s���,C�*�1�ez��M���YgN g�  �Lk�7WW��=��x=��MZ��i@�xY8��Z���R�tr�bi&�XQ0C �2�K��.�m��X�q�z�'(�_�Ck�ʹoa)"L�x
�_�T� l�ZnV}e�8t_���×j�}��|&<zFʿ�B�*`f�d/�9a�!(�{��+���S��c��S"��-�#LL��;��DmxGB� �j$��`P��
�%�8x�C���/�I��~���񿊲�}:�K�h�0:+���Y��Il��_�\7k��iJ<8��e��փ`��;g{����9�� K�����E귝X��Zj-{�`)OCs������l�n�� �9�Q��Cd��w���^�C~cy+��<�>9Ŋݾ<˄�f���Ƭ�?��ւ������	p���E"�+���R�^H��o{�4������N�����eR�T�;QpG�A�>��̡�H�:7)j�w���i��Z�z��/�UE�s��Ȅ�f����}D�r���F����VG̮�Sv�p �;Ki��D�&�x:j8�|Z��|�&���S7W-�d�W��јߡRy(�H�_.�����M>�h�^�3yߌu-XF���?�c��E��D`牽���Ap��N�V���(p�����R:�!����y|�(W�o�{-0D�)���|�n�&@yqj���E�6<yL~��!�n*5�F�T��&(nI�0�,$����~�96�@߮ w�;v�M�Jd�n�7+Ur��ؽ	pd�ݝc#�@���R�����TS-=���?�� Ȕ�c��6���+.�ܱ��N8��D�f�q��4���CGB��o���HR01��I�/�s��f	���p�������g�n�������u����M�C�� ��h~uqG#ad7�u���MwOJ-c5�N�l���k/d��`����<�p���G��{��ϕ>���S�������8�i����z	1qQ~Da��~a�P{��1�������73�1O�f+1G�X�S:q�@yH�s����
�� ���6׈e���W�v,#���x�V�;�Ժ���.�=�]�IO��f��CV�Bӱwvil�"dVE�d|��TM��3�H,gn�[Xw7���~@n6W��&j�X��Q�;:�o:>�DQ�Xm�{�C�4���q
:�C�i9vDW|z�pes�EvϞ=��w�铋�R�ur>�.F�^<?CH�#ָ�9YG�d<3�%{���Eڐv�������'n���KjˑVj�*�;��82r���� �߅���$E��\e�wr �����f@0�=���0�Y�q�0�.�L]S��Fm��xP���z�:��6���Z���Y���)�֗V�c����<��mPd1�o/�+�7җ�َϑ��ըA��?��"���w���$m9�U�N�.��8��yf���]��/,5�`�Yؕ$V��t���08c��t�Z���B�� m=�e�/� ��P ��A��/��#:]@��4�.A�@�
-]�>iUj���Mn�B�/$��E�Wv��Lz�J����z���rOL���ժ�+]��ȸ_��C3Of�9��y�$�o���-K���xo��w!�������!�����h�N��p)��]~`_���c�*�S� 7'��>O�e� ����TK9.��t�c� #x���ТF��eC�T闏zƛ,Ov�7��j��[0�,�BxC�ݑ|�u0�*w�0u��\��D+䴚��J7�. q���^Tᖝ�y��l
��_�7���Į��c�7�P�(���s��<�V/$����r�n��.�@*�O��R,��������*�3e;~ :�1����3�|3 ��F��i!������������-h[������Bg�%Rw�ݱk��q~�S��颸�{P7rl���ȑ��υ]��<�uBDs�v���d{_
�q��l�ަˀ�D�3����<�����=�P�Ǌ���7BQ>(G0t���@|Et��4(�ʾ�	��W&�у� �\E���>p���ڂ�'!5�ֵʁ�Xh9�Y�/�k��0r�3Tv$�ɵ��:��D�@��h\��L�_�s8yГ����Y��r*L��[�>ĜF^%��{�X�m�=�Iay2W�N��WW������<�a� b��ݠ�߼vT���v��SG��E<�N�\�$�=����Ƚ<����ƄxpUm
�0���t����.J*�$A��s_�X�Z����R=�n.�أZ���!�>��3�.K(QԿ�h:'����-�z�S}�3�<Z~�����<�\H�����>�{:���^��0J6|����rA��Uäd�3���\*�`z����O�|
6\�qQ�4H��w�
���{�2�P� ��Iԃ�(û�\�	�c���ZfcJA
s�s��{R 2�N�Un��Mv��û�R���Dd͛S&
�HDfsy���lS���=��),=���/�n6��fV�W*�ꚾR4��Ҧ{��,�W��_!��Q�zY˺��]
�7�G~�	��"���E�;��,��h,�qn�A̟`N�l���ɹt����v���X�!�3B0ɈO?��O̻�s�&Ӊ<��IP^��]����舰0_�l��?�fѫ���*��һ6����L]�4��J��j2tV�t5ы��FD=~�l5t/���U�Iօ�v���2��s���-�L��eܭ����#�d2ڢv^~����UO�6Ͱ�3ڽ٧��P]�I	W�9A3o�H���-Й!�yGoT�(�������C�Z��i�e�#��Wcy�!h���/J������J'x�!����gs:t'��I�sc^��|c��ٳ:~Y�yɹ�@�c�Xp�@�>�r;<�D��Q΋��.� ���j+�������$�Q9�����t����օ��@�b������*��ʨ�(�	������>�ڑ�� �?���<]H˫���%��$x˶��'��hC��LQ�p$�])�t���S�zH��2�D�W�Xn����4�˭�6Be��#w#r\�;f�"�N�$ʲL�v�����t�%z� ������2w;�X�]�g)7!d ��t��R��%�=�'��b"q�[D�Y_�|.d �����u���uR7MxE�Z��2�$����D�7O`��3���R�me�O�}������p-8DI��ވ/BI8�g�g[e���"7��f7�K9֛jX�h��V�yЎ��`��kv������;3S8�~���dհև����"��ߚ��"�2d��!�v�X	K/u�/i��W��exc��D���%&�"PL%>eg��&]��i?�:�5��8Dw`�3d"��f���yD@��F@$
�Q��U���G7�E/�p� �!����br�{��V�$�"P�y-7STӬ�=+DhU!�O��Na��3vO�7���bF�D��A�$�q*؛O���|������?��adT���!��y�S�d�u�`�}W�������ȅ<h'k�SZlS<�#���є���7ѽ|C���<����3� �d!ݪ¸���ځj��h57񦆅���p�NH݌����J]�8��+K�S�0�����~'~8w!�n�@�Y�dѯ!���&������ZA��0�ţ�;�M}�N��OV�Ъ���j���uZ�| ����UmO��eXLو_�-NZ�4g4v�B���p� U�c�S;�8�lkB,��pU"�'b��$�IM�b�PGu˾yO�����!h)�`�I�js�5��*���,�s��Hr�	qM�?��aW��%=�}[Q�� �λ��W.��_�	�=�7���?������9�?�49*�A�)��S�/W�Y5F�����Qǋ�\f�Q�BuhHhi�BsI�:��8�1D�0p�"z�0��7��X���Tb���}��{^�s��hq�~`�p���W��ym� OD%�k��2�����.��YD��C��q�.48����[�5�� ��d})VgU�cx����N�~�[S�m9P5�L���n�2e+����&ʈ��(����ͳnq��#�q���!���K�(6
NJH�M�:�%eu%��8��ݜ�r`�CX�����E�����(�a�᧢FSơ�'��
icf.M��=��bЎ�r��ѵ����g�\�H�L��������IY�F�k�����>җ<�C�P��Y8������) ��m/���ްW~�BNS��YU�!�5�YI���G��&� G(�R�8�8;p��E���+�ú`_���mx���G�b�g�@؆ z�a�l��FVz�	|�o81Sd�x
�ى`^�l@i`��!c)#Ɔ��!�c�q��HE��M�ۉyE^�2�=_�+�U�ܧ���ߤ�|f3��]d�A��W_C�nd͊���-bG�39�,1[�@�K��u#�;�EjIH0�٣�"�w�\��R�G\&Ι��/X�i�ֻaz�$�#M�y��������� E8����O6I��8_�}�tlC��a�<�;�Nݷ��j����.��ʄ|粻�?�D@s*�0��n��͟\T��͏���
�17�L'Wͭᖪ������*,>��eUy�� ,"�%[�TB�ﾍ�e��#?������{�_�+����ʢ�=�Hz�rI<,D�&���8/�#J��±��>;�JL�A��OX܏a�����q��HX�Do"�ΰ��	Kþ�O��򗠊� (��	�^�7��G��^�N/IHk<�nO�X+�� ������6�!�<���O]�!S=��eN�$�J�r�m�ߘz
��Ə�Q�y���3,��V�n����=��QEg�C���J�;��m�D���]��L)�<��g�-��&��7Kw\¸?�oq�4�gP���(32*��y��layN�B1�b��ș��c�[���9�+�
F�؏Ġi?:��Q�>l��^k/��@�Y�Սk`g^?�v���T���[r U^���ݘ4���c#��,�����x�cP��نJj��/��
������&��
�����6�r��
�~\�9F�n�k3�vr&�ƿ�&���D/V���I�i��������o:,��ύD��{C�i�J�?���CHI��o��L/3�����֏(�2(�_�/�s�8C��.~�R��lN��K^�
�_�l��^Ƽ�I�˛�[LY�I�Q���E`D+�v�������xzi�iՏ���Z��KI2uH�$���(��b���K�E�
�w 	�?G2-W�O����V��ڳO�#�g|�8m���=y�?X����}��~n����*2Q�i6_p9�p��	f/�ׇ�����3� /]3a�j|�aq��F��&�-�C�!�����mpA�j��6����Ȃ����~1i�o
��yF�68\O��	�l�J��FQ-�7D{�2���>�/�C8,J����zH4���d���͢9�/�J�����x+�뉗a����b92/�>=I�qoٔ:�I�����^ .�Y�]zγjS�N�q	+_PR<5��k<��Rn�:�t���2�Htb<%�F��W?�L0��A�+X�3%&�����|�;�Tk	z[I�Fu�D�Y��2�q*�2@�'���0n��5���Iִ�����ٞ2�CdеT��r�8�.��;�Nh��2'�����q��4bYU��׌���Z�X��D�*�H�W�T~�:iH]!2$�l�eP��zH���i�d��'9Wkm�/:Aq!��m$>��65qU�x�:��ǝ�Rb��@'���z�Z&	?�.�tc}�"ۥ�o��%�74d[���y��4M;K���{�/'�4�F�N��B���&5�ý���{�'�ܖ�dsةC�j�`����G��@u(���Jm��6H�'lz��R�w��8���z��*UqH}l�g�(_��b<�=�tq���s&:��$פV̥�:ĩ�RTC��S��r%� �4n�Ł�Z(���s�<��]E����ܙ��X�����5��K��YC j���X�x{#Db����Z�&����h��x*�T.ЗN�2��Ĥ�;�2҂y��}� �Nv�%w��a��]�\��-,~�u?$�鬺]�$��oa�c �E��KA�"��NR�L��41}�(p��pKRټ�n\�R}£�9��'���yY�[l����'*��t��X�ڡ�~D���rm���*�I�yP�=�?8ӆ�.��i:�cX�3���쩡D��+��$11�f�m��!�n
ʕ��k���
�w�~�=��Fnj�����".����+ȏd��h#f��N�e��X�������s�h��W�#�2�d�;���Q:
����G��LiN�
Ī���~3�.��ԺN��5~n(��Ł*�1o�`'2Rw��\��x�gl�Gy�m�]�������Sܛ�b���2>L���^�w��ZR�)g7%���#LA�|G=l+ޗ�+iԳ���=S��w�#���\������ @�)�5�B�iGL��,���5հ�#����*��|���&��7�zT�����6���+�}��T���s�>�m�D�_�UQ5��w&�%1������' %����0���qߓ�L����$�D���K�QW@~@s�qSS���@2E�
�cx� ��]v4�c ��
(\��e��Q���`��'��ox)�J�� B��$72����FfZ�{;�#�?}�j�(���&��;�1���6v���P� �`�.���F�j��T}5�L!��lӀ�u{��`�B<B�BdO�0؝��¬�X�F�@�XZ^�PF�g�io-�K�L?��v�3������a�t��7I�Q�{rw��n�k5��R������Zu�*l�7�zE1���`X\z����X�Ҩ��C���O����tіR!��l33�v�#��(��������PI��!34�ZXt'F/��fW�o����.�YGf��Y�1��x��ΐ+���b��טM
���̇>��3��D�G+�v�!W� /�#Ӎ�	�Y��	J6�Jߨu�&1B2fx�<����9R�>xH�udp���N�"��I�����~j������ь�=�`}�}v��M�`��A���'X��S8,Q��.0��*�o{��e$soW_��"��X����Q߬�$�y�L�X�� �Y��l����}���p�c}�����ϋ�yi����B�1����˼%T�|�t��8S/�7 ���*�Ŵ-��ˑ�W��Dr4~�kQt���k���=�t׉8����|Q���`dZ�'H#%��+�g^�2��RDR~�︭(Rn�l!^��	���	�vOn��m���H�n��G��0�zl�=ւ'^k$�[۷��v)��t�ּ���|;�UO���4��_T6  4���_����K?)TB����Q��{�@形� ڗf�&b� ��{���UoL�5�6��\w>���J�o�]��n}��G�H�Y"��*�)�)*�4�fkY~�c!���e3Z�փU@�M�B��p��`�?�2$�NZ�K
�I�l�"Gz�?�B�dT1����<1��s'6A[�\��6	�q^��$Zp�U�lK�Tf�;C�KDA���0�[���96f*w��LP�����ȷ�P�e�Ƥ<2�٤���c���/+���gA|�n�M� )h�2?D^+���Ǳ�[���툏����0�[�t�sq���.���:8� ,�BZ|���E��h�_	�6���N�؏8ae9�F�'�!V�����]�k�%ٟ��G{k���*��^��k���=;FS�I��\`��r�i�&��u��q�)��R���Y�Z�a��;j$xQn<mK��'�z�d"R�+J(��o�L՞���q!|w!W�A^�M�+G���
��V�\pwDhY�n���������`��
�KBT$JQ X+@��8:b��2+:���^�4w�J^u���*o�fZ�����a���7'�*G���`<����m��]�=dz��;���dMhJ2�/�6-�,��F/P[97��pf퀜�䱬��y��92U���~��V���oS�wX� z�·C�T��#m5�P��aE�1*��I���-U��m�a�Υ���gz�	<+YX>�!�ݙ�v�&��db�\R�Tܲ����8�"�##��:�NŶ@�/r��0n1��yt]�q!0��&���O�'��uc�R��E#��x&Y�=��߯��o��d�:eh" 1�\�*�-X䍅G��Xw��ͣX�LY���ȅ�L�Z ��M;.M�G���D��x�`_��Gw�������rA�db�7}<��\��4jh�������p�C���;z�L�
�E/�	��mX�;���ĻsI-�u�s ����*�"����r��!�r� U+��Ս����8�gk�.���a{qV�
��:�V�A��?��Ê����|R�L'L91lP����8x��+�ӁmF�i�'h�B2ڌ����X�X�%�QA�����G�V�eo�R�y�ј�֖?t!U���5�p�Z��PI�k5v
��	2��,�~7mZ|%P���
�����-�0E�b�)�T"e@�g��ˉ�aFwmC�J�R2���FO����K�����{�����m>�w�4ۿ���h����U���P^~2�U����(�YY��-uv���a�c��è}�g�AR�4{����G���T8�qb�4D�"k��8��ϧ�3W^���<��RJ����8�!k��%�C()���e� F�O�p&l�b[��%f6�
����z��U\��:D\�����L�{ۂ2M�����;����t��^dud�F2���Q��Ao���0𬬫���F6����+a��V+������ցYK�u!nQ�:���G���)��L�G�#���yK�-ti)+j����|�qD1`���hb�,<���u̧�Y�h<�D9��y��1Z��,�T�5��3���S�n�����v�5I"����8�ݤm�s�gx̌YKtL{�椓�ne]�Ǫظp����Sm����I�5�?&PT���!�ڿi�u��g�lY/��9~����'�=}ճ�Q�Ҁ��{2��wZq�ul�����ۼ�
�if�a�	�P��7�_��I�}*?1kGi=*�~'5��Z������N�Rb��"Ӌ��g��Mx�8�+�K�����}��LY;�A��� £y���[�[�;:.���R*l
?��9��rK'����xH�D�'7�>�u@C �0���fC#)´�J��� &o�t�����-b@���>&u�0���b�JP�r��9�e��a�D����s���u���X4vA�M�(�x�BQ�XO�N�J�&@�ÕO���C;��ѬÀ �BN�w�
�b���鱂�^d��-��[j��eS���*��T��XV�'��=�y?YL�-̢t�ᥛW)����s��$��a�ъ����eX�+I�A�Bڇ�h���5%h(y9�.�&Z���Xi�'j���`[rA(��^��mr�ש�����"�è_�~�Z������������nݝ���a�'1��6O��
���eVK��k���`B�` �i�F�
ĸ4G��B5��S[�s��`� �dHU�&. lB�xQ�E����C�f͕8���Q�p�O����P(��C�ȿb+��,Pا�F�*9m�����x"���@v�v�A�m��-�߮oc�ۭ�e�
�� 7(��ǒ�ޜ�[�~2� Ϗ���ж��&�^Hsq��s�HUp���΢`S<O�SG�Ȁ��w��1�k�|ɉ���m� ��RYJ��$aZ����&�G���R@P�a�_����{a�9�F9�{O!�z��K�8>��w��,J$���
9�f����_������Z[ѽ7�����r����c��{N����.vDT�D|�(
1��+T �K�WR�l;�C#H{��O��vhAoȮt�6�O��KL�,�B�/@�<��9�-PI܎�{j�ա@��`z�a%;D$���mFL�ja�&�N3�s;FYD �P�0�;�f���[/Ym��=���R��:�}r�NBˏ�-����yc����1�G��Pnr|(��r��SE=�-'{�SP�����`��&����t�^?�F��ܞ �o���;|��	�`�y3�ޱ���t���x�����߹\ٮ.���� -�΃y�F�w��@
������2�Ϯ�C�D�d掙�4̎�8pU���t�ek�� %:��O>u�8WaAQU����_r^�;OG	5���3b$E��H��ߓ��,m�P@�I00gwu@����3�Ĳl�>�Dޢ�""�!�@wSO�On���+~����5��~71l�����<�;��#1׼d�/Lgu�|.?]��].\±����:+>�gg[+�Ya����1ݒs��4�NX��y�����,�s��#ɽ��I�.�AH�L��ݎBDW"��&�M[��q�cF�!�%�^�vl�(���U.�sg�v��n0��v�u���r��|����p4��#�>n�x��Q�xv��c鐴����g�����BZ���񯟋ۆSi�֏"I7�d���LМ�/!���?L�0�6K`˸+.N�L��+�e��%�+l-��������w�s��i�Z'��M��9��Fӌ[T���lT�9ĶO��G��$�G�s�"My�؉�\/����Xf���m�̠�S~6I��2����!�;���ȤCi�=xc������%�+��O!TO����])-U_a���Z}��\LX�p`�Sf(����؞�3a���)�����B,� 9���7tOB�ɹY�^R-�Qa�P�`*�H�D���-��quK�����1a�`K+�x}J�Z7b���jb���xW�!%T�+I�V9��� ��W*$��`�s�-P��b<xk����=��j�-K�������UXB;CkC�ב�v���G�~SUC:߃JR�3�8�3�+�d���[�x��` '�eQ��ӱp`�Wɉ�z��9�mҫ]t$�Pl���2�	�v�eU`>%��|S��O�VL{7���	��K*�-�Ձ~.a�X�8�"� ���G�����$?�&&ֈFp1��,|�� �~�H����k��������J%�Y�ܒ�
V@ť���I�V�D���.J٭�AS2hU��4[�Z3i�Ŭ�	�"@"/\�U�W���D@���ά����r(��31�j���ҕq�߁$�:+��[�W�u�}8)����H�f�� 8X���m�u�o@W� ��5[�]��h��7'}x��dC�C�o�i-k*&���F vИ�Z���]eqb��}LCś�^�^��/*�"����3�����Cx�{[곿~� ������i�K�%u�j��� T�c�L6�����"��b�l���hG�jr���N�=K�͊��6�y�2����q��O��ҲMq�X .(�ۨ��N�0��X��%������0���)w)7�*�mF�"�1M���C���z�<�e�hE�Ws���9�Xkr���v�L�3s��-rv�����̪ttC>��hK�2)9w>UΗ�����ΊX���b�����W-G��s$��?|�)i��`����d��P��s�v��m
7��E�����n�:���5���i+�7��P�rr[�%E� |`��׃~:��Xr+�y@߁{�T���745�����r���8����dV2,�s���t���,��=���t�3J��V�*�w03 ���fL�}4��T�_��L��[�9��� L�[�0;�+�~�V��۷����C�GAt�k����mJ6�"�+�YG���#a+-�L������&e�a����y璠��<�P��.T�t��.�Ӣ%�=�3�I�^��J�,��:�td��rq����$�^?�xq�ԙ�b�E$�6���~Ad�D�x�?��B�hCs��f����5N�p�h�9N���3ƲDЕ<j����z�\�:�

�x,rњ}�yb��4<&A,�!�H���V��)z!-�O�mk��&#�����er�U�,6l_ �D�>\!�������]��3?1�!j��3�`v^��d!J�g�� f��%��p�S�*�[��<��.u��+2�L *��E�'_] (�V��yZ�bH��(�_��,�Z���.�7�w���������{��`N�!�O�zfO)��Q����OH�^�ԥ�m�%�^�p+C�C�JE��NE��v߾��bG�~�1����A��1��{;�S�d;�9UͷJq?����Lo:���R�.��˽��Ū}P�g�6�̂1��zS����`V�Y$�Z�#3\���A[�Q�c�G-Ɗ��v|)�54��p?�k4
=�\&����AY��s%~���)���أ�B9��!+򅽦1H����=R9e}71����i��Oa�Z��vg��p�z�4��I�e�tz,��CH1����i��v(#h��(� &��~������q�P_2�m�{����!J�՚U�]%��2O8���6�c��P@�}C$�I��V���N���ʬ�B�*>�#�M�  Ӻ+y O���'��s�v_��S���>��+k��*�S�1�s4�$ǎ�d|�ΰL��]�s�5����1%VM��E����~O�S//UQ��6�\�|P1s��|Q;�暈���?`�x��N`�F^�E�Z� ��|D6���]B�~���WQ��I䧌���Pn��:���z������:���m�i��x��9H����H������Y��/�@�/Rĉ�Ö�� ��L�y�܆bXfpH����6�Rb�a�K\t@����Ɣ5v�w�F��W@鎕m	��[An�[�������B�G�ٟn�Fз�Z ��FɏX%}�D`�B�FB�b�&��o�V]B���1>*�����VT]#BwB=��f#�)G_ ���(.7����&>x�K��P�]����*�y�;��U~i2�/�Ӝ<�+͔"��C�D�W�a�x>��,a��_�AQ�f�*�A�z$Z���٠�.���Ը����z���qm�������R�����u�@�U�޵��=P�$UxG�*����k���#!w��ܝ��g�scI�p]@������E��>_$k�T;ނm�n��(&��%ĉq�\��>����q7@��Ԗ�a�}��b!ۇ=��h�ЎDVɜi�����S3���Q[�@�;�e�\Տ��ULa�fB�J�g�o�u��Ѻ��Q��U�7ɏl^G'E2짛J�V�:��\�{�P]� ��Q��a�0aw���;gCE|4{���כ���jK�U�\Lw�{���e+JY�Җ�H�$�~𶭿	�����pj�u!��S��x�-K���(�03�T!��L!#d�;�O�,�h9��2�Q�O)g��;6����L�,[[�x2vU������L^,�"�gG�Q{}��L"�6�7����UL�=��-T5�=�|K��"[W�J��^��3������[��E��B��T}+�������ҵd
��nN7Ui|~z6�<6���/�{�u�6f@%�]�M�`�_s����[��GE5�K�e�*�6�������}�/U|�u}����A�й�0b�N����]۝����O��T��vǋT�?7�,.�'4V���b
@NC�^�DT"�����_m2���� x��u�,g�]���,8 [s����\�7��`C��G�̨��1�&�X&SH�H��?&��+�Uf���[���C���aB<�g��{���sSJ#1�0�~��u}@�@= 걗 �GE8 �Z��GC҉.�j�%��F��E-��ӳ�p���fE=��%�#��6,G�pwW�v�HI�*k�{�&���x#��т �A OAKH�=����o��;)��;nj��b��r{��֟L`��Қ����NC���Фi�Ɠ}���:�<1���v]F:hv��n���'IGB����c+ծ\��)<��'���S���� �hs�' 6��1��j�o�Lr�ӯ1�!���\�jO1YU4R�v��:Ac
GGA��t8�z�Ţ��W���vpޚJZ}���߂_���z$3��S�o,�km(�Ǡ8A�~ ��qS�X6HY2�l+wѳzl
�(f��~�Ni� �E]Pqk@�,�^�s��wM���.i�F����6�^ ��wC
�t X��~�s�[j��;���E��E��f�v#ʓP� kVz޶I<N�XF+5�k��H��%�X WGI�b�M���:*}� R��3�sVN�Ad�Kх�e
����ֵ̾i�4TrYћf�e����Kqۆ���&���;���63HU~�X�	��3�>h�G�
@� ����RF�8
Ŗ�E�S,�#�o�����o�\׻�Q���#F��K�v�H>$�x�'�=:�H�܀�=���f��)��ӿff9czI��Z��������HP�_��P	��e4��A���u��=���6i+�@� ��S�(�����l�R֔G��=���t�祇����}��0������&~G$jb/!�=�[�G~�0�R��)BOћ���ޖ�ei\=p��xdq.��C"e��YM�ы�7��s��į�����v���z,�B�I#P��l���O�'��ù����⧣�F�8?����.`�qǛb$
��L�S-[`;뱻��t���-Ӕ �ݎ�K:�U (|N��f'���o�wJP�Nw$����:>�������X�O�W�Wc_F��V�b�'��ڱp���@!-��W�z�!_�D��Ii~�pn������z߭��1��~�'s�B֮[	B����vE6�®e�B��_U5.� \"�1�t��=�7<C*�;��|
�}[��8>	Ac
����7?c��1��wo��8���Ԟ*��gM�K5�kl���E��w��K�$�#�Vw)�z�S���h2�!�	���C
�`��E�9�%����맽��R!d���I_.Qp[���w��w��ZU@Y�3�n����2�^������n��/���1�8����n�@���H�ݰ��:��k �o\��bpD��'� ȏ��g\��� צI��3�K�mI6u�L0�i=��K ��XG�����(�~�t�n�Xh`����-�m�R�Iw\���)�"4�Ἴw CSV倷g��e
�KEh�^5GD�m{�!��b��I'��c�oF��W��S��<q��x}eL�-��Ͷv�CP���|G׀W�"H���)$���0���5Q��;Z���A������e�R.��p@�ʆ���vB`���hΑ�ޗ�6[A�(m�2�����t,1ɠթ�|u_�b�P�1U����>�玞b^X�����]���=C����s�^�W�¸�>����]�!jG�VЄ�_�5�yU>�0�c�?�W�3w4l��Sz)���WU��B���W�)"l!,c��=g���2�/�g��2~��i���`M���9�]��w�&�]��(M8�3�?α�u�,[�yr�֟��fy�,�>P5��#���H8�5����x���S�Q(!��+ ��=��&���US����zZ����|\M�tv�ZΙ!�� _y��6�{�@�_w~��gp�L�jfO�����JSg�+QY��$��DzL�5��4�Aq��[5ʣ>�h��=.�zx�����L���,9����c�9�հȠ1$�.��U���f*�D������T����a��/�*��+~]��|fʖ��������F�;���G���ｉu�7!L��5��P�FMF�G��l�q�K����X>`��ީíPJ4�Է�|{) ;c�2�x8��h������f&9!��^���OT�� ��U]��Y�Hc: ��f���vtC݉@pJ-��R��ϐ��sv�L��yϭ��ϟ�����H����e1�鐪��V+�ӭ$�����f��51��L+�h���)��o�.�����?d9�:[�:��a�mR򟡄���F5�'V�rB�����N��*``I(�7�b7:�ְŲ���l�~�JK|)��ZJ�l�����y�l^��,./I/��Dן]�L�˓�b� �x-���
t���v_ f��t�yu`��&�1�ie�n>Dw�q[�~��s!�	?�dx{���&l�_�yʈR6.4��Y��J� �b�@! �\���m��&����^��=��o��{�3I�:���c+���ā2���Ac�Rd�#p��u���H�Ne���7����8�.l�_�KЅ���N�3J^]�*-����=چ��fdNj�\;�Ŧ0V֔�N]pr��~�މō����"H��z���-�}�O!�F+��
?�n�~�z�js��٣A�Pt3��9I�mtI=��)�ƄXn93DA���"�}N~��uaw߸��?]�K_�*�;@��΃x_�Ee�tjT�}��0mM��y���_��͹HAvY�36�m���- �!"N������/��?��X�r660�@��~N1n���`��vm�2����`�~�.,�Wޙ{�7>*�C��d%"`���R�ѡ|��TJ­�t|���)����z._<p�M��ڨkb�X�D�o!z׈����nS��h�ܱ��ښ��ԡ���A����ܷ2��H�v8H�����솯D_̵�RF��2�C��Dق@����h���eep݉�b����o`�2�^il6�2P�nJHt`�q[0�$�k�^��>�&|@�>�Վ@�� qg���}Gt\;��xL̟��v�{?G3n����T^���;��u�,
���>�J58� 4� ��|ԵO#�:����Ð�_�L�7�2�q��M��c���0ꁋ9M��C�8H��-E��>�#��W�f���Xb�(4	�<0d��_�zNt�a��%twVG�<�_�q��v�����)��z�',���2X!|�a#C���M�n+�2�*��Z��F8�:����'�:�}~"#��/dvs�`^>�]�skR\�4��y��Ha-PY�yK�>�����) ��LL�_��k�d��i6������N�;����y��tD�t�"�5�|	�ٵk�=�=3�����3�]�o�S���f��̚,���gT�'�Q$��!�|�[ֶ�}������[2o�i�ߴ��U�0_�n�
n>d�w�zE�A�q&��a��k�:�ZՉ�/�j�(�8}M}'�y�� ���.�a�')lC�ϺĴ���ox-��dL�1sZ���ϙ[�i]ښ̽Qϔ��s���M�y���+	5`}?A�^���������Y�����`�N�(�#��6�dl8p,N�cc�q���Ru��y+|�G�z]�_���q���1�i:���W�J[�mC�L�M�p�;=/h�nu�:4��Ŕ�������8�H5�A�A���Ň�\d�����Ĥ��ʁɅ_	����#�r��c]��o�	@����P �"��y�p;{�񂁻[t��'�%7�m�v�b1 	���ʗ��K\��7���}ꚳU��į+Fԛ�ÅdiO#\�e�
�D-�׺D6Üoד���Ee|�����w�Og�D��3�����&��x�H�N����
����"_S�
ݎz+���nՇ�-�q.��.3�ї�p�
�?v
mS����`%c�V(g�^�`\�ј��Rf-u���0��ˤxP˫�D|T�4�aʹ6�� ���Y�W,��?��Go�;ډ�JV�B�y�;i8���4����Ґ74(+�����@�H�=���\m�[A䈿(埾^M9P�΋�̡�\�����f���]h{d�W�SR��d��
��i�4� ��mj��g4���$�xA;��D-Yd�N��xl���y�S�s�l�l<�ͪG���4�Ve��KJ���eIC�@C��f2��n�4y T�޿H.Z|̛V��a��-m*�)_l
���%XA-r�c��mct�'��E��mY�~�n�M����lt�ݺ'dJ��R	��ӎ��u ����$Ʊ�K�B�:�u��OS6�#�Ղ�9ݪ�Co˦0���H��|̳5.���spB�C�i7�:��Ǻ���lcd+穥�~F"J�52�G�K������fS����C��2D�J;-<]��a ��$���G���-`2�-<�Ǯ��EA�Y�Ų�5�� ���ft��*�zš��Zy�(hL�ܚ����ESZX�mǨ�*n���]G�0���Y�=H�o��N��y�R��jGҸ�]�k.��Tvk���.���B�º�{��4Q��g�i�;�T�FF�E:�D��)X�Cն���<�޾�uaE��5,�_����J�0��*��UA�z[&H�.�B��=���1���xw�P�F�q��44��D1�i	����*hˋ��C�[y�ڬo&j�u��d��y�u�c���Qhϭ��Ŀ���\��;�+�)�1�=R$��&
>
�w�7�L����B$�\H� ����λU�8�m��9:������� �ƴ��q��&j�(��P��.Kǆ��İ�*��"(:_����t.�b�D]����(>��L�?�~����}�IO@:9% k����^�Sΰ�@�F��x���<�a0?-]Æ?���p���"�"�=� ��|j84�+��le�ʹ����a��ܪ_mt��a8Ea��}�E��"�d���cAoCt�}��t��}��h
�\��$��`Ibj(t�t4��oH4�EI�����Ŧ�$m�8�3���jw�o�a��'C��j�.>X�-x�8W�Q�����O��ѥ5�3�v�'�,�`mR��V�X���E�Q��P,�E�ى)���UKm���N���
R��H�M�k�����C5���HF(6o�Ȭ�aT�w�U �'%�mB�����64�w5Y�:|���UB�+�%[B�ԃE\x�� ����	�@븶ݖ�O����@�[}�iڿ����������[4�������;�H=��Ż+[�#�m��#���DlBda�_R��j5M󬾐��ԭ�|D��h�i!����Y��BF�g���Q��;E�zR5��[k��� �M��HQckL�����s�/B��3�x!}�5�Ǖ��RA�0:J0[rPX	���A4'�ax��yk��jkR7�<$L��ظR{'������ +�����q*�����8�}H�y�����1���<�h��Xޮ�"�i5l�'���G�]��a0���nGɵ��Q����{z���8VTle	�'RK��Շ�T���達�y/����5��U{>�)y���`�:�=�N�7��|��7�>��oh^�����yv[笍�+U��O�J�mS��҃V��b�GMa(p��W͕�#�O"k��(�I�D������Bqs���0W�C���U�@���.עT�,$<�oʝ��\��Q�n斩o��J�c���w�{v��5s�&�z�|ZrWӅ�SS�S\���/�qUq�+�\K^��?���O�0��.�@�5[���R,��CA�O��b�9���������D�jB	��KY�}�"X�Γ��=�Ze8 s���tt��B'���M����Q�n��0ލ?Ֆ�^z���J��a�&w�<��2􄋫%��QQL�H�M����S�c�i�e���|e�!^y�2���c��6�|�����E*T���)|٨q�(JR3ZH�����'��a�ٞ+������sV��x���<��ZO	2���9O�a&�־��.�ϬN-�"+R.�\S�xp�N������W�d�B#՟>��>6�U^/��<|�bfޣ��`6�%h�.���U�i� o�F�q����-�� �;)9�9��%o%��bIY��F�Am� �".�9o�o�w�m��nci'��@-7�]&��S�'�3[�O�F�M��t��c���d�r�?�U�F�� ��|��'�A��Y��&W�'

X2O�0	������/�3 �ђ؄�^[��?�r���������wBJ�<qL�
[����jp6�Zr����X����'�0�[�x;^���X�|�DP���`Cn�'�E��~�����kx:1���\���v؏;(�l�:��H��x�Qh�"�-f�,Qъ�Xj`1DTС�z����� 7	�y�m��ķ� �k���GSa�D������[�PZ�n�*��� ��ĮO0k%D
�e\�GЃ�̺6�@��J��D�n�@��o�H�x� en��k�/��1���4��7���v�ɀt_��~�t�/�����yc+)I!�$���f8��2���h���(�&rg,X�m8 �w0.9̟tQxHA	�!�r���l�?�"n�*�$A��p�Iz��|@�N������Qp�-��cn�+u�E��Zc������uH�K�3L�٭˕��r�X�瘤t-{2�3	<�����UK��U��G�y3���8|��
��>2���9�z���������r_*����8;�G��Q9�RG��Z�K������=�V|�E���Y:)�Du������
����Eu%�Yw�����"ìփ�Ь�N����|���JX���x�M���5������-yk�D�FƠ��n�fwcvYq��6�>�W���q�\ke1�v��;z�J���*����
�K%}v��S~gF�4�@��@��څV����q��#�)Q�KeU�Z�y�^���>U&*����'y�?C>�h�3:{���MY9�A�na��7a���/	�&�G�aT���}q(C���o��{�(M�:�]����=�qn��:7�2^�$k^Z����kY|}��wt�W���L�h(2-�F8��\L{�0���l�z$�m;�jY���E�]����R������]2�o\
�ι��H&���L�C��g�p̀�R��/�3?��q�:p]�H��r���Z/�9��dv`*
Ж;0�\�?Vs�vaKD���#�����P�R�c�kQՆr�(�Z���9�u���E�2ܓ��g*������5�yx�S�9$���.VRu��eG�Q��P��8Z��8����E�,s5��11t[���'	�"�`M;�d�~'o�.��
����7���t�<�7�p��`!z�Lm�;�b)L_L�j���'H��J�]22��4.��oO�q���mT]��֍p�#�O)��CR8�3L8�"׋��!xe�}�S���;�'���f�
^W>&�.-F����@����2�0O���{�盯����T�ba�s{2����S�\�����Ѷ���9s+R$���	G�,ǩ��2J�hS/��	�Z��^��l�{�Pj�Ĭ�R����n�`}�2�X���7IyI�:��CuG���~Et��ٯ�0�k��^�:ʣJ���7���%��8y�l�,�Qm�������`v�(WƟ��e�.wf�;��Z�.#��}X3*�yu���/��|g�+���g�THMv1ӕ����?R0�V��^<W1��;�Z�>K�[�m������/v��Ü\%�/�X;�=������|�p��obJ^�ˢ�ב��ÆW���S_޺�2�K�Z�:�9�'+�	�4���71�޵����߼I_�F�GiX#�4vJ,K����ϭ_���{d��|�s��p�[%��.A�!�r�.a�X�I�Y������n�mM�2�:�W�	=��w�9J9��B��z�;J�C.$�(��4���|�����&�c�߿a�rx��J^Һ�f	�'R񮐨�K���_��hh���{���� ��ɚt��`�G�:��~����3���s�z����LG6�9{D��I7��1=��0�ǂ�*|U���� �jbE�>(j��v"K	�_ʜW���ޫ�X�{$g�Յuó�Mb�x�Z������(�D�*��d@�?���[8�h�mo\��ƭ-2�>��b�	o�¬���nѹ]�y4��o���
~]q4�ս�g�b�p�#�JY�SRm8o��9"������eq'4�]�U~c�c��E|n����LHF6�)�v���~������X��������z¨ͤ�.�L�$jes�OE�u�Nט6tT���u��m�GrO�=ɶG������tgp�$�����a���
I����u��%Eq e����te5�x�C���xvc@�1s�b���(G����1N��oMȈ>�bM�R�_!�a@�9���ōv��=d�(2�i��Դ�6��f�������B"��ǡ�����^��������}s���A�������I��wL��>R���ſe��B\�:ٽ��	�(J���_�k�?����_e����.������>p����Jo}(\f}�!I��*3������W-Yb��O���R���iߋ���	f���{�H,��&@]S;n�fE��mT���K ���=f>�Z�w\�\1�.��r.��� z`5�Q(�H�ޥ��=�'lT�>�A���\y�X��)��V��ѱ�Ġ@T�b:K���NC&���`�����r�����y���l��{㟕N�t0��NQu ��1?B�:��'��W�����%�����y�X�{kw�iَa�|!�����ƣ~�Z�"�9 m:[��U�°�w����R��.���Fa��0v\��X{՗^�M%Q Kk;�Ѓ�W�|~8,��d]�C�<����sUkOz���-Z�)	�yBy|	�k�+����h�pJY���Y8��ƌ]�N��3����E̴9��N�
.��}ޥ{�"��d���q�����E����,�{X��܅�e��S�S#U\�r҇��mLR+B#�ͣx���_�ٜ���r$%5�1p~����cO޴� ��;Ǘ��iz�EVI�4�s����h�@��<���ȳ�8�.\�u��(��a#s�κGu)�P�*��e|65M`��o�\;��^��؃�m�V�/X��΀9�h*4)��rD��,�`���)�f� E�J�NNB~F���^�Ճ"���Ě`H��e���RMkΥͫB��˒.����wr*���{����r\���Op�uuI���$[���ܪ��;�����c��#�ӿ{��!��"�,���W��:M:�ճu2��ZǦZX������2���������>Vf�q^$Rhpv��k��̥L�Y�m10�Ը%s ��-�e��O�f�K+�<�-k ;�����kpi��7���c;3�vJ�]ß��U���]�s�I���x�8{��
)���wX����2	0(��}��������l����k[>ln_$(([Zއ�O��m�e�A[��&SrRs
:�?f�vة�����'%����8��Am.��1l��`�H#t8f���}����"՗x1b{);v�7Y���+s������ �u�P㔾���-�}ePn7�xųE 8Q@S9`]ؽ�b�_`Uf��ۺ��6�u ��������Gn��p��0�ˏ._|xk�6ȫA��/�{�H�] �N��Hcp
���٨�aI����*�h�LT�2�q�i�\Sk���I��e���BG�[�in��e挖�I 4��9ɐ�J�!����5��	Z�C�V�L��G�_ 4k>n���b_f�3�9�7����Rr�TlK6���w�k ��$2�Ls�Q/!�7֦B�p����V���]r㶴�x�(�N�⻿�Jg�h��a��?"u���[�$��	
Ls�F>y�Õ���zL�s̻B��~�-���Tӹl4.�t�U���Т�1M�i����c�d)�~��/̈{�^YKr�8~:����Q{4���u���d��i��U�.�糺���/�9t\S3�jKq�?y<h�\^�k�����!�V�O��Wㆻ&�O����5Q}��81���Z�*�����Ms��\I�i��iy�*���8��i$�h'E�K��m3Ԡ-�m��=�* &�sص��c�J���tOw0bdcl�_}�*�AXi+Vk
0�Xڱ�8q�(����C�s�ؗd�n��O��E(�������,׎׸��{��rUe�i�]��(ـ�1Z$��E���ny,��X\�q���n
���'���o!)t����8�r�S,h��}����=���b}G��X���i%��ϸ%;z�Nk��0�E?T���=##��h��h
ӈ*�g���z�f���^!�3�5P�(j�~
��7H�H��[�<3'�C]������3�۶Zy�J� 1�/��E�J�%Bj��m�hEH�;�� U��)� ��gY��#��N@����N~Ҳz1&��AR9Ҥ�95�J�{#��	���/	f���J���\�8@b�N��kB+�12 �����PO�1�� ��/�Ć⭚�P@+k�;'zv�9_7u�.]�uZ�#�hv�R��H�,Rd��\�6���m�!� �>er��wGH!��T3�l	e,�oͷ�IME��jx�A��R��2�*a!q-�Ef�,z3_�B��X1:�r����'�r\:V��t�j�SR����G��*�>��#P'���(��4>u$!��۹�$�`ۺ��Ʊ��*Z����F��덵�U�[5M6;�ɝ��xD ����h[UL2|�֕��c6q����w�ú��d���H�(L�N�د=oc�p��a{��Qa������mI2q�
�oH��]5�o
΄Aؠw� !�޳�L*,�7w��n6w��#L�.V	�侻��{:=� �D�G��`e(Z�ρ��@��BM
X�����!Vgm��s��x^ƅ_�����Y����YL��ؿ73-0������e���p��7�9bpǶ��|����CP�nb�!3�98\\\՟)�oa��X����%UE����d��BB�5��}NOY�� X�JW3�gӒ�&"��K�a-���U�c��1������q2J5	��߅�G����xWnֵҬS�@����c&�w?c%X��䓧t�=9޸������G�N�};�a;$�v	k�J���Of�'+�	\+O%\=�+P� �`���`AoJ<���{���S��Y�p�JF�������H�9���*�$I'{������r�l�ĩ����L���&�XB2��W8S:�u��b���F%w[8��z�f��%73Ņ{&,[�O��/e>~�q��I��ۨvI�D9���d�J9�֕ո�<J���-dw�v�۴8{c��	�0���[�lnȜt�����E)$�n��H{�0��f]���������\^",n��M^s��HR�IX����i�U=��|uO�:�];�Fƍ�ʷ2I��c^�ߏ�}(䩰T�� ��=�o����C� ���d��A��E1�-�jQ���]�^�I`^U!��cO����?�N�Mh/����v���Q���I�����j�ljQ���/�L+�u�t�F���J/ �a32��g�,��X���s�kڂf��	������5`D�5s5��_ڿMA>���c�K�|��đ��G!���������������qd��*�y=���w��{����AUcoH*k.��$`���U7�.���'��R�sf��^�/Zf崷��Մ�T���n����.��!�J�<�q]��ҋ�v>Χ5T)�_/�c�&��rh��$i���4ȉ����� ���u��^7u1h��,׼��=,�
U�a��P���!ٮ��8�6������:�gt���ǜ�r���틦ħ�^̐4e2���%��Q�ށ��=�N�(
�� E�A�r�ǘ����_�T�#T�A2sq\O3E��`��	X�.i����T�m��.O��elJp�z�V_]6E�w�Y��ӻ{L2Ґ V9[�e���������`#�+wi���)>pr�WZ�x��)�vϢ��N������%��I�O�;�;\^Vk��u�WH�|�|j���Ύ�� �QE���CA��<��j�������L!�לׄ����/2әfd6�S3kc�9��x�I�u�?�RdXFL̑ݦ���^T�/���r�5�>�\�1�-V'��٤m״��oZ2�p0��=�4\��I\E{�>�9J��K���-�g̵�ԁ`�sF�t9t�;α�E�y�?PG�{��t��I�O��v#�j�^��퀗��X�+��l�i(U�E��\�ٳ~v"�Y.�P��8�|ΓD�wNM����CYc$IV.����)6f��Rƞ���@�\��S�B���>\=t�z����P M�;@"т��@[ŭ iT���T+#�.���p�rY���V&0�y#cK�J5/"w-�S����%!�Q4k�@�K��2l2XN���ԠS{��n/V����0�]�a����'��B�a�P�������MW#�^��Hx����!V��Bab<�I��W�&d3B�d�7i<��NrD�*����(�I�"�{��BBH�	lz6���s6��}uJQ������dO��$E�]��5�E����s�i���D��h�g"��� ��̀�+��1/���	p�㿌Q�u����aP�5(֓�{�r���}���`_L!~�He����L��M�C��/`KxNH��Ț�5�����g0��3��_H�E��������@༠�=]sAAC���ȥ)��<��z�Ѡ=x�H�O��m	4�~�	�̑T��5˸�Xn��^�GNRzN����%O�=�L���Vz�t)����9�Z"�܏q�2�s��p#��涅U@�#��4������c�vC����`@B[y���^��l'ib����s�b
IlϚ���Ú[��Y �ܑ������!5�c~ t�Q����_1��}�*�#-+�|n�"�D7�\��4U���@	Бĳ*|��o󦋗�c�R��������1<5�qhV�J(�Eū�d6m�C�� �/h^>Jm��b���Q]A��d�xK�S�c�@�yDO0m�5�^ʳ��Vl�hS��,��(D�*��I%�#O֞��sZV���S�s&��+�?q�]����gYsΓU��弑�b9�"�e�Q�0a��\�Od�(
&��z��yD2yC���w�IR[�;և��ڤ�S�Q1������>-�Ɲv��AGFO	�A�8�]��a.�N���B=��˯�oȋ����v̋SR�7*$]dl-� }H-�?;>�ܖs��Q[�Zpg��|ym �����y�y����F�ʍ��:X�RW�ս�ˏ���-iTOj6w(���6&�?�ʡ'�R�ַ���gl�9��zU[ĵ�>՘>�r۔C����!t���r�E�AHس>�J�+/>Vya�������H���e�}�+�K��R�c�S.vP:�\a|��	�$<b��>*02\�J%y=�����r�Hce�ݹ� C�3�A�Ѣ/�|gbg����)G�K!����4�4z)i�8���ZW1 �/�����m�8���� �*���S���:IJt�n�������lY�~�.�A���\�J�J���k"�	5|���X�j�^wS�x?��ɂ��B8�RY��󠔭G�XZ����/�0��r,�>T�z�g�J?�.��������1Z�k����������/<���c'�3�+�
Z�6�n���5��Y��v�P��#S�:]��5|��X��g�?c�&hM��]�����k���U�m�Zr�4a�@���d���8�'5~ӌ�z,��G0S��$O�$^[��\$0O��Ύ�0���.����M[�m~��?�[5ʻ����$'`��<B��)1u�ey�S���њ��]��ܠ�B��YO|���6�����7���&��A�_�E\6U`�VE���\C
�_�Of�A��%�V���ҘkWᠰ��IxE{�|n�FxѰE��KKA^c�Z!���Ãt(�k^	S����x�BuD�漋�,�� �Vd�6��w��ԄE�.��&��ǜM5�N�w�Tr#�����	�v{�J@�� p(<���ِdsqB��q��&��!a[Ɋp�'��t�/N��&�(X��y�q���k�MGG�����xŃ���ly)eO`��&��ׄ!���I&g4LB�Q~��,�	uyT.������C����5 ���ˆ�)�����ݕ�<�֚��}�c����2�D�`� �&���l�kt������aMk�������� ��-�S���x �^�t'�Q�M�g�uAp ��=(�3�Ԯ{7AH�sl��,R\_�3��`]vby?�U����]$̹K��T�c��,��~���\Z���Ko%u�,X��8�s/osa���b{���e7d9J��:��&�o� �`c�\D���MH}�u`�s=l�V�Wyta�H]N1��
�+�N� b윣Ҹ	~�a�Һ��w���Q�,�p��r�5�4N�seu��Ғjي\�$������/�H���˚��^ NM02uxA�1��@�-��H�/d�W�F�w%�@�y�j���h��}u`!�4ņS[�۔��f�}�ZpI}ıC{�3�y��R���5�DՒ����ـ��AU���:2���n&�M6-��L��k������C��+I8ŀ;aR���`'�vŎ��R�a�T���=��O����	���8�4�yŶǀ.�*Ҫ�����,�G_���ޢ'�~X�N�OCTu���[��F�r%���a��o���{X��-��K����]�ba�P�%w��x�{����qZ[�lL�a3���c�å�k1G䝖������ϕ$'�2���:�5P��f[3\[ݥ�R�Z�a����-�^:�I�	�������]j���˃�y�
V���V�m�/t0��f�dH)@�r����oY��Bdk���q�t��J���ٻ������4)V~�(���L�=��~�Y�<�Q���'�3m��3�J1�\(�ȃJ	x7�+p�+>�!��s����y��f!S��B?;m�/�v��i��jak<���N}p�\�M�'������t�@V�r��_�B)��]��i�V.<rۀ�ܨ�z��d���Gb}L]����ftz��$�&����0B��gV��)�ZmGՆ����]!���^��2\8����+�x�w�G͎]��ߥbJ��Vya0[�9���Q��j�+��4]hS�T�N�8:�Q��t�8�.B��%�;�i�[eZ��*I�	ķ|����-�DE5l9M�A��:���'�'ѻ7��S�љ���1����Q����"Tg��/���fk0���r
��̶�d��	����v�`�lQ9��jv����9~����q������A�o�@P�$��}g7��mV4��Е[�{r�[�����J6E�k���8&�wgͮT� ���1�=�Pd��n|� �W���ʘU��8�J��әp����P��f'���4��S
�r$7d���(�T~vTPH�z�6�����ol���[��c3v�~-?i���]!4�0V!�.�[~�Y��aeMd(}�k�_�p���Ta�h��8�M��c(s��x ʟ���2��Цw�1��)����A��z& ��\�o
�@�3ƛ�I���L@�'���e�KNFJ���x��jt0����+�|�T��YAc z �y�[+R�� �i.B���}�k��@��C-D�V���Q'?BOB�\q�OX�o�ׄ�?�?�7�|�l4M?Sa#��E��`#b0�iNR#T����7� ��'5=kQ�Q5Q�.�t��d�*�!�|�8�y��$�tȓT��it�T�ڏ�$�_���������{��hN�+/� �3x]� d�31qvKr�\.��;�	�Q�I��/r*fĻ��zW�"˵��b�\L�n�N�w�X��k��\-��9U��B*w	Zȡȩ+>����N$��ε	��ށ8����S�����������?i��/$	����Q
��P6p�u�;�n��NP�H��YVb���a+���2��[M�h�o�%*0�u�p����$f����Jc����= \�mv^�%r-"W��_f�,�둠5��8%�]�bQ�*���aC�'�W���́EJl�t��B���;J�8����	#ީ�7ſ�k' ^@k;3J`�e5�o��AVY�s��M��]�q:��X�g�n�y��lo$d��[FiW�tB�⳿^o��i���jÂE��i��Swv�ll��e��a�E�Z+����h�ۢ3ѷ�P��x.h�[xH�j�D���l.^�3�
�C�ӗ{'TAM�Ӿu���;6�zj�����kǣ�N/
�`+4�80���'=�ܟ/���f��1G�Jf��X�x)i?�O���M�%Ml�gG�\�y;˪�k�>�2!M�vj2`;FN��%d_m�cǬ��(��8�-�@e�2�L�_�A�e�!�Ğv&��P̌jc-����=k�46�̎��>��{Њ)� ��4BF�����c̆-W�S��,��1.`7Z�J�=�����bh[�D�8�r�_r�=�z�v��?��d��$Y�5�F�`������D8�-�i��I��q��'�NTr�7��X�I�H6���#��=��G�{��l4
�aK A� 	�bOX�>�6K�B!m�TZ�6<p\�s���|}B�f'Hfb��X	��ơ��j���o�֩���򆣘{x���L_�ڧVض_�,��t�t�DV��7y�f&�7?^�"��`�Չӂ�.��h�L^�o��5?�Ӿ��ֹ9�=,���T���Y����N6�:�^��o��$&�Ǆ��z�5��D$�'��`�+�g&�\�m3�e�
��
5[��in%g8��+&����s��Y 4�4Qek^����CDL�u�<
e�4�V��%Ҋ]̙�6*ђ2C��� �U�7�Tb��
tm�Sd�=�2�A�r�3��<xs��5�!��R��Q�T�1�r�U��'���D`��{Va�2��"X?�'���9O��#���;�9. 7�R^	���O���`{���{��� ��������>g���Pu�Z���*l�4��k��#Z����%�@��N�T|�V�߈>��`�y1C:vu�ƚ����s�-�a��	-��f#X�#Ñ/�Q��%�D2�I/9�wh�	�uH�����T��Ȯ�ϘY�.���ٌ�#o���ʛ9�`�C��o����y,P����n�rAC��ώ��ߪ9�3X,�YIMwj�L8GN;R�g����I<?����a��O2�]�NC��E��U��.��F��@rw9uy�T_���`����b^G%��>2�'��]W�S�'�4�_v�.����5v��u�{>�^ɅvW�F��h)�E��f��qN�5�nv)ܟ��z��#G}Jhꄏ�ށ`�U4��I����sD4 �S�L���讆�QK�4� �zB�	L&��Zj4E�)VزJ��/���I�d�l����n��KvS����x�[	�,M;v���q@|-5D��qu&�b߻�B��j��ʼ&���x�w^���-m��s7�}���a�LUs (���@lkb��Yݯ�Q��{ǵd"�4�;�t�g�k+B��@S��q&*��m-u膿�ʏw%���C?|�߫|J��ڊ�c���	�m��; ;��J}�IHDB�h��ǚ6	�����?%�t]����9 ��R��:4u�O^��&iwFSە�������m�˴��G$�]���?sa�8��Si�������{"f�\��M~\��<�s�6yRF�b��v���!�Q�靸�~VU�)TT��rԉJN���=�7ԋ��1��hwnt��=��ϥ�v�T��Û���}��J�ژ�bS(- �4���"�n��n���k���U�=ԅ0M��A7��%	K�j׽�ܧ-4�P�+�9�~7��˖��8> �"p���8��[�U@�{��{��l}_��W!j�B��N�k�PB�¡��/P�����D7��'h��?V���VO��<�3d��Zx�ܒ�� ��y�(s���/E��j��D\�q��-�x�����c��V��;��ٜ���@)����f[�Ҳ]��Ӓ���-xK*��T�2$yY�Txڙ�q���E[������p�D[��F�7O�Y�s�7����7�:v�I�ڦ0n�b�X$f^��^nm���c�����.JL���۰^]�e$��k�U�����N��{�+ƃ����T.����O78�E���{%����; @�=�z¡��m�Ni�t�[}��L;M�y8��' �`H��"�c �x�@�+��?1��͑�jq̙~cNz�krd�P�=�_�S��l�-�tB��"x��K�Q��Q��Ge�w1�	g펻;�����2-���#R�R���ScbCtJ�Ń�Yѻ���0�j�0)���;�b��Z�ۿ�m7v��{�"�p	�j�n��
}i�X��$%��%�	�!je^Ql�!�U��,�9�̢�:�V�g��.�#u	Zj����Ng
���3Z�X�Y�$����#&���z���X��M����z>P��'����&C+}��`��D�e�7��6�Ğ%��q�TH��y��8����=�>G|���KݔA���u-��R��ҽ�<0Tk�n+��S6
�f�i0�+�R��4r����;*�ػ�7��6�@@Wt~Ͻ�'T͞�����U~\�q�Cl+�N=O���.��-��-Z@]�2}�����:1l�x��|�
;i7���0��
;�ׁ�����Kɬ�K����r��a�;���0���޷�/�=�n��2v����_h��dp[��\�h�D�=��S�:|�8-�d�lM�#���ᏮF�EO ���>r2e�����,n�k�1)��5>���
�/���^_�!����� �c:$LZd��5��z�ͻ3�⿡[Ż?e�W��,%����^�"���y�ۖuMPA��92�e[����܆6������l�7�;1�V��E��ȫ ������$���1��+�I:�v%y��S��E�[���R�ܺ$�������v��Y�%d�6� <2e�QA�`"�aS��0$�P�fi�i_F�j��zN���!�s��r�/�OR�&v�Ci��5H��T����\�%�;�!�1���Zrv���7�t0h�k7(����X[�!\���$M���J�%f�Զ�p�y2��=���G>��\��ĮY��2"�`*`Hڸ�C���{r���!OB&<ŗ��kX�56�:�|�P�]LN����h���+t�T�:�O/׮�-��:��#/�Ǯe~k����N�Ux&�BK�>����7xi�A�.�圦��K�ЪD��Â�`����v�e��ӻ�L�ƙ`=��DX��}��+r�p3L4�C��umT��"�z�̜!׎��"^�JQ�Hr|ow��pu����UDz%[�����砛��"tO�V�vI�i�^Lo�Jo��DG!L�'w͝_Se5GTg�#��� �ɺ��fr�� �C��~�W��Xsk;+��G<�uH;����\@�k�؀���Դ����>�Q�r�H�9UTzC+��ڽ����nO���2#RM���r�2�>�e3��4�qQ��h�$̬�j+H�g�������b�V$W\+\�>~�Z�T���D-����8�[�,ۂ�*�d�H�<\�����"}?g-]?�2�4G��5����,I���� �qkaS��)��Q�䡕����f�+�,z.1����j�ϐ)ܬ�/�\�]�\�� �˄�hx���IMڪO����d�����W��xA^/�ϱ� ��C�=���M- �TQC�ݢ�<��۞��7�7J�LI�PQ]�hֳ4��b���$#)��]�c-k����6ZvU�����I	�
~�1��ٗ)���<�2Ga�P�� §I/Ɖ^�
�^9i$��H-��2t�K6-��N���#q2e��K���o�(3mp;��"_�\9�J4��`�|��\�b�0{�t�G��a��>��M�	3���#�΁�r1I�޶s�*W%<w"�q�;f���}U��Z`IAz3}Nv��2��<�S���.��A�[L/]V39�#�?KeI(�a@n�ф8�9m{\πL�bu*���t��b@Z�Ga��q�;a��,T��6�S�ih)���P�����NNЃ L\ݡ����]��}�6��@�n��	0VuY�ϛo����W��tL R�7ױںPQ������Z�1ྛ?));��4ؘ�!���@ٚ�^ƥ]H�cF����h/Ù���c�� H~������B�����[�p*�_�7���@}M�(8j?tF����[����1��#�:2t�^���R�҉����T��J7 ='�p|�D���@��
�G�Ay9"2t���lR1	� �����"�M��{�Cݛ�%���O�6���xg�Ƌn�9;d�[ڔ��9���6�>$�n8�В��v�p�A\�/��p�� 1�H�8�,�h4� �ue~]&��8'����RW��&uw�J�R��T=��ߍ��C���J���������M\�S`�9���=������H_V/]V��s��)�_q�B����N���2�B����9�&J��$��n�i+�팞��ch�:�����1�<�}5zO'�k�/���~��<����쉯�`�N���a��6��\�]ʩ���(?^��`贞Iom�q���	?�c�BJ@Ʋo���%$e�5�a���Vѝu+�>Ra��{-���1h8�� WΣ�a�d�Ĝq���ꫦ5�%̥�W�N*�gI�(������	gi3��qu�O8~���K=ߑ���י�(�P�� �
��zy��D��wi]���`����	e�p���qΙ?���p<�b^3gR~��U�d�)�k㗯�G�2�0(�Y'������=	6�=?�W���N�l%���4�E�.��1��*!y��k#���K�lp�;�n"��ؑ��D)?�V�6R3�}��f���zV	q�8���޿ӫP끡�+�<���~��;�3�
-���n4g�\��3߻�f���3$J�9R��ES�[��j��7�6���'��B�*����D��z��E�h�1{���N�@xnNo?F(y��̒�AP_���)�����T�Ge��?L�`��P<�'� 'J���sd��<c��!���/l�;@�hD�`�Wb���
�������_H�x����%!�)�z[�*�PB���=��)iG�SfL���ic��_���g��sK�L"O4�j=(b5�ÒEz���?��e��},��\q��x6d�d�6D�W^�ǭ+EmM�8��a�p�<���.����M�\�e�b[���bc�!Az���&;�|��T=v�ڶ�0��|�+Ɲ��e��w����R�jp��A-.�����;f1#z���C7!oY�%M�5���<�+��}�rU���Qz�?MH����G3�6�����nm��q��b���@V�T���D�3}vQ��ZY��Z�x�O��Mx��f��md�hܠ
��~1/Ma>��,���&����U�B�O¼0B�����I��{���ZcB5����lq�4�Q�'u�G�N=T�۾�;�e��;���P��P-����ЊYH�w�����?��8==�d�rex����w�.��7�#��ysu������E�+$��~��n�6#3�R��W"�,�
\z����~�s��˶��CX:��%G'Y
���w�"B���|��_�f����cKl��%B��e#����̀�����%]�hj��~=zv:�k��N%���:y/ᑸ��X�$1�k���Q��"��֍�}e!5f�^�#<�7We�%��v�Jyj~�{���	�z�屇�/M����N�QA�"�)�,;,z�Jt�!RfN_�����	i7'�;/�a�:�:r��[ӌ�=(�0�#'2��ʦ��@#��rr���[?r�x��ŖL��i��2���ݬLٲ͉�kYm�e������ء�A�5؞X��/N�h,����==ES��O�Č�� ����^�b]�������j6�x�q���B�����1���np#�k���Qfpc��ۑ�C�ڧ�*+.�F���
�|� �֤8�Lk��:�m�����rߋ���sn��v�����$������XB4�A��1[�nC�E�nְ=����P�Z����:R#����r�����t`ժ��
�"A+�N@H4�����^��x���#���O�&���Ē�F�wq�J��|&6�|���k�X�q8g�6Co~��ZbH�Yi�Ȳ">��ҜJ��)!&��6���7D�ղ.A�LÈ�!�z}=�|JE֑���@���ǽ"v��)Q�s��	�>=�C�2r�ɺ>)����4���{\Z���M��o ������L�%�maI�d2[,�r��T���^��ڥE;g q�V��n8�(��ל�3@ܳG5ĭ��)�C�6D�b�����i%�(�`�>�.�ʼbμ�Y	����h�5�.�5����ԟ�X5�/D�G�v��a����2�Yw���=P-�*k���F&7�"0sel�͇孁�	�Gcw|��(��u��ܜn"���d�uk��t?x`�5�60�G�_�z��H�P�Ϊ�x����q�u.�/�M�-�k��8,>�15z4,���K�/x4��[A��a�W�k_�P�yP�zw��#f�v[)������љ����;��fB��=�z=o��p�@{Dn^L[�yC��w�'O
������$�������T}T��/Ac#z��YԹ����QIm�u>����&���k����^hE��>Il^��1�Ay�Z�2z7)-���5�~�I����U�@�gMtgy;����N�����K 3���Z����헬�9�)C1�#�됞���7�P%痑�q���B��������lh��ؔ����M���M��~*yT��p�7�Ì��II)��Q+��f�dl�נj	m팵cJzR�ƶ���Ha���>�%��p	����C]���}IQ�ֈZ��l��1�ׇ���A�Xj��ь������\�<k���(�9a�OuT��;��*����2�y��&�E3�)��h�̮�Zf/dqi�-�W�-�*X!���X爜Uc�t׈V\z1�u��>"�EN��l�z(:����3�{����?v.��<*	f�C�D���M����v��s4�C�uY:�y��2�HP�y��	�&������������'�x�o��WA�5mƔK#�X8��u�M\_ה��>���H�h.A;Y(���sn�^�k!#�J���F����FՂ���-�%��D3�WY�2GB9ԭ��cB��d�rZ�i$��L��֋��R�:1�Ju#䧼FP���^� �h
X6�ѯ�X�M� ��1�Y�����6F�ءʁȫ��zc�l�&wח���ٿ��
����%��wMȷ{���hw83�苤&�զ��I1u}�a�[&�j=��PT
���h�Cʥ�є�- ��SOQG��>�C���O[��h���ۤo����C�G��f�֠�M�'���'�p�S�o��I�~w��.�Zc�b�4����#Dv�PR�%U2�@��!f�:�4[ԫjLqZ�_���*��ʡ:�YОg��#�w�@�R��8��]�p�i��'��#�*���#��N�F�Gq�$�f4of{a�$�Wȧ����s���0ߒJ�\�i�MqL�?�/u��n��GT��p&�Y�_A�B�Y�Ҧ����`�-Q'���9�0�"�)K�"�!�f�D���)����B�O*��>k�8��F��HE�U���7�z�KP	�q������2��Vx�n�XW]��fg�C��G�i�j�0F;X���
�i����@&�I��s��(�pd�T�UL��ܽPV�yө���$�4�rJ��w{ô�=M7��I�í-W�D��\{��~[r=L=i�Hk���A��&G�{�XBY�w��y�1������EAۄ���ԁ�*�f60b*���o6F���Ub 3I�>���G��.�4�t�s� L�G3�'Z��Q����"���/v�)�E�\J�D���o�%Hg��=+޲���B�p�wNA��E�(�ve�[(�,����I��,s�!#pvsbVj����}�����x�o;GBY�'���{�{��;���D>!��ͱt�� �KO�>#��-���8��V��7�������z����N=I�~e,C�M#��Ú��Bb�ó@n˯��i�Eɏ����������'S�Ph�o��?$��9�5dH2�����\�Uע�A1�ǽa�U��Uݞ3)#�� �s=��Ȧ&��J��4rFE��:�Y�IL2�$V?��b��{��5�~�\~?� �z��4�➠�L�vy%�d���*�#�)I��2����b�N��7|#�?��j����\��R �Ƨ���b�J��C��f���R໌ƶD��;e����c�Pv�M
T�k�#���H���`��&<P�9$(����aG����ϯ�Du�ױ���.�>���6I�.�����杼�P�(��O�F������rd$F&G�T.1�ڽ��F�A#,�s�J����Xp+,(LCV4�:��sx���Ee��r�Wڵ��Rc����4�ۺ�y��:j�C����e�I�P�m�sr��6���b?�7Ua�sI	U�c#��?/O�x���k�/I���F�[���P.S�T�E�5�c'�B;����'�ih!A^��Mf�&Y�
��4,��MD��d=�Q�C�����������Lv��2J�����at�b��qԘ�H�!�.YPi�3�o,6I���&�Wra�l�����d�vxD2�5��Vh��`Z��32?�}4v�d��Om�O���e�!��7���5/�$��{)_�;b<������>8�C���cEFD}��(!Z�_�����~� � ��A�8"����|D��a�.�
���o��H�Ϯ���ߌ��m��[��4��_���͗�ӈ@ +��@�����6��5)��A�t��u��o��W�yhf���]�d7 �i�k�$h�\ߘ��GGh93��^0�V�I�k����uyǇJ��aɈT�:��W���F��vM�i���
�� @������~�d�g�h�_�ձ�����b�_��8ڤ��{��P��O��)(��𪙘n�����A�����8!��=�/b�^����~󎯷d������yr岉��՞Ʀ�n��{�t��F�����P�`zbP�Q�v=�"�g��G-�j-�"��2�K�}2G��dg����j�c����<�!hpl���w�a��%#^�䇰=DC���q���멽G�B�)A���U���M�H����fT0�)��s�9�L�Ţ=�h�ݍB�ض�!��C��z��0 
]�3��Ǣ�JS>G0��h��X!j�旰��/҈��Ł�b@KlrjO�45�h�v�a=6�Y�U�MaW'^��'ŌyeeR�E�x$KIr�Z�d����\�6��ɷ	����f��g�%�C FJT�z|!�7-pW^�qn���8�϶jοyt��G�h�_��c�|ToJ�f��r���X�}*�H�3N�ֺ��q7���J$+n���� �<�"�|A�V�pk�@��_4��`���5/ȝ
����HȭXh�;w@R?��%Z&��l
�1w��UK���e	�:��� �UR�G���s��D�;k��ڸ�֋�e��O��aE�ͤ����\o��a�}c���z4B�(�_���!�iO�����V��K������M
���:�q�FX�����iH�&>���)y?"��d�4_���'���#�4���?S�tE��@��#J��@�i<�g}nVN��{
�N�W^J��&s����J��6�v��,���%7��:�i�<k��:���k�@Ԍ�,RF�E`Q�If7m�1�w��Y���4�MH�k'�2��d�Ũ��_���g\e��Lg��;�U������v�\�0%J.����漅�}�bxBB�_PFz�u���v�/��y1x�c��8m�����5H5��D+��$ٮ�_;�%�Of �O�˓��hC����-���~F����"�����^�%:�K0<���BΪ#@ke���N	��*�vT�x��+��U?T��Dn���c�N��Sͺ�ͱ�%1��Q�jؽ[G�
.%MؠHD�7�B^Å�̧Z ����0�K2���t�+�1�r8Is�m扉��M(e�~����}ï�Ɲ���L��s)���s���Qc��c�n�kc1^��ɼ(��gY�@�T�B���K�ds���Гþ����{�F�A���3ͽs-���Ϭ�۬t�b��k�u��f�}�Й'��&/����*a-�����ֵJ�b�.�˭����b�& �y�2�A��n��H59;vK�P�0�FO����:ht<.F��v[8���.Fr����;�#���_��p���YQ�$�%.��_�!l9Wa����x)o~� �[���RV�h�׿�/�JT��ݎ�Rd4j��,���U8#C#�hU�,��wLL*W��Zӡ�TPu�4(�l���1�wr����P�~�m��]d7�y�Ӵ�nO���2�	���=�&Pլf�����ER-�q*�W��9�3��Χr��pE;��[�/j7�F(7�Tk��VJ�Z@ X���3�T{)�P��4�_D��v

��e�eu�X��w���w�k�*N;�(q�I��J~*5E��fO>�����t�,Zu�5*� ����1[+��j��,4Q*�h�c�L"&N�������2��(/�ai�<�=T�J���#�����r���h8��P[��P��PD��ճu���j���¿S7�����¦y03�g��Dgn	2֘��Ă�H+q�@�ĉ{��tF��񺒮D�6*�h��5��0\�g��kǍ2�����G�A��]�-�����O5�Ju�����(���%y>��4���-1Y������[��h�9HaT̲�:��"�X��0�������q����B�9�z-�K���h�{�Y�x ^4���2�6�:5x��z��0�э���Ӣu~R�צ�X)�;υŜ���g��� '9%�\���_�F�~���G���q�F���ʐ�����3A1�)3%N�'_��wR*���T@�%El�'�K�dh�|ޝ��n9+Ku2�co9E|�q	��p�ǧ|*E�ՠU��[.�k#��ԕ�4��1ϕ�\��W�^��tG����[��w���دy���'�#>߹�`|�h9�b��;Yq&5��0ۮ�'fv���mrz��E8��Wƙ�^���'�U�XlZ�<�eIF���.�A$&����:�w'7�܍q/u�eO�ݘ����:��g��p|�����N�֣^(��l��p�rP���?��}��g���S}44y���Uj�C=m�O�r�>C	?�l��ÝA=X��:Y�/�u�3���n�2Qz�\.@o:�.g8�k�)Z^�O0�#��c��1;���T�+���7uU:��up68���t�'o���0��dI.֚�dy?�B�it
��a���⹩Q�yX���z8\��ҋ5�L( 6���"��	��[Ǌ]�|}�&! ���dk�.�r��Ƽ���ke1���gF
b���?��nu3>�Ŧ�5�l�c^�@���k���M7����7	����x:I�� �@���\b'���u�H��u�5ͬ�h�YćFys @�Ǜ*rȆ�&@��%��?��i�[��1���	�//<��Rx�	���*��]>��9�%6z��:B�ͭj�JB����YR��FA@���B����g�~�[y
�)��B�7\Y�ce�J?v�!���h$�^l�2V�MP�~:)['dE�LIg��������!�d_>�}!��o0��䏶1�B��V�&:�<���x�S�'S�ioO��2u]"d�o�'����h��ByQ��
�g�����\��jL���o�67Vܜ�Bg[��>��F���@�-�	��N��/PP�ߤ����Bng�zN�(��+��K=Iȇu.$�;�莁`�n$���$�C�(�v�F�t�๜W��e��)H1����^�ɸ����7��\q�t�>V,C]��(�KL3��3oJgz�ܵ��dd�Ib@�c͕�Z�@A!�����,4������hcdkq��z���A{
q4D�8O�Š~�4^2�[t���?m\��M�)(�m�$��i>i�����~%S* k�|��ռ� ���.T�BbC�
�M�R|� ��b@�Q�V��K��������s�8����RSq�_mse�h�B��vN�Vi�*"˸{���_���;���Z<�H�.9S�M�4&q���:��$�l��&*��ڲ f2G6�I���g�u�L�ƣ&�)�<31n�E"�/�ɭc��%��� H�Q��|�HT�>z�E���<2����ċ�l��R�[ gc����N+��.k��ua��h��_�Bĥ�I*�G��x9#Z@i]�>h%�rB̉�����'Ҩ�ώ3
@H(�nPQ��Y����M�[<��;��5Q�No�J;�cOI�97�@��y�msc+�P�Ă��Av=�-7R�k�ym9��tQp��9�E*�O76��b�����U��~���	�@H��Q�O]~����*K�S���M^����/!�54�.(,1r/J	Ꜿ[mF����\�oj�6T��K�����e�9�+A���5��]<~RX��
5C�N��B���]x��������WWj���.fU�����t���������KФU7Q���r���I1u>>=�R#�B�Os�����M�><S��D��`�8|�_:N;���%3Q�	Jd���Z�o3,�Ȥ�鿌�l���
F�[{
���*��vuwK"��ڿ&�S��&s3S��D�k�tA�	/fA����m��S���S���X]��$��+ySM�%���S��y�Ef4����}ؿ�I�
1� ]�x�.@�l��#7Wa�v��rW!S���f�[��LA��P�qd�=������6�;���]_� � =L� I���J��ˮw���;L��We�#Ӧ�Ƒk����U�!�:���:x�(��z|8��5�Nꤶi]Su32��Q{�]e����-�&�����͟�Ɨ�	�v]Rm��Yx�zjp�v��O�@�uO���UT�e&G�h7�ɪ�������P��h<8��$�P��]�0d��DZ�'f*.�eSY��#�v�`\$)��F6��j�&� ���Γ�&6��ꩭ��a��s��՗JE������?���� ; ���D"���(J���m�H־�}����C~����8��� �V���B�
<'xhX�����)ʃ+�"�U�vZ\ч�'���1%)�3X�L8[�͓?_J�A��9YA�k|�n%'+ܿ���b��I9�q1l�������k�$�����bG����Տ�q��s9�y�����;Xh*��C���T��R���a���6�8����&�$.�1��35�+&����Y�w�B�?d~��F9
�J���y.�A�/��''���
�� �W�q�{�Ju����mZ��1�����,�������4cۂ80�X��F��?I^��S�l��96�=�$-Z�� �����4���,�5�x[��f���ɧ��A����K��#��� ���ⱴ��S�������(.�yWOǳ�%T�xR��#��G}lu�_���l�(�b����KJP�Us���9F����Kq��¸�bR�m���l�=��H�9S�&l�m�r��?"F��N�q(�z3n�ɻ�Jክ3B�7|?��������88T���?L�p�����nc=]C�)R)�LW�cv���BO�zS��Ĥ��c��RNL] �h�<��Z��S]/�,�+�c��H��v>�x3��;������(���5�B2�M踌��m��򷴴��VJ�CN��FH��@��{xT�`�����ݑ��7֠>|4�]	�u̙M�ύz�X��`�]:�o�j�ww�_��	�����%P��1-`5Hۂ��sw�V�.iH�B6�C�W7/���??Q�?o)<\1ʨe8����L��Kz{���.r�?��86�M)�;q��L_;H���e�v�SL�H����)�����T����$x�N�(�hAr����A��x�y#Z��^�A�" ��T~�[s���9�@�n<�[�Q'��e/7A��R|HC�ڱ�b��W�G`SS'��m�|�]�b����&t��1Jb�8�����`<��L |֒�$o�\2�Y�����e1cͮz����݆?������-�^l�,m
�S ����>V�~aY�����9�M�v�{��qo���}��2�^1f8O̺t��z,�o9�L2a1��C3BY������[���6��b��U�̘.��}�1��%��ޒr��M����:��õ���ݩsňJ�Sb���t�:�s��S��)j�� iđXBV��h�h�T��!�8�C@KW㕘���6&���J����)���C�lwcz_-���Y�-&ױt�'��)�����o���������}\}��3�"O��	��l��ރ�f�w)jq�r�_uq���N3��
 �
�{���� o��|}�3 ���Q<�LR�x ���'��@��5��x{2�葉�ˉ�;��AU&����Ϙ!<�������: ��8ձ=f`^c�m%b�&|�S��Iδ^o��̽G�v¾��s�A�!	�J8ę~�@��k�_.4��v��Nv��ޜ��� ˫��Ԅa]�3�lH�)p��,?o����n��PJ�#�ij� !���vE�O���g)�Գv��Ѽ�Q&����ȩ�qt�$C��s�t�
py:��#ϖ߰_�P�� a�Kq��S��ppjGp�Kz��Ȧ���^3�%��돶�gz��{�v×6_V�3�cr4;�@;��H������g���޷œ��ѺޝoA��3>8��/�^JA q�x|۩u�Q���8$[ͅ���-�bǕF�-׽81ǀ�]z�?w�
ٚ2uj�nN_������G�hp ��V�i��`�&PM'�:�M����镯s��d�X���G�
��A�i Y����[�ZܧCq͙|?i+����������m���3�'ɰy��Cq��A8ћ�[��p�`���F�8��')���M��9�k(����3�NQ�קĕ2Ξ�Z0t��7�ا��������[�5�:#��fNB^��k[� WÏf�)�H����=��dh��n[L�.E%?P��Xil(�����M��z�����2��H�ۂk��Cs�kI��ğ�!��a�4�ҿ�M�� 7�̊�a�$y�N�b("�#�3����](��t���\�K{%ք�[ ��>�9^	��VUU�5Q��c�g*����G��&�x*���nY(<'j�<������>̆���t&%jO�o=��T��f�H{�^E�ğ/}�z�I��Xcp����#w�/DJ�@�(��V�lmҁ��ܡ��
�M�3��e�QJ}P� 3lb?�+N����}�E^�8d����cm�t(\�a������}���;�)fz���'�����"'J�KWΛ��Ř\�Am
_s�kh���W�M��uz�]Uk~-�.��En��{ŝ�u;r7��1���E"�:���|�W;K�hI�c��zh�i�C
G�^DsG��*]�RUIl�Č=| �E���~�o_���|��3��1���Ry���3b���&j�ͨU�)��r�>c�șn�E3���WzZ�7���T�t��������͑�s��Ʈ`�:\s}����-0_v���� �2+� ep؜T4'[�9r��_�N1PPK�V&z	�jV�r2-��Ft������m������	�dZX�!L�]r�!�����!�Uߌ�u��)��B�R�]�"�yZ9�ۜh�`E��x2����?�����	G{����= b�ѕ|0�*��n���x�$����1� �Ͷ�|߉�.����6����Kŝ"m��f���+�v{��^��<8��ϳ[I##Ɨ�Z�)n47��t��>�+�֥��S�=H����1 k���+�f���Z_̍�y��N2��J���^�Gy�Z����}{P2/�s2W��{N��3�A���5�`K�XU����%G.��x4Vǃ�'�x�և^�$o:DE�a�5Tf�W��8�t�C��▾a���uE����vTk`z��e��/h���L��]���J6���� M&%����袢������lT ��x;G��(R�)���'Z+�Uh��"u�>��튕A��SNDލ #���Ƴ��C+����F�gū�i��d$���ȇ�5i����s;�B>���j}��>]R��9ދ+s�	�=�w0ڇ@�<��m�֖
9�M�;1�?�iwPU�6��2�3@{�*3��7��u�c�����ꌬ7܉�b�=}#���i��]my�;A��
�GG�/u��n�+3g�g2sX�F��5�y�BW�P�`�9��T��`�q9Jd�Y㫋Bt�?�R)6�� &�j��K��#��}�~������ߋ"���7R\����1���;��v���1��}!�"��..��3�;!Z� f@n���c�c&�����6�h�X����N���6��Q;V�H��{��Tg��zy�V����s����u��'iH�ȣr�4�uS�ٖ�3ED�j3��i��@!�C��HI����ZF�=�B�Y��J-'W.'k��:�.A��w�QapY�x;8>��iWI���2�P��:�&�-@�u�FWZxv�>�F<ƥ�f�U$�xƚ9��ʴ�����+:D��@\������LTb�I��f����M�@�������{j�c�k�����7�ɗu�/x��냈iC$u�*��}�|;��L8H��T����M��~�Ӕ�,p_�}��]d���^����&w��v��@	:�C��t�T�*�HJڈ��}i�L- f�ܔR�ku�d3�k&XCZ�%n��cA��P�}�����L������n��eT��؄�����)�E����G��,�!c;Z��~��|�?�`u2�z-d�zT���B���eym�K}����6��u�� A���vt
`�������J���!�I���$x���|���1���>p��
�Z�m���BSlK��Β�872}���A|���u����x�m�b?(��-�)�Z����թ����W(�.�te�R��C-&UwN�8+�W*��:���'S����Sa;	�Y�|�[��p�ȧ��J�f0�U�Χ�BNn�m��Х��Z��ŗ��.)�m�|��@��T�r�lS~��s����=׳ߐ�5�ȶ�E�am�b&S���a�;_�#�tx��DYG%g���L+�	k(C(rƧ覷tޅ��׫]t~�Ȱ�I/n�O�
J�!��S�<�����N����I@)�V�1g���OkzB�`��ay�C_�|��pw�n\%��m߮lvL�i۾��e��6�@ꗋ�U�lf�*H�xr�!bH���'�U�\YቍTSw�Ϫ���d.C����܆�����X��a�4h���Tne��� ����̷gs�N�_�[��DG%�� e��:� 8���~�����k^��c.@;���v�j�5~��5t����2>�6�"Q[Y/r��%�M��H�]Y]ٷ�H#����k�<H�Yz�=�m��ɸ}r}p�L�Ņ��rѯ�V����P����b���9��sN�,��~���r�e�b�N���@���pb����dsߣX,�����@j�Փ�Y�a5u��WC�ڕ<��a��#Uv�l�������VD���t����/[�ܸ��0J�B��1b[P���9��Bjտ�g+!%�� ��Ѽ�W5Q�J �Ҵ*����0Z�+j�ȗ��, �xnN7���dh���	x#р��XR����ϋ8�����!��l���Ë�g��4�b=��[@�ݜ�_M�)�l�/'+!�p~l��E�_�9JZ�����]�.�s0����($8��*���̆9h-������Eg����ѱ_�������3&���=Q�P�hփM=�6��6 bؔ���w ..��.��jzE�I���7&��S�~�����p���Uj4�"ٱN�Xc���@ej�|g�s���9QMR�5���=<���`�`\��	��� �`���i$Y�.�͵-z ����$���؝���W��;k�(��s�3�Z'c?!�-T�#Ț�߂�2o#��r���A�LpVYv~DC�9�U~3aʐ"7� �r���复�c�\(�w�����/>�Ln)C��
αS���d��/�`��dA��%t���� ��,�f��'�GZ'O�1���G�_JW=���^��ɕ��PǱ���$�Kf�e��5��5D�w��(ȗ�aB%n�[��:�*ئ�N�T{@Y���ֲ����i��^��ps"�]�i�J�p\oǼ".�1$�)���@ҧj��<�ʍ�U��m���#���ث�c�����y+P���, �����3�˨�~m��ݲ�3��jn�67ڢ�k�*�XS���a�6�/`�=�`}Z�Vͭ��O�=��M�=ó№�͞�<%B�)�d}��Ln͒\c�4Ơ,k��������?�ǖ'VY�1���c�n2p�Np5�Ls7�}���LIU�av?�K���y�:E�Pv�^�nt[�#��s�ͬqf��z��/f0��C�D�Ł�t��|)�m">\����Ū�G�����Z��F�K������G�D���W>AjV�����f��?��pZS��[�VJ�_����c�Gb;�Sݽ]>�%�}��I����G՞4��E�X��;�7϶p�!�_:�{�'[�85-�������4I��&�B����:L�� /����	�G��<{�u��:����IG@^�H�3}ݓ�Hbps��J.^�Y��_QD�Ѹ�R|	��Qm�9cZҟļa��nft��@6S��hD�o�wVs>�|�	z�1��x�����7��~��+���{2����L��A�*V"{�EX��ρgg���5)	^Cn��.��u�P�U��Y�g9�;V�K/ߡ/Z/�'�y%���1qE�O�!>�hf��7zqƚ�#�w6����Z[�mx�b�}׺(�r��sv��0)����T��V���YU��ޣ{���� ��C�r@���u&Z7�Q��g����p�m�� ����@!���ԙWNH�b��QYڡy�a��;c��z��;<P=b�Y���?jM�J�i��#�WYof�����5�.�p���2W(Φ֪�ƒ޶��	z��F{g��%.>|x�"u&3'�0�^�a^^��cn�w����a�������.��s��+?]|1R��`W�ӂ�H�;�]�w
�.�Zβ`����Y�!yp�hv��
��"6]��:�������zB����`KCmhSݐ=�@c�)o�����\lb��xﺉC�N��h*����I�����/����)lĸ	
=4Et}���$�j �7��l��t9�'h�>cc�ku��b��/�o��'�R�P7Y��7Rѹ4f�6Jw�9ꞎ�	�WKw؟!�Id.$��55��=F�wK�t��6_u�~�����X�ٻ��s^F;:�!�x���11�t>��Y��2��oݠ�ہ�Y�a����q"5A4Vd�W,:���î���M��9���!2�ι!���J{�՟�y�Ovݻ�C�JBf��I����QX	�0�����A�l倠*O%�=���'$:-�Q���t��}]HTf0�������E�*��� c�,�.S���c���#�1�#�C�:�$���}��겻�K9�����5�$�[pە�ϯ`�:��m^ٍơJ)0��\U;��h�HHP�͹���JEL?�7�*�O�'�r��j����S���ZK7XVRM�S�Tu��Y�����V
��T��<=�m��t8tO��H7ΫU��hlh�ޝ3�������R������>@��ֆ7�}�g�>��W��ꥧj�%~i���WǓ#<�C�1����#��Q��č�"�à<�B]����l�59C�Y��O<��tqX��ʗ�O�7i��ʺ 	�`�}Q��-�+�B|��e���
��#\4�h�\�65���mCa�8���rj9��N��ocȯ5�!���Z������$1ƀHO�aÁ(������1��=o�GYQ�0�������Z��>����ԫ�3hf� �A@�����t��ĩ�i����G����D��=D�H��@��'�ёL�1��|�6�X\�&�(e�O��/�w$�lb-������_cE���N⟾mDy��Gd�=hb��FW�yd�d��W����K{sϴwÇp�<д?3"��_]e�d۱����m��8|��8�
��d��L�u�3B�������ٚ�Ҽ� ʹ���^��0�-�u=�y��0�˻�J:߳�聇Td����@�gl�M�����س̄�g��S�X�
��8Q��&"v� ��K������QQz�7m�T����A��w�cq	2���0�ex|q�Ro!1���:wv��`�Q3l:\�k��㐤�.$�T�� �j�y[�A�����Se_P��jl~"t_�Kl̍��&�bXX�> � �����51I��"s|"���y���ѐ� R0GR�N�g9Cv����[�b�hD�Vn"�-:���s�%��ѩ����G˻p7c������m�c� �V"�.X?��L�y�#�\r����\����S~��	9ř}鐂?N�c")�ӫ5�J+�D �n|��Xv��,t��3��6�}uM��x��i!ҹWF
,�&��y5˧���A"�ʮ\�Y$
����S��3o�=E�7.��X��ϕ˻����g?<�}�e��Y�%
g�x����]t|�����ku�	�`�u)��q�OņC����s���0��b/U��T{yb2Z?�[���O�D�e����7Ti�������Q��S�of�sFQ���}M�t�P
;�Ʋ`�7tm��D1��M�tE�S�1/����r�� ��T}FM����`q�����JfVG���ٔ��3*�|��X(^'��q$	ޏ/�Ǚ@�%��󝵟 �\�5*�^v��a�����>8����6�N.mhE����#����Vq7�y����癵nK��ސ�Y���Q9��ߟ�>cz��<l���G�n,�EI� �B@�[꽥#}~1yf�{�>�Z�N�`���~�4&�F�r�Z£��ͫ!O��M���zYg��9^*���M���jo�� �i/cz�r� i���v�me|��?q���8)���$t���Ȣnڗ5��/����V59�Z^�rD����p��ޚ��n�V�8qc�S.@�!e�)�`���"[�%������pB��_4��]�d����4� �7����X��cm&A}T��,�-�"��m?�B�Sq�Ƶ���4rl/Eӎ�G��R!ϔe�/�T$�HQ������S�����6������q��r*��(��oƂv�q97t!B�UޑL��P(
�3��`� ��5�:�Y����%%/GUf-���Ч�UL�6v3CO#]�D�Ħ��S��$�>�����X��@� �q�C�CJ�F���o���#�%�����49�~:u�I�i����TmM���������Ǥ�\�͒f�JlV�y�e��.���=�9=���|),}��m�FgE���ڮ$����_SuD7�1f%M3�4�z�A� f�гj��]��Bv<���_�3]&%�r�=˖}�Yh�ޗ+x��ۥ|`.�b2>�*����Yp���wD�U���/���[�*]�瑏bs�߁{�h���j��a�C�A%�n��j�[ ��l;�e���P;#��P���6K�2�L�ȟ����V$H�����Si.��B�Rh��Q��o�+/Q���'r�J���XI�+�$�o)񃠿�Vj#��sY���q�,���t�g�;��_��1��ŏK]���\'Q�_� +�L&	�y�t�����r�Vz{�{��������yM?V���r��
��GK��2�)���|���X�`i|Z֦�z����""H��
(��~�x�=���7���K�V���@Ԓˎ]�; X�L�O�����ч-��4�uJB��o�P�gU֌A��'%��)�H���@� C��n\��R����㉆d��C�� @N{=va��Pl�Zg�J�M�E�qg���\�.��zj7̻}R;,�?�
d�n#xx�77?��Z�ϲo�$�-�ѕڣG#8}
��K��=^��	�p����N�4 ��s�l�ӥ\�_�կ@=@8+�d�Ra��&�����
�1�7RO��G��nr�h��B{��ed��2b o�������#�y]�w&O�J@���HTrܟ>B���@�v�l#2ڝD�%�cO/��`%�vz��4)X�iH�3[_Ñ΃%f�P�H�8bH��.ee�/�������І	5	�.�1�*/��߰;D�y��tJ��S����R����9����沊`|	5��`�:q������M�m?��n�h�6whL���.kՄ1�Y��e �o�qQa�Ώ��ژL���4�sgt�>�6ӉRo|k��A�دƉ���^����}Nc����:C�W��P0���8nѱ$�KHv���@�b������~� <�Ć��7�����>fه:� !B��-2wxjԯ0�>y/��}Z5���5�V�4M�x{�g��M\SMʹv�����Y�1P��]��[y�����ӻ������BIe��X0qt!Z�)KY/�U���0M��������?�	��+��T�r�t�J���Ԟ�r�u�@�G�,Y��z̡��b6h�-�2�-I��]4�����c�Ï���{�F��o��
@����n�f�ߧ_�����?�{�H�6��蟜����������aݎ�������'�!tc���Qݴs\x�wT�.���H����a���e�r�n������X��ԗ@&P��L��?�0&b&��EG�k--���;g\՗$l�\�Հu�J�+$���7$j=#��FiO�7W��B_�P��=w�G����6�MG�xt�v�Bޘd��qo� )��y���"�@]��{�u��db�o�r^|i�r旘Rg�n	L�Ƚ����6X����c�z�����CV��H\�Jqm���μ���xN�`�/2h�}v����!����3H��Ol�ze�i�Y8<Z�y#��$��{����0;�����
^�Š��\'L�k�f��=
;1�52*�����R�)3r緬�4`���VQ�P��΃� {���R����xƔ%�q(r�2�3	g��	�.�ӹNyݚ�@�[�1~����O�`�'(F������7d�ʞ��{ ������-��x���`�Nb���Q�v"�H7���v�$S/�CfuEJʒ��$����su{;y�>��RL��$U�6�V���{�����.�@QQt[�=)ry5!>�ԭ���dw��kMћ�;åWX�s��z��d,p�(���C���-�c����`�C��ז&�ɋ#aA!��rHb?d�Y��me��O]����c^>C'�P�^�K�	�Jg��+6V����P��%ԵY�K���������.� ��c��a�ϔ�bv,�^���g7���}�鎿Kn�w�fL��*N�%YZ�#Ɛh�ڛ0�"�pJט�o��@�l쒍�1+cJ�F�>~��5�d����7?,7t��@�=��c�TEk���R�HW6���@�$v����F}�@c�Ĳt���\�9�F\�O߈_���E��c�.���#Z H90C mq�-�*#�]���-3��/�.W/]-^�+�QI�GH!Ny����-',�^D��u� �����Im�J�8�6���gw�	y����e
2����/�F�ֱ���(א�t͕5&u��d�`mj�>?I�Wlmߦ��יY� --���p�_����#�]c���L&�U��2v;�{��n����j�Vg�Ĺ�E}�[�x�����宽�ĸp~�wj�`M!'9v�%���Wq��
5��L�� �;!&WB��������I�X�����E�[�I ��}+kg�S�%�OKxk��=e�l0��� i�.|X[��<5�A����3���_A"�v�i�d�Ǜ�ɺl��j�d�J%�𨧝�Nat2,f��v�ǥ��cѺi�0�P���H�{L+
IZ�U��._�7��p�����(���dt x�MTk���/Vi\�V�l-y��1�'#
"9�ӓ�7ݹ��&���Y��[�Y�b�����b=��'lvˡB��ߌ��!Y�DހQX+�ulf,��y����)��fB
����|��]W���G�����u@�r��}S#�
{�>P��߈i�X������H H�t�{���3�2Zcn�J�}�'ꦁly*��C�k����}�5����d߇8G�����W��
��=��֨~c��)��햕�-��UF��+�������|o��������Ƕ�i
�8�S27�����j�0u��*�nR�*m��L� <kӞssR��pڄ�M��W&߰)��{فg�I����U�!�5_"(�K���P���"􇚆��A9�1��'�ޓ�_�ę���zs^�B��(P����z9�4��Y �v3�%S��z��TSO�ާ�}xnc���z�z���	9 ������= A��t�U�rb�f�-}��Rl��g:�?)A�S�ܢЫ6���C��m}�QX�s/'����V>l���7.��r�B�%� {a����\���7_�y��!�V��)��-L��V�
6�ѱ����[�S��!�~^�X?���vˏ��!eq2��YP<j�|Rv�Læ�9�\r�K�t)eZ�����N?OF&�hN���`����}��ܷ�}��}��S�s8C�:n9X�x��B���O����ݧv�mqN�Ui�g):��2Z�ŚQ;=�d2�ۉ��/l>(-�BM#ċ<���{��I�,]ڹ�!��Q[��y�(ixg��ِ�6 ��]_4%��q0A�y̎w4�~����-�䀆�Qx���P����i�)a{b��kYM��.��[�}�2�g�s�[�
�ی~z�@C���|��SX��[އ�]�y>��pu�����	���_�F7i���i^��CDh�P�ez����%�D��6��d������Gf�����oZ�-b�B-�4K�8$tY_.�_Siw_J���X�n% ��Q^4�#��֦�f�qPX���$HAs�����&[CiQ������E�u�A���3�]��PU��v���g���k��O%zb���6�����2R"hXx�Fe�e�'��C��I���)�v >�����ZB�QjA=n�!<qׂ�m^Vkn��xy�nye��9o�����,ϰg=t�kLO%P.؃a�H�v �-�g�'�CR��?+P^

�/�Z��PL��w�i������i0���!sٽ��k�6a��-��ג�B�Y����x���#�\Rz����A���젻
'*��Y�XZ�&�F>�����R��A����{j�����l�	^�:^�4�z�'�[��\��EPҪ���µ~�Dq]�Y��rW�]�ӕ";@��q�[v��Б���������54�CZ�K&#�n�f�9���u��ۮ��>�I����5��sɨ��`�9oyb".EƔ!��@Q� ���� �s�M&S؁@LHu���Ψ��\�H��R貄�@"�;K�8T�^�֪湥"�J�}Y�.��$�q�m����t��x?5ь�j�ϏX3��Y.�����Y�u\��Kg�<���y�3�r��2��b�&��s�|zUUk�)�=;H�ä�*���j�#�\�9�����y�Nqk?�"X�/��� ꎏ���S��3�S�g2�y��_����<{�T'y��,A��ږH��f_�������5��7t�b����j�P�܇}b��p쑋	�B��P.����Wa��fo<���d��)Y���}�Lh����Zz

�6�gkب�K��V�'��Edុ��	��#M��(L;G����Q}���>f"����@h�;�Q���^�����98q�⸉���"��:*��A��P�:J���ʧ�}��ҵ��(`�7��ﴹml�5��֭�s*.��u�  �⁏�x&hSt���,��?��Q�X<rX޽������*�})h�����~����8h:���
����Qm�̥D��/~�}�Y�V�Vç,d)0����C`aL�)��SmsZ"T��Rх���w���l5vn��\Q~�r@8�"3?��[�&������?nv��6]Ԣ"����8>�Jba���x�i�-��73�κ�>ۈ�8;A��$��Tz�;��o����"U�ޓ�����o�����qh�00��m�V8����v���m3,��&1�i1��L�#��6Fׇ�[�wa�g�ºX����o��:Bj��K?�a��V"O3��X���}nJJ��{ZuN�uڏK�<���ϕBǡC����rDС�E�ϙg>�l1�Z5���տ�˦��`�MHK���`��	���i���Sׂ�i@+h��,[��V��Zh�Z�X�4���(@�[�_E�tY؊7��y%y��ܐ��a�S�EXB�,�Ry_�>[k�M�$F���T�c�E�dO* ͬa5���m�1ID��t�-�T�*����ݷ�w9��7A�Ų�8G��R�W�z�/[Lӯ�@�+����4C��	�j-m+;�9�7n�O�����ۭ"�ڑ��c�2�&'����A�vN!t����+Bꐉ�3��<�Ս��n�,]�5��*L{�
�&�X��A��ʛB��;�m1��*NC�0;�.=e!h���iz�Y{riB����Z+~�.V�(I(h���jRey�����۬�X��`��j���쎧��_���hJ�����~��hN��G����!*�ڵ��[uر�1���6�_�2m���T�z0��Zmj��Pa���GE�FK9հ�t�3,e{�ص�I�+�"��DqT�]�:�`U'µ�M^r=�CɥdO)q,P�Qk�D^D�B��y�ɻT"�,f���ra��Jr��Q.%�	���>���	/g{vk�ثJ��;��l*��$[l9q[ _�Dƹë��YL�	/�X�9m?d�kI�"[6��I=���$똎�*��1�������$��}PmT�����WsiEZ'y���.�lO|�3�Nf��K+�U�|&��x�z���V#㾎����5,��L+	a)'BN�h&�0 ���g��*�����b(���c������@�c�3��ݪ���k�}�����s����T>m���/@-SbR��:�<�E�ߞ����K�e^eq����S����Q��l޴���ѱ���n���w��b5��	>{�ʲD�G"r^D��I���r��!�A����(�Z �_�=�_�A|_-��_��Ӄ�=J����ۤ;Sb��>���BG�&&Ac,�/f�У]�
��9��-���f?���� F����I�o�;����rk&�)���~H�-��zF�\Z���0��MY8Fϒ��w�D����W��PG����hq�lr�2�f
T��HOE�H6�� ����PD�����:&�*"����W��,�Hk'K��˖�F��T�y[�߻uT�շ6&�8
 SiIuG�v�^i_g��_'&ґ6�̛���k�t��NJQ����!���"J�+�-s�y)������鍘rJj�P���,��D�m�?+�:t� j��e�R[��%VPy�9�%Ę�P� �i/ڻ������/�;�\C"ӻ���	��3��'�"�_ug�,��xa����)����1��<�����~6/N�c�Eb)C�ir��	�XY����h#0����B�X�<pY%,WB��]��vR�J�B���	{�Wdګ�<�C����&x�M�o)uz�
M��ѧc��q��F���B��XKX,����
�xܛȦ
�^ɶ�(����92_y90��cN��&��1�7���:�7�O�D�*��Z�grs��Ժ�K�<�����ך4���㓘�������'_/G�g�3���9/�o`|e��M��B���Љ����(���Z���@�HQ��]���E�~6Ӻ���$�kd����J����? L
���J�GAЙ�$�>0�F����o:	�-�>����#"����A:?�b&��{�E�א�3��)#(Z����0�1���\�l�C&��r�&K��Lkawuf}2j\S��c"ɣ��O_��V���~�]�>S�\U��;��I����D-��v���'r���l:9�\�P)�T���Ru��h��"7��?��5�B��J'�x6���3��Ǘ��>�WpTip��*�n��T�,���՟)v�g�lJ�U|�:�1Z�oo*
���ᦫ�8�'Z�j�ۑ���P�
���X�!���>�o6�iMH�&.���@��]�62��&�+���w9�����Iɸ֊����W�`�(�ÕVt��� �_ ��}k����;���UQf�ԾJ��0+Kԙ-e*W�FXTL/*q�w���O�t���9�`N�$�][
�c<dEғ-hWp��?b���J����jԎ�QҹC�'k&1���P��s+��6H�Z�t!�:�1����$��a=���j�ؐ���i�J�.s��o�y�	S��o�U�m1g�t�R���2l�P�>O���(nU䮀�Dwa�|)㢽��-_�ULl�$��{f@*�*Z�$�S��j� ��j�=�ğ��퉏�Ϻ�iN�Yk��4)��t��x��A�C���/�v� �<�\����O<Y��e��г{0�h]n�h��!ZJe82FJdnUp�ϟ�'D�#����6��2��2b�O��}�t�*0��#?Ԯh'k�]Ƙ
U�O�����^0���ܞ���ٹ�췓�U�{I���_����9�e�!	��QW�L�At�>��E֊�����d����~��8�΢k�����8
k}Vz��9+�)��T���* � ~:4���_��1	�.��	�,�Z}o��!Z����-[/��f��6����9¨���N�Mi�)1]rRe@��	���C:�6ZZ��K��ABGg�S��sq� ��c�]�DZ� J��6Y�g�eEyV�_�;4]�лi�A���CK��)�D�G���ѥ	�(�vl3n^�8��Fa7֫=0�����'��_��Y6��� �����G�K~�dabkޙ���Q`�@a}�����>=y"�*�=����C/�<����9ߢK���3J����o���L�\���n������������+t%�l�Q֩����8g���� �x$�ic( s�$�9t�pC��-PƈR�W�8n�	��
�*�Q��,G�
��>��J���%,��RQs�Ѐ�;+�\���]��j�χMt���f�_P��Кi��mp�V���D@孇~���
:i+�*	��Nz2��T��z��0��<P�wI��t�e�/j�a'o���9�ت@7p�D}�I֍o�T�K�e�|��%0
����s����]K'�DXT�(�k�T�;M�J�x>�g�-woe��:l��N�%��q�&Ůxd��}�~S�^�o�y�
-H�E�t:Ʋ� iE���x�y3��鲲yU�~��:�c��m5a��=^�P �6�Ј���F]#�pֆDS�¨1ދ�l�(c�� �5�ܷ�dq��A
(��a��h���T]�wi�?ݱ���4qϴ3f{C�h!Y&����6�F��f��1�*č��Y�?aڛ���LF<s��w�BN����������=vfe��ۇ*�bO��0�O�	�JEhr���:kO�pOk��"b� M��r��tV�<��v���Y�3�+��p�(�%�S�a��@��Z����A�On�O�}�O�h=��,\��Ġ��b�3�@udǵ|�p*涾^i&���ۗأ�RF
��
�L����7��ܑ�y�@���>؎A��Z����_9����18�q��K��O���ʐ�w��S��w�')�ތ�M��VtҺ�(���Y��ҩ�2���[ \���V�����R��(.�����e�/h3���5�d�w��� �{"�b�5�� �sN�UQ`�Z�H�����2����
�� �c�@��h�9����q^�Z�Ma���x��L��!T\�T�v���U���4U�N]��A� ���!�M"އ����W)���"�݂���:�6���W|B�t@�DL�Q`<��f@̩��SoV�`v)�#�{:�E Y�^���g���юx�P�#LC2O	���ʪ���1ir �����) D�g6�b�IΜzs�H�M�J"a!O���g�"�6������T�����g,x6?��6-lc�' ���!�����T�7�ʗq5-�����lХx�1�a��2�{,)%C?)���ߙ�� x�M�g�����`�8�,)�(�kG��ǟ`��A�,ߐ���VR'3��(,P����Յ+��aƞ�t��s���>�"�\׫�8��=�D�"�,O.=�ʾUw���ޥ��bs�Ku$��"��X	 |x凧�!Y��]j/"���3A2��p���c�BzEjr�A�[f]�P��|�[�激ܽ�q�f�%���SMKAQF��J���)̉&�x�c��9��0w�����L���2A��hχ�L׷;0@M$�����SV�R�����gf;��n
k����O�J��(�ݟ�Ɯp�>�n5S��7��*�5~�U��8���*m�^(2��T�v��r�B�Zdv��8T,���=�eg�'AX�xF=���cA�k|唩�J�ć��4��f|W�r��X/(�h���Twe�p���m�*��v�PH|�'����<�#��m&ўkH�B� �B�Yak[����C0L���E�JK�Zh���C�D4�����LD=�
R���v.C�,�Pޙ6H_i};���%�FJ��Cu9��P����."���S�!�I.2V���7�q��yx&Amv�Y�:��x�p���ؼm�x�{��S��2��x����+��`^$�������eOC��I���M�'ߛ��d���Յ ���d�����@T ���^ߣG�����k>��WS6	 �d���&z)y  ��a�0���7��G}��y��쾉 ���O~��	�@�^D8� ��ó�%��g��٦��9c�鍀rrү������d�8��������#���ܶ�{���E�o����!�C\�@F?�{8�>�]C�fk��0�/�f����C�%(AA���^PA�Ug���k�HZV�j�CH&j[��ˤ�f�J�� 3�GY� �M��>��=w/{�e����)X6!6������{�Bb�.��l䀿
%oJ����U�x��aA�xw��Y�Yc��X�Vq��kV$@���u��2**���D���Z�����t�����26s��W���Rd�ޥ��f�n�[�	o�Plt�,���1���T�D� ܅��r*J�R�ŏEݦM+i$z����:�G��Q�5P�i���\!,�}�O���H��/��yÝ4�C�Y�a��E9��\�����I�C%�����Vk���y�G�q���W�r��{�r�LN�u�Lm�L�_���������a���O;!���{�C���ں"�� �L|}��ӱ��}v��/�]�M�Jo�b�n�)�ի�qٕYl���5�����)q��� O�.󟾷앗���!۷�f˂��v�JH%�} 1F�i��v��E�K�m@���������c�s���F��,�-�{��U����\�,��.���Z�sb 's�a��oSS��u_!��c�
`��s�J}Ruo��49V�c����:�k]��VQ���	����V�%1���i,�+��=>��f���$��/��J�T�{���51k�X��|i���$DL^o�0e7��~�b5��}��L���ks5=�X6g������i#l�Ar*tXeǞZ�s�]��o�|B�X��J/���"��	�u�&N88f>� Y �$��"4�;�Z���z�E7t��e�*8��q�g�;�P�t�2r.�S���,4(.�GE�?bfPb�F��-�~c��ӇC�-�v@�#���oa��[���kJ(�o�R�TN�^i�h��O��B�2.�T��)���*�mI�E��k����:^2��#*]kz�&@�_�H&tGD��J���u�M�Z˳���1����F�X:98��'lO��3s��:�P2�������Uv��=^��`�nG˝��C��g�>�k��jE���e�ZH I�0�˭���z�ͯB+C�����Z�}���:�����6���� }�zl�����k�$#4x�,��=��%��9u�� �\��U����v��kOZIK�p�*�[A{x �]��QIfs1#u��Dѕ2��@`x+q��F{Nփqt�'�k�!��4Q��_�d7���%n�X��"���Hwj�윌�>��LQ��K��z�Q.��D���R���f��+�1۳g~���o%ړ���Q��b��z˄Z�����Uu��J����n>�-��䩎-?�_�#��-��nS�v����!8�Z
W��h�/���i��Ǹ�a��tI]J�{P5X��\����Ag��H!2����!���v/�0�x(�7q {��c������rO�Qз��ꛫVG>���2�_�`��A46�E�ê{�%%�ĸ����-'����^��a �["Õ��֙�&���L)�4�ߵ�G��0;���^?(���Ҁ!�Rm1sjeeCS?e��_��m*��?|�c0���0n^3h�"�3�mm��a���49@/�u�᱀�?WK��Gߨ�����6쀡�I�����_A{ZV7oy�q8��7c2�%��'�aݢ�6C�%e��1�D1ab���[���v�����d�s�5#㣥x^�ۙ�pbb!.k���lӰ�סT.�ԥ�2�sdg�v��r��WT ���k�H�	�B*�O�EH�/����K!
gO�2���:�/u��<ao�kz��r�6�wY);�wG��!�E9%lĕ��Z���{3:(ȡ|Vda~�]�Vw��-�ʚg��e��n"=0��l�rv�h,-��%"�^=j}�Ύ�u�l=���=���v'�07w~�����`�N���1�M-��H�K�ʕ��&)�`�}���/��/��4?�Ϩ#����˴O��.Ǧ�h�m�;��	҂�dx�K���ygKT��؄�S�o�}�`���C}�]W}|��
�d������'-�2g��D� y�TǁJ��p�_��;�ƹ��$@��
L.�z�B}ɧ����������Vvu��9���Щ3c#|�AL���C�=%^A����Ӧ��'�:V��-;jW�s��� �p�Q�!�D_��8�5n��U�T����#��E}?\�Ш�W�Y:��jpd-wn�>*���.��kA�'����a	[�8�Vo��x��w�=	��"#�[�،���\8�N��K��8~8ϣّ��]-(D�.>q�?7H,�ˊ�_�~��������@DL����!��J�;��O[���w��OQ�:+���8� ����6���>�9#
x����r,*�ՠAdN7��s8*���� �1�+�?Ё�Ǒ�Hv�t�=��u�%�6-�/xx�N�D����@!}�l�EI���B#��ķ��W"i�O��-:Ea�V�UYpZ�b"��|T券��A�΋ԡ��	�Nws�6��J�A������t���q־دIH�5��Q�3�TL�rU� �q��N����zs�*��AO��b0@Do�*b��ZE�9�?����΍�*��j��s�y��/�+9��Jy��e�k��`�!n�����!�5���DF�<���q
J���<��+'��9�S낺8��ET�L�'��E�W��~K��cHh�[+��Y��;���R�"��t��T�X���$o�ND%�H��n�_4��z�߿WW̾�L	��	�3��bT��v)�������P��e;��x!Q���?ͣ�mƄ
�s���^��k��<��W�/�"Ha3k���X������R�7i�Ji�?ޑ�2'(��>��0F�Sw�u�!��F�i*m�q���\Rw����S�WĚ��ұ*�t���(.u��N��:%�@@p�7�k>lӞ.s��VJ9f��p��+���/��(6J�g�׊�ى�E�z���t�2�<�l��k���ZS�Hj�N��QqeBw;(�?6I���`�A1LK��\�c����QB5����i��}}Ȏ@7���Qe��r�M����xJ�'���g��{�e3c���ͪ�h�cB�zW�dm��j	}��GG�=�7 ]n ='�PT*�UJb��4�j5�35ޚ5v\���)��Y�>���mh�Nj��#@���F�W�!���)̔7�75�ܳ�%}�tA��ݶ����1Kܩ_�Y��G��#
�'�?R9�A�f�77���Yƃ�}ct1p.�cw@<��Ք-�k�7Τ���b��ݤ������]P˞]�F��#����3h?���3R+a�Ճk�!q�C�)�Dn�nY��n�����1O��6�_�a�P4�H�t�K�"����,��/�ywCu����ୱ�䣹�r)p �OC��ii�0�a_���q�|���(���]W��s@��c�����&��F]�P7�)�F��n̹w7}&/$;�04a�-�q�3��>�7�����b�/�HXK	����J�OD��T�ꕲ�3ȑ*Uy�I�r�ugo�dw����A�7Q�S@�tR��[�9�H��A�}��Ȫ�˱�FS��2��������Ce�MT���AH��8�aD>�:SH$;� IL]*�>�8 t��t�	vb��[/����T/��F�t�7��u<�W2,����y��S4�*/&������-{�œe���[v>��oNr ጖+n�y�_�{�_]B*��h��P����zu��wlw�%���>$ 0^���7���,*ITqg���4���V����0 ��,��E�Ј4�A"4+�?2���@�"4X�9��\ے3Zbąa9+�'ܥeR� ��L��ϋ�l3ZB��a�p���'��aI��`�����'�ml��s��5���~L��Fu�L@t��Ss�l�ZHB��B��ER�=�:i&U|����Í+9�)0́��$ҡ�{#}�[+/V��iXjO5yrP6�.wW��-]�1p��&.`��ƫ���_齅I���@�`��@���c*׺�%���`0l_{ȿh�Jz��y���m������=�J�)3�9^�Z�U�E��I�j�Y��k�[H�GLą6ey[W'h����9	,�f]���+8��F�b�����Ȅ3f,]���ٳ���� ���EU:Ad��Y䒬������/Y�Ҿ�VW-M쇼��[DLV�i�1L+ӛ9T@�MĞo����3��c��������y�4�".
����-�7wV�$pX����S�
��ir��ۉ����2�wh���?��K�9�r��f��l��� H��6�:)}���6�e�_��B�y3 ��Q6�ɯ�U�?
�\)��k�RD��SN*��@}�0��h�`�OB
�o ���2渇y�Cg�O�p}�u�T���]�t�h�b+6��vXcD�<�/�r|���A�:wh5ܕL�l(�]�â5�q<�'zR��p��4,��;`�#h]j(�J"��k*�;�`.0��ZQHTa*�Z�|�$ZϿ������m6�Rq�lX˃�(�_�}LhA�Y����lP9 �	=nZ,�Q��֪T��P,���Db�����9�qީ��PY)Z��$3�J$0����H�%�����.^@nr`9��э�<.T�8��ď��L�G���������*�Bv-�3�R�4��|��*�o����OKI�:�����w4��|g{���j��D��>���Jc���3���>�H���E�_�Ɲ�깱�ud�0
�ۭ���O!�	HI�q�g�eJYȿ�L#ip���	��I�w���=G�3f�;�z�*@j�I�����W��0�ׅ�on��*�IzO�.��1H��"-Oq����Y�A�)-����+|u)��������� 6�Nbd�٢v:.�}��}(�{z( MAIO, �7�}�nֈ�����/�"����=ޱ���FUgW�Ȱ4���ʤ�Av��x��'��ϵ�j�3Yl��Gk������ $�d�k�@/�A6C�&���1���[�}r�'ʏ bZ~e��k9av�Jb>r��ԟAKF�[3%Ϸ��}�ܙ���Xk�?�z"�q���@�'�9R E���}i0��is�qQ�47�kыx
I���Є�5uv���.�@G2��b
�XrN��	����%��]�[ۙ���ftU�a��ΪaKpق�4�.�`�����v5�b��3�	n�6�kj��?�}l�~6W�ݜڻ@`�f#u���0���Eyq��~�nP�,���1X�#*�]7l�^$�PM��䏳������r�ȓ� l�gs�E�r�sN��(ָ���kO���sV$]Hk[��dWcaЈ/Uڭ�Ɛ>����w`H����L
*�S��<U�%��U����|�Qb'X
1T�}xHL�h�f�G%�syn��dd��C��S�����E1h��p5�_��n��x�3���ӄ��P��g.�+aПv/�%~z~�������5Zmx�v܏4�(�XP����\m���%����:,��1)���,�R���x�ĭc%�#_�`�O�7�9�G̹/�Y�kc �4�A�������vu���Cʓw�/��3Ջ�}.��@�=]F�p+�� ������V�!ʃ���/�	���zG���8#s���t����hřqLג%{�2�z�&zO�Y�F+;�(�`�ȹ�f�4�-��i{6�m��ն�m�A�[]#M�#;��=�*��.����� �g�<!��IT�] J��Vk���:?��� ��Ql�ስ�ыT@g7=n�g���"I5�\��TVp�3�k�س�����,1y�F�`��f���|B0qԴ�rU�stte�w5`ic@}�p��72�k�f,C#^���D���(Nn�EϨw�{�\���5l�e�[@����<S��/	�����_��
�U�F�p:r���Z9��_�e��4��O�
yǱ�ǲմan�1�Z���(�U�A�}4"�GMk��i!�u7�9�,��ɋsr���>�k>!$]
貄W���u=9��ߍ�=Ě3�&�b!F�L]�!v�E,Q��-l���ȧ������ã���홍�f��Ln�f�N�0����{�O�bT��_g+0��4��Qe64�?�w����5!�7W!_H�{z"��͘�X|���m��3�k+ �Z��]+̹
y��=�#���ӄ��A�I'�ڐ`:�l���M�W]��as����^�EĴ���~D����q���]���+�pt����'(�z4$Ρ����ف�'��+ъ��ƨȵ��>�HjR����M�B<~����ZވG*��u��w�G~Xۯ Le(����¯�dB�%����S+I�,Da�TM��^ۖ��S�<F3j_�"�����g\�J��\XVe/�v#uI[k������͏1_oe�K�(� ?4�G���я5~�YM�(R��98ajQ
�����G�D����ޚrel�S��@(&Ǜ_�����+g���n�lQ��۔h�Jw"S�=V�4�3=����!��o0�ȝ�E߆��X�\9�T8�ݽ?��ƈ�\�_��τ9�	��aB�����p6\u� u�Rq#�둏�K]&������Z~��l�0�#FM
�Ή)L��ؚe*GT��ߡ6�c�w�P�L�k��I�d�Sf��QA�6��`n����L=TBM�t���ާc4��}F���䊧wԷ��G�2	����Kmԏz$U���E�=#s�R�@E}VR�X~�[ȫ$�|1�Wr�1�W�(
^{�����GK�f�2�P"��3L��(Cx��8�c�Ux$�	��&�?�����q�\G��<�8{Ֆ�&\���`�E�Ӎ1�5�9J�@������\�Ǡy��z��d�s��N����{X�Q��g����n�٩p=������=t�;KStp�F8� ��Rq+��.FL�#��4��Ez�$�8u���?#<<w��~N�(]j�N"�H3���ъ\{�n�0@����4�l�s�F��E���>v)�(*W0�ga���G�ZM�)�Ps�NTԑ�V��_��*�r�0~k�2��{�ѪX�H:%#�����|�_=q���²X��
.��DY:�|@5|\���iC�C�*�MϷ���\�z�D1g��CI �L�$=�m��f��_�����,��")rU��	�q^��Z��_�-�Dܑ����L���-��ý�?L�K�a�o���d(,��-�nDg�ڦU���=&)������_����;h4ie#1|��n$l�Y*����@L��Zn}~���Ҿ2��zX��>�7S���C׬�W��>��U�D:&K�U4���^����u��K���X���IV(���]��Eaqp�^:�񛣤461蛩ʼ��t�V�/1U@ϒ��'j�M�T��;�a�P6�ˋ0�ʕH����;/�����@,��U�,����TŊ��	pH�� �����$Z��"RY��P`�jp̍&Rf@�ߧ
�%R�$-����|s�Nrs/�h��4A՞�<�7�:tEv>�`���&}�$�a+,Q�{Z�#rv��A]�y{�T��r��$��9�b��穚����,;��f���?:�,E ���'�s�'J�$����$�{�^�[cw
YM���0�۞��G���c��b�1����Є��l�oj�>u�lg�j������:H�cB섂Kytv�0�iO��e-�,\Ԩ*%�dsĖ��4J��D̔%�2'�𾳏;�ҳ�A��)ؗc�C�����\=S �K�
���r����J�4�M���3�����6i$�J���0�p9��m�Ґ��@���,d��+0�:y���Cg�:���!����`L,���\vY�L��$��F^����\�pZ�$dU $;�i-�a-����X�3��(��b=����fNH�WZ�B���F���&��է���'��I�Dg�+����<F?�m�ASd� `#��L�%0$
[G��ц���W�����6�.�m�p`ׄ��%QP�����?0s�I�D�]t���f����_��{�2�Y��V�A$/����-zQ�NH�r~O�`n4���i���l�����"�]�?lӱę4 mΘ��t,R*�S�o�}�1�������s�=�Yb;7��y����1*I�x XI��r-R�d[�w�mAd`�Z�ƣ�Rͺ�>@�1hm��D�q��qy9#�w��I�꿁�elؘKU���g9)�}}=-tB/����>U�R���P>�e}���r��N����"��0H��M���h���Za�6�A����FQ��bq��$�"�K.,�|�9(�X��yJ�U�	ɚ�o�0���%�c�
e< �ƈ͔y�����[�����#�t�e*�w��Y~�wZ�o٩g�u ��(r�Å�$f��lD�!�����Gf�(��l��P 6�X�NI�.Z��p�h%&E"�'bsS�ȵ�����=�~��$JX'�`�	�R=$�2צּ��=:g��ܫC�o�	��31I�^���6�n�Uԛ�۰��BBީ���*$A�삉7��?h�����Y.��Mt�FC��[���Nx�jn�"������n<���M*���F�I�}Sb�;�,���}z��lj�#?E�,���	�(MW:z�������eiӧ�Ū<)،�\���cw���*p(%�
��HM!��H��X����*&k؝�d�������:�	�=���9�5t��CoItGj��lW��%L�m̇���E8�>��LX��d'�>3��a�R0���3�0�;%��E������-h�F��TR,%Uy�V��;#[ �ۯ���3Ra2�;&�0bt�>���<jN��������c<0��ﷶ�^|<Ici��~д�%X�7���m�yzͨ��Q�h�<6u퐺�����Z�[7�x�N��dB" ԡl��%y46�b��#��n��o������+e�AzdǾD�+t�#�!�u}�eC���R:�p���^�p�����RH��
 ��\d�1���+���gOǱh��'j�6B�X��o���{u�^��$3�W�P�H�H;��tRii�^�'2���Z�߆i�^i2�K���)���C��h�L�蓏\*��H�Vh%�����"e
�#}f�v�PkVՊ+֚�0X<�|�iHYf-jh��ּ�9t� ͎בW[K�G�l��e/����ı�J����
�f�E���BX]�b��g�TKyl������̞>@�ja�xh�����'��g"㻞��~j��.�zO�ᝋ
���%ߕ	mWI��5ä8| ��>1�5��_���\<}헯�ۀ�}����,�*J��O�(����Ǳ���Ya�'�R�~��e�ظo���-��V���2x�J��{��މ���ß[*��m�IR����S�cd�SL�/��Q
��F� [��r\.��E�b�p�h���2a�:o�j:�-��~��Xp�/
W���,6��3��A��_l�Hn7�Uy;)�k�8��V��_�Lh��k^_�Qm�����z�1��>�@C���d2�ܯ����x�uDEJ�dO����:]��<�����_�2���c��#��q�0_���
�Fq!�]��B�l�l�#2m�+��c(`�;X��B�i�X�"8`�"�?Fr���f��ަ7��6�����<��+�U��`�V=�?bA I3�M���*X��a*)]���-�l���?N��K�VI������ط���h&��d3̂�InHZ"������(�O�&�����������vIC/8`����}��G���&v既be�ZE���9T��ӡ���1]	���l""yq��u��+��-�c	�0G#��| ��Y7k��oSý��7 �~���о�����&�W�����x��ȟ)@[~�'}cǫ�8����,r�^�z�h7
�*�.sTOl1"H�R�s�W��ŲT��,k̹�Q�/�zz>'!���vj�˹����:���	���7X�P�[3̰_�]ե�E�]���ӐwD��Q�n��,*a�I?�0��h��@$�	I���z.}�mF@�3֑:1�=�����<�c�����؇�����l�u��|	��U�5����Y?G���F(�0�y@�J�s4	3�M�zE��[K��x5W��ZlU�$L��*G�R3C]H��Gd�C#����4)t�/�&���b�"���n��XC�|:�U\"�>s�����Ϋ�~'l���g$�'��ݾ�̿�DD��V�3i��Y:a��L(O[�]�u��	S�E�2"Id?����X��vU�����L��1�cI��XT��#c�G�����7v4��۔� �*�vp/@�z��D����h:��=0�N��P�t�(-�E��P��V���m��<';�=�R?��i|���gb��g�� �C��\�cA�"1�����Rœ�D-G���#Y�bz�`8����o�%��4ٰѰ0_Iބ6̏S�?o�=��Xwe]f���;{��������8��̥�9vI߿6�Q�����ۤ�3��"���g$�vZF�@�GA/8��i
����0,���A��ɲ������n[��o�r؉��Ll3^��U9%X���K���pOaPf77N��_���ȿqV)�xm���y�~�L絔����u�G��>N�� ���&�ؤ�)Ҡ����d��`&\�.�xL��wՈ�v��À��;QN+���ߟ���";0Lo�HCs�F�����xZ�cY���:[��.��K�j�#I��,��d�k�����6��ф�.l�B�������D����x��i�Uq�����\�o"9�h�~��]qW�6�!�ԭ)��<���oÕg�;P{	�Tԫ�y�>��TO��캔�h����:�$�W�W��˅�p��9i��H�F��O�G�����s��?�Ǻ�ш��'+�CT�O��λa�z����>�3��E�2.�94@�5�g��Yh-���ܳ0/��x���<���;���W�vP�؟e�И�3f�S��Q�`NR~y�Od��i_=�𦐹���{����	���>y��s'�;�3�I�2����y���Ia�<��L\��T�;E��L�����nu6�y�@A��L��2{᦮T�����4�$�bY���x�W>�&���sJ��[�ט��_�Y�Jc[� `�f�_�9w�P�s.�Ouq�yhx���)�i�����TB	��&��y\K���� �3�ҳ����5~z�N��G���K������Z5��|G�ԝ��T�'~�l�m�ze�1F0�CH�z��p�� z�X�yϴ~@v��:VVV�p�[ ��B7h�n_-�;���x�v��/��*~��Z�G���0��x����!��!�J��<U���L׽�ts�2�<@�F�]�3����QN�C
8m���N�[>�f�0�v�(�O��T4� |�`҅��`/�nJ������["��j�����Y�����'�m��:8,�Y(��+�u	��[sޡ@�3�9.d������Z���C~��R-a3�FT�)�\fO�urIt����?�*ꐲ=����n5���9U`��%pp1��3<�\����h��{ӔRGdTI���1u�{�n�1q���� 3MV<E������_�X9�&Ŷ��e�=�&�� �@����?�Z���tt���:׸)�"�Fb�b���srvG��G����h�YaZ��Vˀa�U%���*ʄz�1��W����e�>��"��$j�m9(�7�G(�]Ĵ�pF�ʳt�>�@{�ν@A�7z%�'�D'�b�G�����4�\�pΡm��C���P�&�J��2����=.��#�?��F`��D��G�R�%Qxvp��dz����]�k��>��o�o��Z��YPd��������&6�P�c�)�$�贐'ªa^���9<\���q�&8�83��'7���]�$�@=�Xg�4��Ou����KѲ����/�~��L��Dʽ<-{n��j~GS�<��9��8�Mq}����-��	�ڬ��!����*w�7��:@�Hsy^i�Y���>)?u�=zxf�O�`B���g��.0�&a���׊42*�/o��(T�4��Y�����e�'Ix�h{�1����3����X�V�-�h��~���x����P������zl��Fv���R��8�|5ܬ�e�~<FCg��|�$m�OzQD��)��X.��g���{��<2�D�S��/F7$K]��t�HadSB}���ڋ�&Is��O �c�l�X�,����
oL:�p��1	xiD<�<u����J:}H�e�\U����gn�}���R�.A��nF�^0�Ky87����,[U=*�R�Y��W��l?80D%5j�/� k��t�>;��3��<"�[�˭L����^�q�	e�?|�TE
{�b�e�PN�����Jg�c �D��m�piI;��+$�7���u|�U�fd��n�Q�fm�9�7W����\�?����9���8r�	�Ceۢ����6�X]�Y���u������?=(Ev�Z-�\�p�rpH)	�c~9D��Q��In^[VQ�,��/"�;0�s��'�.����%��p��@g>�M�zo��'��W�8vJ6�:b�l��1	���Θ]a�}�kĝ{g�\0�����h%|Ŵ?�Y> #���e�`���d���J��.5�p/�P(�h�w�CQa"ۓO����v_�:�7j,���dM���X���,�a�J��ӓ�<��nj��-P|��ٱ���5]�W��d�U+-�0B���_ɲC�"�)a��f9f�'~Qk�>���3V?
����許y'x4>!\�Jp_�g;}��N'/��D��U���d�]h �_3j�6`������36HŲyL�q_�6��\3��ݙ�pG��mm����<�����guȜbH�>�$�p�U4�j���H�f�V�!"\��n�a_�8��髸$��+�v�I6������OU��GHj��@J��\:l���?��E2�n�9�қ�d��Vw?�jD�,'j�Yp���"R��H���f�4�w1�����gw@�Y�cvX�1��C���C�i��eѽSM}_��^;s(o8F���#����RU��3�ۦTdvaF��}�Q-��1re�*�'���^�^�N7�ă��
;Σ�=O�+O6m|j�����Wt�~��_���Gj�u�U^�JJ�]H.V;��O�k�d���}�K*3H��{i�]u�VO5�*��1�EO|&�ԮfMg����<�r��^�m����k\�25ˈ�&_�T���o���t;��~2����Y�)/�	����^������̔�K���X��G�z/���|x�-Sx5f����+�_\���ڌO��a2SeCN\G>�5\h���Y�C.E��v��nY�mG:q�u��N��|�tZ�v�ʫ'�w��\�Rl8j��wVA�{�}�S;����_�趶�={h���/�lH�5u�7yaͭ��0���0�>�W�V �Oי{5Ǫ�.E�0a�"� �п߰�5T��Fd�ު����k�sݷ�.L&UԞ�[_��}h�LU/h_,�.o���z_(���P.P�؇ _���UzA���9��"4���JG
O���9��i�K�_� ���d��{*�WѰ�a����F�'$��J#��5��~X���r&Z�iנ��u�L�<�M��@���}6�� �w���O���sb���Y,<�ĴIv��(�R�E�W�Ԋ���9ZDw�RЮIL����q���Ķ�a�̠�7�YMS��S/�����.��!�҆)�d��6�+��?���9L1��q�ܗ�&�%d:.PG��7g[2�zP�:���u�8�U �m'���L���gЫ��I�M�U|"8����)�����c�����E���
��ZE��T��\s�R1!�anY`�3t��R��X��x����n­$����z���!)8�����Nz�O�'i�e}�k�Ab9!/ ߣٛq6��oB�Cc�n�p��I#I\�4���C���ǜn)�un'e�bM��W�*!ｧvo
�$ڭ���Vg����^ \�WmpO�6S�D"(��}׮�+㽣V����� ����τb�J�=_����M���Q�"����[�LK3�Ï˂��Ku	�	[<�8��-2��5e�GvAU͚�>���C���$�E��LF��a�)YU��R��
�yM�~�l�G�����y](��⬄��]s=m������'�UOͳS��tϢB�t}��,7.���U�����*r��*��Em�Z��K����w@��e�}}��eۻನ�, ����H���]ܸlVG!]�j�J�h�/�ε��, �H`�ǣ:e�z�ƃ߯4.%�!]{_�\�k
��T�NI��1�e�t���f� ے�`*+��Q ����}��0)���Ee�ӌ�����*r�V�ME֔|��aSU�%�:T=<VvI���X �7�؊2�Gm�R
�D�MR�D =������a�� VO�?��)�O�G�G�s����r1z1-s�e��ݫ�f����Q�{v2R��ܻ��mK��ĩ�p�u2"g���I��v`��� G���̾RVa��q�;e}ǆ���� YZ�^ԣ)����F��[�{Q�d��f~���<M��r*�ƕ�x3R���ܽ0�����wѼ-��\�g�4)n���
�^;�D9��lA�Ǩ�CБ(�����PA%M��L�G��C�/��9�[�g����~oJs�+K�Lt�G*&��!��{2`�53�0d���vR]��e��,�%���G+��;�O'�;PU��x���o����z?ex�d^����V�3].�?��J�����&ъ��A�1�M:?���>������}Ǣ���u0�6G������nMֽ������U��t��a=ʳ�i����ʴa֝/I����e��s�Y�7wy�*c?=�/��:��<�4F���FPߩd����H�*��S�E�
W�BԳ��$w�B�>�&�<�0�'�!���z�#�������"v�;^+����̨]�o.al[X�8Z�giKy>��	J[�g��f�h����1^�y_��Oث��j��!�&�Z�h�{��erq��a�ZA*�+�%V��-�|#$�������`e�Em�S=7���� �J�<6�
	���gFM� />K ,�-O��OJK�9E��T |�^��GB��U	}×�v���̊��9�B�N)%��~��=���y�kbsC�҅�_��M� �|������0fS�CO�Q8>j��c�3ݮ��΃�;Q�� 䠻�{�e�3 ?�b^��m�?@&��V2�f�T�*H���� {=���%��O�t�wE���56Y�7 �A�sӪ_�@��f���4�<^�ױ��-��Z��k�×�L��laG0�ŵ�
y��q�a�R���G��I�d��q�iwE�h �(���9�K��s����Y[8)��Ag�n�w���d�^�#� ��u�����Y2z
�_�W^�����%�#xȄ���`��>^�dŰ�����D�vv����l~�G�+���cԪ\�� و��b��@�ZR
��G/܇�Nž�I��2�n�u�$�q������X� Y�:�w�W&o�:�uѰGU8���@�?�<1OgUX)?%�K��>�AӘ"9�,�)L�O|��$��J�d�C����p7��(a�)~^'fC�o9V��d�J�-��.�t={��d���ISZ��v���Z�����wF��ʒ�T��r��jl�?P�:�b%�z-�����y�~ѷF�m��}�-5%$�@��o]�Cn����A�9u4wZ5���� ]	�>�� (�m+E�.IS@Vf��ew��$#t��o^<���CC��f�� �o��o��u������]���:���	��.��	˘Ocs���C��H�]��%X���p|u*R
�K9��)�;S�\�6�!���Ն��qnQ������a&Z��5���T��b{,�]pq��6��ڗ]t������ƣ۰{��q%����|�og�I@AMn���*:/Ja����lP|�Z�s���!5��kɒ��)꼭)��{��Z���]�����nmI�t�Y��w����ΨaX���6 ��H���U�����E����^CP�s�"-]T�#/9���U07^�{��-�i���(���P�Di��Ytx<���C�{��MDs��1aǌ�!�{DF��Ҡ�DHbT��vw+�[�r�!�t��ٌ�,��U�8�0eѽ����'m�Xt���2��r��/�Q��]�١T���x����bx�l߭���f�J�q��G/��.Y��H�>KA�S۝'��+0�i�HJQD��#>�=n�z
�됆�!L4�-ܴI�Zc���Ռ#�\��׆��F��u>��2l��A*3�n��?>�� (��^��8�r����Qks�t�"�2�a]�Z�d���W�>��3�;f��O�Lp͂�o6PO����0�hW�.����b�v\G$�KEbWQ}\�9/�`�7e���߃�=sätV�/&��1+$�pRm���3 �����!��TT���hi���8�6���$��Ir'�Oy{�^��;�snC�����C��b�	�R�գ�u�?�63�!T�ѡ��~�Ğx4p0!��`�ϲ]�UŉG�՝��g��Qu����q1�ez�� ���lH S����Z��W�PJ_��
'S��3*)=)�!�d���m����M�S�s����Ui���s1�=�~#���h�m��K5#�N��M~�;^�B�@�خ��K���Sm����j3��hp��Rkg��֟B��~�*�����D����y�P8#���$�A�Hb��WN�|X֢v[��j�Q*9z]Zq�XvI����`@��'t�����vGCh�(�[�Z�x;h��6dwO>�Kn��`Kd'q�go�H{�ئf�hA�kH󎺨P�}HR�� �U��}������KyT�EsB#s�Dޞu3r2� ���b�'x#{�N��*C��~�jjCUzP�#�f2���a<����
L$��W+�Ȓ�xi�0�ֹ���7%�𯕒�����1�5��k2��#��s��:ߤ�.�C=�	 P?5FbM���xV�%�DER'XN�#N�w���g�(N���@E�`G>�C�j"U>�����N���R�y-K�bx��0�O�sS|�Fl��sWe�[��?r�?�^́�B��������[X���4�ESc���6,~.��r�l�"!��J�]`����&;����Wj��XQ���T���y2z�p�'w�d���҄�&�/��@wx���-Ϋ�ok����د�~���ރ	�4mo�Z�#�z�0j���Q1�XE G���: �y����3�7|Cq��(��ҩ<+��r��̱IJ�g����k5��U̅�0t���j���H���D�D�E_�W0�yU�AG�{,����7F���C�N�����h���C5�6(��x�>i�6�Oز�J��?�,���<cL�bu��Qg�ߕ�V�C�;�R{�[���(�igY��b6Q�#(�0�"x�`�l���P����[�����	��wmV�A�{GN��i���I����1���mu$cXSL4;�S~:RG2�*V�o�@�(2�t��e	Ց���B� ۶�`>^4M�W5^��]-J�D`�ƌf��$8����uY� ��j{q�Go�ǲ�96��_�J�<x���%XV��f�%~�T��1S�J՛/�gN�d���c����PMH�4S(�^����)_���2��D��r=�DZ������e�A<���_)�wr;#Q�n��w����q�X(��4��ࡠKx�]&M`t��U~P/�v���v
�
�:}��uAW�$T�,3�~7�w(S������~f ]�]{�&; �R��a��sV�+���T�-ė*����$ '���8x�����g2|�|��+�:_ݞ�Q[U�+�bch{6�\��c����N���6�l�Aii�4� K�2J��0_�#���8�c6֕)����a�<8 *�Wj_F��Xn謩�con�Q�R��\��u��rӁb� ����ʟĻ�� �R�'�T�>7���-�����H��|)����\��[%�6(�".�����>�\}߇?I�H�Ћ��%�N&� ���y�/ДN��t�T`�ǽR}v�SU���\%y2�0��L�
�z����*ho�e�߱Z��O�t�{�J`��qHr�	|��QJ���_uHs0}��25���p���v�'3Q�,w��;��3 LS����^rU��v@�2��ȫ�nfH_�N���2��u�<rv�%-]O����"�Q�_�;�E��\���#�n ���)I����OLd	�S<tt���u��3��-2��vL1� ����
Z�8<�a����{D��
�T`tD3>amqJ�_�x�|'�E�)/����y�(���
i)ˉU�j��s���>
�4��	� {ћ��o�kx�~��>��(����@US!34�V��DL����U�\n.j7�1fݝ���I7 � �ɾ׊͟ù���Td ڳ������)��M�f��3��^2,�H��D=�gp��H	H"7m���v�k�f�X��%��wO��������8l��ZKM�ڕ��[�Ph_M�o�:�%]<:᫉2߀v��(�9��c��u*C��?@�,�����O%F��J�/��C��̫ן�ͳ8�s��6�L�鑻6e�t��݀q�Ux_dm������)���]���²ɨ�8�M_�Х�#����^yA~�R��>�n�����=��] pD��ߤ��1�yI������~=F4@��d��4�6(һ��=&(1	N�nȫ�H���Z�Ы����+O�Z�E��71������(����]��H�a�U�&��2�u��$Ѷ|A��:�,FQ$F$YU�b�~�X�jn*U��Ojs���_C�Ys�3^ΤmfbJM�������t�JNw�����{�`d�":��¨��z�(V�;8M"�������L�B���a�|d�4���J���tC�*ք1����w�\91-Q���@������˷#RB��ɏ�㲀�} ��ݓfǀn��P��\�Crv�$���lW��E�]�
G:��&o�.�D�wL�z@~�Q�䝓\���\���֔�N�[��ߕxw�;J4�H�4!�R����XP(��C[��&`�X�"�@+>u��qmՠ �8�Ҵ �IG��;��ɕ�Vu�vdW��!SR�dsŰ��c�x"C{Q��e��e4|s���܅�����1��$��/�[�$(@�{�t�O�eō�p~��������K�?v#����X;����Ōk�yy"�u����9�+���K!���oP�2��V�P�J��k���|P8�Pp�G	t=�KVߗ���&����av~kd�����E�\��������[��!���	�-��I͸�M�|��U��n5���
 �6ail:�pWF�&I�]ǭc�U5��Ҷ��2ܢV�ݢ��`;��Ku�ܮ��w������'DQK�g��+�,�I- �Fd ر�:�i���I]�}(3%���]��n�DX����Hԛ@�u����@fnA�\P0�b7)&�
�`y�Rk��fos[����J���������F��0�����v�e�bv3���E7;�b������|��a�7?��~����ߑ�+���VG��~���2sXn)v{���/��(mT�A uO���]���3�F= G�N��+�dn����",�r��~��D:�h�l�@�a�{-6L�q�Eu�Fk�,��7�Pռ���:���4������ʂ@�!v@�c���~C;P�������,���ۨ=���,�5*��od��x�X���j��`��j�~Ó�HN�}�Z����6a�-EY&X�r�4��lk/�[-I���A6.Vp���K��U��пj�)j#�?����#F�zx�-]�(o��^���!�m�8;p�[b���6����ش�
t ����We�A$�2�+"���1ot��Q����|_,�K�T\���x�A�(T��[����5��v�2&p�=�N�
M��bԪ��$��к!�Rk�SH���=���GS�/��\�d�'�}ǣ&Jd~s� �m��*XWI�v����������lR��K�V�$l�m�︙��(������3��.E�e�:�̦�]�N�Y�a@�q)����Ј�Wf`��]���4��(�$7U��	 \�)������KG֮� �{%{.e�"me�u�U�正.�̆	�"ٟ�6#7��N�� �x+ݥj
[�nK���;���\����́i����D���z�V%%X�;
YD�vd��?�*O��g ��gp�1�P��Ix��pfm�fQ*-�'���ȥ���Sd/I�9���Co��mNVr��_hHR6*�Z�b�UT%�Q*�Ͷu�>jr�~gL6nKg0u���{p� ��B�]��+�pCw�0������Ύ5K���r24� zxy�>�~9�ߣ�i��-�����o�D'���M\��}�%
`B?+���b��/c~���Ah��V��Px�@��H�s��N��YZ�+�/�4e�~O�I�v�� �]���t�
�&������:��t:	jZ���z�P1h2��-�X=�	X�H�HX;�k
��u�ѝ���*����I�IP�R�������ms��zp�S5��H=oK�]6��Z@үc�����~lXel��r�ـ���2�&AODAPSFq2j�������5ƽƟ�- �Z`"�/��1XJD� ё��Hؓ$Je��$^ ����^^��岒k�c��<b���t �?LP��Rȹ	�N�p����l]�F�Fs�L���xA� �h6��-�6���[Xͩjt���G������j�}p�>��~�Ca�tg(�U �̵E���zl
�R���&0Y���O3Ub��#E<7�X� �З
2�h���� 2�C��\I�vO+�� hl�h��! ���� N���O��V2���X�č5$ߋ��{�n��.�Mt�/��Z`��I}�h�S���i�ۙ/aR�~�p�׍�^O�'$�D�l��w- �ڮƯ���dq��Zd�\�~Ӵθ�I�1z���M�Y��:q������':�;z��E
��{K��-��!�p`�7y�N�Q�'�E���%g��֘���Q�5z0�-�m�Pg/J�aS�\�����XL�z*�D�	8��k�gCy�x�%lcn��n���#�����ܨA��Q�/r�`���J}n�����q�)hy�_Hf���:o0_�č���=c��4����SXx PJ	��.��"�����8��2h�ΐ��7V�oGP�Í�N"@��^瞶y��r�=�ٲ�=a_�6�U����kE���
�kۉ�N���ڟugs��X��g\�9�Uj������.$Ƚ}n찼NOG��1&"<�}�`�lFQ򼊰h/�z�"���n�|ͼ��;���g�˺�|o�Z�BX^5R�_V8�֞y��5J��8- I�OR^ܢ|0T�'I�s�t#Z=lwd}����>�R8ZȒh��t���c\�_�G�U!�Frכ��(�dh��Hg!m�
!�"����t;��d�2|0�y \�;�{�B����/��U����GZun����A��Ӎuˊzg{A@ҬBm
(���k� ����r/.��\1�F�ev)I�^4���M�@�-�V�r��^�kZ��R�p����2`��eyf ���v]ǐ��k6�ﶓ���@!�ԩc�UAa���A'�w-��Ci�c��{g���^&���g���Ҍ�yym�(���{l����U V���X��!�eQ�0d/��#�3t���eRk!��f6Bl f�>h"Y����Fh��ՔǤ�S��~�e-j��H��!6��+��\�t���~��q�rS_�� ��=KN��?pI��*^vȱ6?H��=1]�2�x��Al����va��Ccძ��d��k\^�ܣ|sg�``�BྣΡ�!�,D��4�]R���gv6�jJ¾��?͑O�ʑh�H�еuB4��k�����(��-�B �'�\އ��4Fo�/{*�T4ׇx�_�_��(e��T�*��jy�|h(��������3I	�xq�{��0�W�H~Op��H�r\���<�k澞�����Wۮ�J�"�-]o�5���'���݃�XE侻R��T@l2��޻���vr����9�C/��]�)/b03	l1��oEζ@[���5�3�(c.N���ɒC~�"���E��wьys���s3Y_-}�e�I0~V|�O+g�;�y�[v�K���p]�u��'�u��|�N7��Ů�/Jg�-��'�	՛Cg���My�_a����iI����o���&����I����d��
o��y���4��sC���brؕ���|mF����R���$#v���W������8A�vw6D_�j�B�6��{^!�O�N2���%��@��T�{�p�y(.�q�ej��/�o�h�O<�K�� 
�~	�t��}��/�XxY�N��^lg�3�m\8�p��ҽ��Z�DZ���q!}9��3��@yB暨�sS/kiT��m�R��_�����(��5j�����!����e]��q��'�	f�+ކx�:�4�&�i����x�.d��d%lY�A��/��h>eQ+"4�ҐxB�jp��S�67�����
H�:�\�F��N0�I>���Pݘ?������m�O5ӡƩu�r͗ø��@�&����&f���&ٙ�;jU'�J�����ߢg����/�'��㌈3�U�N"��y
G0�� �'>=9jo�NC�xa-����>�MCJ�c�2�|�a��<��f��٠�_��8�4�k7������i�$����Dw�b 2}A��!�3$&��uA_By�}꽙}�KW_^T��vy4K��%0^|���Sc�2�X����KR��c~�
By�oX{!�Z@���Gsnn_��.�z�C��2����t��ϴ��؏�\�4�(��>&8�\��&�+=6��]o,Ћk��x�I���d��q���5�� #�t�G��yY�c��R����ݞ��!�S�����(f�K��m�ơK���E&032<�]��XʴuN��f�ؙ;|+z�S9^ZѶ�nI�湻�/���7� �����F��E--�X2�&�*�]v!|e�ŒP(׼����L�c�Iٜ�g�?�`A�U��꥞.��c��@kbQ_�@ZkRc����e� y�V�CO��"[��PrA~�����p��S��I|�%,D��Tٸ5�-�9�e}vI��](�o�W����<�O�u�ӣ��%����۾{{�b�N�7%�Q`*Zd�u͘�smP�U ���Ʉ��}r�b�q-?0�dq��!�_wN�N��2��Hצ�n��[��!$��m�O����[�+��v.�E� �G޺�������$�:o���[����V=��X����W�!�̑`Ds��1���h۪��?4��:ևU(;��T_�U�xy��<����AF��׉��Z�NK�gSsխ��o�
��m�J4�4SF�@V���H�����e����TU~k�W����:ՄO*����;{���=�HD�x�o hxݕt���`eLtu8W����J@�LBM�?�8岊3�4-!P�D��=cӏ}�ؒ�4�t�ZO#؇B�a2J^*�nQQ��vG{"E"�<���"X���Aa��)%�t�`���d��iw�����A��p�~�#?�c�t*���񙢞Q%�5Ǹ��c�Wd�7�K�;/��磿�ÅMO{[���t��-������|K�c2��:�lT���<=����[N�{F�ԗ~~���T�J�'Vp#�����^����-3�א��@�,���$Cc�Gt\�VTO2�8��Ģ��Eڤ7}�o�P�q�k�b���}����D��"|�Ֆ��[Zc���V�@��]���d2�N���D���
�����L��4'�a^� +���os��jV>���}uޕ���Y1����Q���8�V9��K��	Zq�?��J�u�?n[������fw)f��l�������$����D�X��C\�1WEЪ���X�%��pUC�{��(��31�"��G�~a*�pF�Ӕt�K�1%�
�D�n����Jx��f�w��ce�])�d!ȧ,�<��o�58&x"�Zp�g�T���1���F���o\�7���X�Øe�ε��=��[6E�O��د�[-v���wmFK��_�4މ΅7����T>���ŰQfb����{�+�Op�kg��"~��yf�=�tU��ϙ����	-)_:G?��}~�)����ē����_��F�VA��J�Ӗi�  � &q'�zt��ӱ�v��ݙ�0�#��{�fP�bg����'O�L
W�f����GA���r6a�t���2�,�y~����ܚs�AB��8-���aW�-y�z���Y8��4�������o*�� �KgiG�W���������_�aC��	�������moN_Wd�{;d���y8>�',k0��p��6��U!�qb�V,�##����{[���x�PF�]�՜�Q�}�~�7����T��yz��.n
b����� ���~�w�_�ZX�凮�qx�Ɓ-���$�Pj*�HkȎ��	�
^���\2}ۑ �K��2��a�Y�����s����O�}�N���I{��}�Q��3;��z�H�.I��P^��a����^ҿ���\�-!{C��|f�[tYuX�ɑv�iQ�'�Һ/�R%V^�<��m���NmY�u�gܒ�/U����),ɚ�ig�;�PA͙d�9���p	9������㯢��,W���_�����:�I�剓��1y���z4A+y�]˟�h�$�|F�/�?�z��k-&�[��6[,���V�H<x�X��y6'�e�i�{�4���!h��Ѳ��(z��p��G2��?��t;�\^�������O͟�є�Q3	�2n�\��X/Sg�J<!y8q��_�^i6�Z�6	�;�����|�t��"y*�jSy~(��yx���wP,׺X��C��7?ƜeS� �T����#m���P3���±�� 8�l�IdAݸ��i�W�ї �p�pQ�֯R����|�c\�K�Hˉ]!#~1��8uUT�Ҁ�[~6V=�pԅ��Գ��KW��ָYZ�f��K���vz�1Ϳ�a<��YWZ���,���z��H(D_~Ym�g��T�)���`*��E%��3��te��o�g?�C4>���eǸ�3�E���2&��@Z5wC�wy��]V�0:�}f)�4�q�T=0�F�'"���
���<�~F��~��h�ꮛ�]V�j?%2�qaj�Ug5vŶ����ﴏ+����@��lWT�u
�����3���	��Q�������þ��t��)p�<C�v$��
+�竹MWa)�.��>8�n�6�Eg���� [4?�r�efq��W�p�D/�%�ʃ鸟��߅��;�a�9�O���P��S����A��%�/(>BXD�XGm�7�*�C�����5�>�iPPy�Ŀ��b�%��Ü���pgI��CY;!.|��JE�����+���|Z���.6`w�߳Z*z-�pZ/�-���(�v�����{{V�$�	1�6X�WM7���%����~+�9��e�ѩ*�2��@e��IW�<b^6���e+��d��4w��>� E�6o+U��8�QiR禵���m T���+��i��q��-�̗�����Im\z%4�7��^c4y��a�}��ur�zvz���_�e���"[�d��c�4��h��ҳy�`�%�I�6 .�a��p��f iw@`/vA<ڸQu�jj�w���|�g`��x�%0�����BW ��e�PP�s���%H� ���t���+�<<`6�珌]qz n�9��w�'����mA��7w�_�n��y+;,ğ�0R�Q���G9�BE����~xK��ˉ�֫3	�.a��ɗ�~(�)D�µ�i��Q_���hK��|}�:�eZ�2��bŧ5-7������v�Q �
�蠇�������O;�K4".�^��4��M ��tuA�C+�zw�C�?sC�b�9�*�.+��D̂~ ��C���+�vY�X�@X�g�����N*�S)�$�A0E�g3�ëm"7߱�UR�ń
�V&?����j��SDXM>fw�ɵN�ó�A?O]'�2��Cd�*/OVRm7^�&MX@�UȬ��uطR.�}�uJ}4���s�D�_��챚�j�c=dz�A�+줙%�K!���m	��x14�ܴ�-�t�72�=�P��o\��� �Pm6�vRW�+�@t�vpT��wkՇ2u�ހ��h)��)�PD��9���,���,0���2�3��i�vDP��Fe*6�TO9�~:tof���-�͉�����WV��[�8JH�+ƚ ��Xe��q�#���s�s
�H�i3׀���ޑY���@ �e���e0�7dh���{�(�_D-4h̨�t�֓ P��0�2.�k�;�K�?Z_g�-<��m��*��h^!��ڳI�(��Z&*���\Րԛ#��=;ۮA���{�LA9��8瑗��/7ld���_M"1�C[�2+����M���4�iI<�i�޸��:��(��Ż�I�6��;=k%�x��5��#o�j6=��`�Yw$b)u���[�)�~WcZF4�)s��`SH�?�����a��X]-0F�f!B+,5��$�"u�H�AT��opE�Fr�-hб4Ō�7���J��+�d6�1se�i��}��o�!�����{��K7��U(��'��b3I�('ق�DR�*��o#*t�!zNpAՎ� d �أnJ0�ʢKk�f��i=���(;��� �LX��@��W��!e�|W�gگ�<������Ƞ5;Z�Vp�Oq��ڧ˒KQ�"��ÙM���S��|Ru	�1�u	�s�5a۩��׋0?�����s��m��q������5��$ҡ�{��p�M�QgE�@�a�(�6'�V�!��M�sx��.s׭�q�9і���,!%��٨��,�\@��Y�|;3,t�E����z��Ÿ�/A������a1���s'a��*y@�He(1��C[	.�qĻʯ�uR �
�SL+�$�l�,�Zb� ~LR���nօ��@v�x��]����#Ubk��#p�[lsA9��]�����Ѭ����ɣH�#���8j��V����L��M��z�-$(�ܼ�n�����4����8����َ�{���6[M4.b|�=���������i�p:���O�0��� %,2�Wu�̀Ԉ\��)l�ȏ�2���4���#8m���s�,&��d�s�/7�w�PӉ��V��a�+�$�ܜ�P囡z �x�S�O����^�a4�1���0+-�	�F�)�2�(��p���e�Vl�^k':��� EWx�q�Iv�=���ۅ)���P��2V�#�zSԥ��zX��~�Ň�����+��k8�Eu�cXʄtP����1������D-|�o�b;m�4����7�� h=i�U˪_zb6����3�� }wc�hT��#�p!��x�/�cPcW�-���%A!8*������~'I�� ��t�j�ί�P򮴤�N��*#Wo�#$kB�E�n��E˙D0���'�ղq��\�р�WY�[
_{����EQ��M�",�JGv�(�H�IW�	��E^�@חW���d`���*�fW������6���:��Ue�>:�b��:c�lo(^�����\��������8�r�^�� l��Ќ��.�;���t7iV:$����E�$$t?�3��NV��gY"u�Pʚ���n�*�]�Få���p����i' 1���;iY1�DU�i~.��{0\9�>�]�Rb��M./O>�(��Ix넋j��a�u$��;�>�Luػ�ts��xaB7{�rp����'C܈�m��0�s��W�N[r�+��R3�X1��,`#��x��"��]dz�v�j��pT�#��8���i��'l�hn���-��]�΄�T��c�ǴB	A�m=��ۨ0x�, �_=�Mx��dkP�r,��ѳ�B5��[��(�� �����f��jф�`��N��0�7��D��yF� ԅ���$���^�0Ӑ�p������}�Ot���O����{�9�����1�f�Wi�ȅ7g��M���Q�_{.�
��e���~�(ә�T����u�♢`J�a���W�hꚂ?��b��@�$�Đ�������d������?�J�b:����F�/T
\F<��Ư٫�_�J�=��� M;{�ԗ������P�BP�&"p|�	��Oޞ��z�9Q��QD�&���^�Ws���=��`�������B<�� gN�ex9������L��Yٺi�G�%^TA�)��R�9.�V�,��SW���:͟p&���K�4���:��d�B�Ԟ�@��9][DX���q�����.u浯\J�cW*KF��n�1i,�Od���Y]B;�E�@�����D܎��h��
|m���1;�&���kW+�.+a��o�%7f�	�ß՞�Z"����g�~�� }ӝ?����]U�%o�E�As��~)�8�fh ���I���F���|ٱ������������1���ȿFo��r�A�T~B����`�)��VA*ـ;��nɒ�)kSI��Ԕ�Ʀ�He��IR�*�iq�{��4�w�
o8$�� �3a����`�,�.V���A��.#���cdJzLl{F��&���Jr�+	�<�.a
W/J\T�pӈ�=�l������f��u!2���'���ۼ�`U�컖֝���o�@:^��r��*��W�9��b紮���J�ޔ��^�j1I�sV>ŏ������V �8�W�$�����d�����_bŔ�z0���f��Z���o2 ��O�����铀��|�u��"��2�QI�ݴqNF�j�P���˯�ǹ_,�A��F:����	���?��U�/�K��H	�&�<�u�7�TY���y������O,���� \vs����Iˮw��5)C2���f�;)����!�^�����Ls�?�����s��O�;���[��Ԛ�w
1oA��[Uƃ�?���"�Pk�Ɍ9[[#3v�z��9���U��y�=������
�V糸�� ɋ�A�����;��|����7��kwi�觥ֲ\��5���\�PR��3��Fp�v��]c.^?i�PL�H�E��b���8��}�c�l-*}�vW�N��Q��Oxւ}�oT0z���������N�W��T��pD`���:�>��+�t�n]f�+�)���U+��D4"���ɴ1@�r��n"J�MnV������	�	��������h�Lb��k�E͞y�B"3y+R�RPM�5/�����g�����b�W,�G��0ʐ�)�٢�4n�a�*\���S��UZ�c�>ulr֐&#��.+�N�pu&8X�8��M�[�W�T�ϸ
�#�
�1{�<S��*���wXu2
@��ot�pd��zp_\���9
ܤ�j�1�t�̟N��.���G�@���5"���b	��o
q��\_	�/� �M!�0�C�4�s-J�8Rws3��	4�0^�3�,��fF��9E�8 q�������hU���/3p�.6^-��]��t�T�E�2��, 8�k���\�l1�D��:���+s���p)�t��\���q�e��PC�6�L��]BZ�g���������>.��0x��x�rxʟD����z���_d:������!?��j����0�شI�5k<@�qK��^��:X���W��rB��z~"�ބ_F��Nv�=�M!�4u�h�I3@s/r&Yy5����$�r�tx�pFG�N��}q��-��\<��
"٢�8���E6�u¯_�J�����Wdm:������y`�/��_� �`� ̵R������`o�?@|�X�G%�%Y�c�E,�v_���hf�?NC�sF��ɻrfI���OEd>��G��QM�����a�G�5�a�<���?��-�J]`[����(x�������'h2���gu(!e��U����K��\�� �j��_ǦIRs
��}���{��B��AڰѺh8��혒�@}Z���hp��藲_ N## ����B���p�-���%i����X�h5��0
���	`��-�ld;�	1����V�p��ӊ�>abB�x|	^���Ht��Q�:Q�CtN����D��'�c��چ����o�ĥN�BFG��f�l��/�?�u<���L�����lئr���BվA��e!��G��2(�Qh!*"/�γh�𿌋�?l���_ę�o���pm�ۮ���i`�с���,
�$:0���	�bu�G\����U(Ș�,�ˢ#A�={�tp�$>��m6�Y/."���vA����~�$��+f���+��T�ᕙ��)��T!���-�*���L��h{�1�2���4�G(MCU.�x2��S<Ɍ1%���y��7N)�ME�����I%�Up��!����k����-�c[����*��UK�؟���/�B�߷�rt]�ɟ�~$6*��W`�.�_1k��h�־:�u��dȻ��K��y�p�@^X;��dL�W�Fϧ1A*F&�rY�b.Ok�Q���!�*�AUJ�L�l�`2��{q�?h�M�ѥ��M@6���p�v#�t��_�hq�`|�ߜ�ْ8����[]촹�p���w�:�����0��Y�Ty�we!&�����d�ӻO��C�jP����m\��$� *�L ��h]$i�2'�9�rצ� )*�>ef#�2�C9zĠ ���N�fxј4*��|K0~@�����Ѫ�b�JD��S�@λ-9�2z5t���\��+�P�Ԗ�U��M���@ �_�KB�]\�P�=蘴@eЙ����d��lfk��^�1uwO�7ǣ*�}�Ar�����3mlzڜ#q�����A,[/(u:�?�l�P8��k*��'��+T喊�W����0k*���t:I,�1�]��r��4
^S��W!�U|v�r*�؜�U�H^���vr��S~
c�\O�pr뀕����������1#w����-�4Q�v�b�8�ht�kN��,_�Q宻��:�!�hu.��xʞ�h$t�M� ��i��q�P�x#TTC�M�"H������!��Ừ��EStBY��Q	:?��kjKT��Ȫ�_�N�~�/ -t����k��c��@s��ٻ�S$�ߎ&W�0S��˝���+f��_Π�+���ɜOil���;�WM*#�jVl,d�3�n#��.����D��:��?����Y/��v�I��`N�������gR�q��Em�<*�W:����̮��:2��6���W�-��1n�U�*
��e�y�����Ms�W����~�1�~.�O�9���g ݕ���zF�l	J�h�@�#�����h�_0�����B?	G���~��y܌�f�	�qat��3R>�ñ����~$ E��b̛�� %�R��6���ɥ�1����/�T$��>�F��A��	a�D��`o�!�΃2��ƈHrY�k�����.�ěA�P.P�z`;z,(3�i��f~�>p�2Jd�uQFcV� ����H?��:-]��4�4�����[�x~�������]��Xqۍ�f*�#��m0E< 4M�p�q�l63}L��񒌺+~n��tzsM��#���,���H�ȬF9mh�����B�^|�rl&z8L|y�i>��Q}w!5oeJ&��p�U��MPsWa�/j��R�u�*��CG���f�\(&wh�y!A(�	)�45��)���>�:��ugV�L\��9��+Kb��h�e�C�%]��뤕2�`Vv^G:(3$��LCTQq�ɦ�*�����!>�O�^���"Z!�h�K[ �Æ�,׶��+$	6v�� ��
�G9�ętƃ��eW��T��f�.l�5z`�܏�K	G�p@�	%�ݘ=�p���|.C�<X�_d]$5����Q����>���}B�Q,�!x�y2f@���:� 6�5OXn���	�KI�鿁2��/��H��G`�޲�����t�:0��o+pw��X��ol�5�?t�v�l-�A���;~;��Wj�����W��_��0�����(B)��"�D(ջg+늍q�Ɠ��?�2`���A56n�����Q~?K�f��c�� n��힡��=K6�%)�k&yK*9˶j�%��r�Fb�rľ�p��`���
mٯ ȬD����*�U�wQ��gQ��"ZO<d׍<��KI'�EP|WTxm<}�#�O�*T�٘��P��[���y|���bN !X��ՌwFMa��u�z�s��jlb��ί�X��%��j��8!�m�.ߥ�՝��<uyt�5�'����h���ɭm�xЎ��l�Ѳ/���j�i�K�L����hr����5k!�0�V���A��_�y�Za��1��;C[ U/��CB�B���<7�G��t�O�Y���_�|���am��bp����&����䋺fN��rsC��S��̶tP.�K�z	�|�I���� j�:T��2g��-G`mi����YkL&����1�U��26���\�8�NZ�j�į��­Ê��j`�!j�cÂ�BO
���!u�[�k�� ���-� ����C�n��z���(pwĶ׵�K�ND�ek+� >����Cs��#���=�$�v��-4�y��+pSgbf��H���HZ�kؤo:�R.��̅v�ϕ�Bg�1���@�뚿��LAZ6"���vB�OA옢
�uX�ߠYM*z�^A�� �
�z��$�M7۾������;�(�\qN������HK�����L���dn(�b�4'V����8l
�j�t�X��Ș%6�!���������B��u�%[��8�5�&x�M��8�8w�}�.F�#��&EO�BNa#��w`���TU�5�I�X�g3$	d��_Њ8�QnM���A5P�JQX��mI���pY�.R*@�U�����M�+�.�lHy|�)�K�����?�*헞�|���D�Ml��o�B�5�[{�K��I+�b�#��]��,�Ɛ&t2~�a/w�61�
�l�#����?	�բ�F��-�-��F�s���ɥ��X��x���g߲`&	-�<O{v/Ɣr���L�D�����I#w�l��߭HB���_zÜ�6�Ԡ��AV��3�+�p��-��d��r�;���3��:����^Ē�o��0I\�y�W�~�Ȕ��O5�G�^�w�,�����6�.��Ň��s�u�y�Y[�PT��Tn�V^тA1�Ψ��
���H��i�Р�̓��aWH��5�N�����J:Kxt=LU|�Ig���uJ�VC��8���{���^b��%s�v��	��ԛ_�m���Xc��5�}w�.��Y*}#��h��Sf;�]����=��!;6J�I���X���)$�1�C� 2'5�J!~�BYX�fm�z."�[�%AR��H�BV�+d*u�p�\�;����m�ω)�2��zpܩQ��^�.���d�Ni��@N�G���SI��������g���#��B��N_���0G���$9��:qj�5t�rxY�
����������v��D�%I�Sۯ`,!�p�A� �L	%bp-C���Ls�n���Ħ!��G��"3�l��>�Z��VŃ��
�j��ϣ�6��M�ݖ	o��k�0�>ީ��-����k��ӷ�1 �>5�{�J�Fj�p�W��Lp�[�2���*�������l�3'�m����%L)��6�9�ůk��h�.!�xb�Q��Ý-�=�ַYi���w����I?uR���>����Dؔv�Cs�_ģ�}�M{�k�/se�N�������$�Gg�:�z�5w�}J@s��֧���x�,� [.�$���`)�.�lr=Z̈Ac*������	Ndċfb_�\א��Y���V2��'�ƏuH/�Ty��\�pB��7��|���%K���n����i�L&�|ǳ�K���&��^[�����!�D��`gI��&�W8h���B�z`�X�T�T�|v��3�� =2l������ג5rhBb*(A���GF��Ѵ@��!���Tb_x��f��6t���j�����UrB��|�3�P��Kz:1�ʞ6� F���i���l��u�7�����Җ�
Oq��p��n#X���:\�D��l�_&��3L#AAQe����F=2B(�>����W�)t��EN�g�r5 �̸(2(ԍߋ�lVL�9��7�88��h	��Rc�N����!����w���K�}J%ȼ��SkՌ���X�$F�������Q�!
�[#�
�Vͼ�XP)ci�"ٿ��-uIp�M�j|��L�,N�GG����,�"m���Хi� /�	�vm���!�V������f��L^*��=����qR���_78���\�Ov�,NR�t����4M�j�$Ӎ�X˶�Z�1�XK��>��B��9O0��<��<��j��sK����L��}�?O��ݱ��j� g>�� �h�h.4ED�O
��ϝ�D� ��!�����<�G�M����v���qm�;��T�>�8�5)h����f{ �)�w&�Up�{��Q�G����/��w��27A,O-�S��6�ѵ�6���XiS늲��f{�O1*k�*��7�љm���Ⱦ8���!V)�L >��;.Q�+�)��D\��CU�|J�J���
���J���]��?.�g�}�=�oYI�׬�~��7�5х�$U���AűO�@#/���'|��mY+�ڂ�{dǆلUγ�LV���i΂H�N4�Υ&9�`^	/S=4����������4��1'�ZJ��י�6��]���Al$`�f��+�,�@X�? ��D$T�A;0Ů��KEl����X����I�ie�{���d�NT���SI��V,ZuI;)>h���[���{�:�u��8=aD��+;)�ڈu(���HF�X|����ӫ�m�@J78NxQ�a�=�sreN�$��,��J;�q>Q�u�m��<9��O���W%�|l�5nuCy�3ծ}[�6�L�%�p�2���8kg�����,X����x��J��w)��mi���$h��!��
����4N�$CK��X�Ǌt��,WT����w�vj�>P���?T=�Ng��$V�����̙ν�)j�|i*!�W���e>q�?tO3`�	 �!^I�-y�q�����O��/ACO���c#�D=�b%����6t���d!O!�>�`
X������)њ����D#L�5�TN����.���Mܙ�!g���[$g�M����]�<����D@T2� M�zT��-�|�K���d�w&�|!�퍣a�/5���En6��[�%�<�l\}	ֺ*gS��,{s��G���6�ш�O�U���N�^�e0�7��V��2<��L��Uu[죔�`I�ws=Zŭ4�E-��a{M-y�L&�a��a�,��.�|x�s�܉�A�J{�]hd��O����h� )ܾL`��S_:� Nܬ�!){���y 	L,������L�!�k�р�2+_�|mݿ�� h�h�_�K�Iz�=��^��E5<�����X�r��S1�[�͵9�OQZ�p�M���R�M��?H��)��|v��f�jb�/��Tk&c�ŧ&��w��[�4j��ƨ# +kro&w��]UJ��c�%8������k�?<H�:̘�#�X�S����t�O��d?&)����C�d
D�z橗�b��b̄��$)[��w,����o4a���NT�69�Z������/S������Omn�ǟ�|��s�����Tԕ-PN6c������K��~���;5�L����xo Ho�^�"j(83>����r��Y,�EH��h�3g8�6c��T��RW��U|�a�:�\Q.g�ى�a�N
�.	�����)[�o�u����k➰�y1����̢bJma :�� .�� �l�wE2e������|d��G�b�ls��S��`�KV�.bNt^ڼ��q���ׅ ���L'�\s�hu��B-����T�"���=�B�D����McX-����®�����+�_��E�wp$��,��Y�L>S�g�9$�f������V!�Ԟȳ�yU��p�j���Lw�!~`���]EM�����+'xpĨ��C]�7'՝��׺�\ˎ��m�~J���;J�y�E�@��m`������sd���e�_����^Z�7Ro�.O�}���^�o��󡈽�,���I��|T�;�S]c��uϵ��[���ը�ٲ?HT��إ��d��#�j�E�%R�q֏��Ӈ���J�QD�Ӡm��,��8��7k��O�m�Sbɨ�X�y��~��3c1"�䶭EuQQ�%&��i-�U��ϙ����Q��pJ�m�QP��C!ҭ˜��sV讹�:4	����Әt��p��^����������������"�a��h�}��!��U���#Fࢭ�gr��~�� 7m(<O<_��Y�g���}"7��~w/���G�Y�ZS-��Cb��9�v�k ��"��J�CO�j����@�:��s(��d>��?��$�����lt �M�{���Z�.��B�x	��/Z���~.5�d���E�kp.�~n4e)�W̠�`� 4c�=�l�f(�@�d~ͤ�W�N����β[*��7�``�>���/I�y#�}��&��d"��qx���2?z�c��\"+R���h�Pӄ��x��'��E��m'9?���1�\qݮ8U[f�ٷ��Z���,�B�x�Q���]F�qV�2�K����Cii6�|�{�7O�}+̂�\���냹;�n���Ff�����6�Kf#��*\�I�/ ~�p�U���!��2�j�{�+Af�����꡽�n�� |n�&��LJ���@�ch=�J���N�-nјb$ʊq�_�X)эzO=��$J�vi�/��7X���7���mYOO��4]�Ң�Ns8��n��ѩJG}M!��s�P7���FLTF��P>�\`y��;ՙ�FS�k����-*�:t�X:��a�R�"��u������`�]?�de�^�z7�TK-���ޙ�D9���1�!����%�oM�h�6m 4�s�2�Զ�����o젦2/����]	�krx`�v�o�O�p�Gk�șw���}�Ing��,�t�w�.�h~��E���$U�
�N�ROT�
v�uI~�B��z%����3a��M3%�.L]n[��J���ʥi��:Ԙf�r�H]�{���UX^��������i���@׀1�h�=dW~n,�ëi���u2°-�'4Y�����Z���@y!��^�^?�.�?�gZu�jm�V�����q�a�S+ ���WD��?ˤ���/�lA�&jIG��bp�%��(��K��=]�Nօn�?��d��>p2���ӨMߤ�8�K:�
��l,��H��u�N��~�`.\S�

�� �7^c@�y3�Cp��@���j"���XT+�ʕ���Lʄ'T�I>�t�ze;��$j���=�K!��e�tW�%�F�0�:	(_<�a��kҜ���k�r�l/��aP�����u��;�Vx��x�UO��{8�B���]{=� ����%�;��e>�#�t����DU�2���(ܳQ�,��a,�w�.9��1#$1K�3�J�iܨ��Y3EpT��	T�2����0��5�^@�ȧ��3��}׺FF�F��aѸ)��+&�$��C�y��e���_Hk'�<�6�%�ȃHf�����0 ݤ�Q]�_a�E��e�"���Őa�~;����+TZ��KЪ�b2�g5�����[*A��lf��Y�i�io�~�ÆȣCJ���dH13x^��@��~p`#�F�}Kî���k�O�R|�+��f�G���gaUX($�0��(�_o;�qbN
����\���7�QĶ/Q�qp؂Tڕp N��́ �a�<�8�����6���?�f��bN��i�(4 %�G�U�?�j���,�a���T�����r��Z������`⻘Xo�[!�.�(zn���^��&
nD�>R�є�i0��_0UFt+B���=�3�pޅ��$���H��v��9��;[��k�Qo	i�����1��&�r�Z�������Rׂe�h�+{��@�11U�����^u��7�h�K9��ޛQl�L|���`f�3[�;½����7B�z�3N����T�5����l�G~^o�m��2� 7����Q�,{�[�����nv���4W��<��Yl����:����&��b6X��}Q t4+dv�g�H����%5VB���ӄ����Atd��(���s�u�o�#ۆ�$:��n��Z���v��2��m���3�yu�N�Qd���F�2D�u �Pl�A��i-�:��x���amQ�O0�L�o�����U�_IKT�8�̏L6ii)~�[�[2R�@ȕ����s��>���N1�E�D���%+T��ͪ\"�/��أ]��	Iq����As?��zo���E�����K��@wϯ?m!���u��a3qH�#/=1�������#��dK��C�y}��d0D;_Ҵrjn_�N�?�2*���=,���)��i�\�_�v푾�U��gՍ�{��+��=j��j�;�gv]�|��ii���x;	B(�%#w�ޔ
N3&�����)?�:<^�<����Y�m��[8�(�r����3�#YP!n�Vvø1f� ���%�
1_G���j��0�M=��?���\�UN��}��ֵ7�;��l�0ZY�!�O�X\&��ҪK*��j|MT:����tE➖�Ǹ�p C�R�`B���2����]�tɘ���n�c�0�[հ���5�|������c����^"�8�j�1�� >؎04��n�K�
_��1�F�c%�(劆�W�����q�+���9]���]�O��M%�?��`�0���'�@��~y; _K̎�_�cr�['�E$�i�`�^�g"�g��&_=پ0]]��Zݯ&��Ԕ���[��*����^Ү�.f�_<�p����%���)����
��O^���Ob���\$R�Y�i��O_��*�E�^SXS��#w�ɇ1�0�o��Y�0�o�}<��*�y�|�y�Ӈ����O���!�WY!�K�
K�m}m��ANDNq�Īi�{��i�A�7y]���3�b�P^v���b���g)·����E<t~,q�d�=�U�l�j��@G���2W4����K"�wx�`��u�Y9����{=���+L"�[Lf�8���~r�s��p���C��lnyn���:�m��J��ܮz|�ˋ�5����q�^��M��[�ۂ~$�nx�[�	��T-����� 3�E�T�&����{�=�w�,j�*�Q��ͼ��򣛯E3���LS�w�fn�D���-O���~u�OTl ���q�P{f��*�����Z��eR�j�;72p�V*"���xK��Dz�}�z�v00��6�3C���OW��5%�kP��gqE��������b��~�a�7h^M��j�{��Ņ���Alg���x�J��v�EL�-��0M����f�Z�HVH�͉��64�44@}߉�E�-�mG�G+�n��G�_�m+�,�R&�
fHSf2�Ǵ�t�t�:K����٠�_��NN��D��3��g��L��V,<CpI���V�z����D)���*Ic?�p|�`���~z�F�0( ��?[��T�+@�-Պ48suXL3�fœ��#I[��`9�a��Hp�N�p�ـ�"��ap��i?���K��~͐��\�hK��X���sw%���DN���15�&�ڤH��k,Q��T���U?u~�G%ۓN�!(�mT퀟_i������ު�lrH$L��hO����ރ�A��%?e��*�C���k>�7�C}O�BΣ�"��e�g��_����۠��Gl:�x�q�A׆��ԐK����2�1�1���{��{�*2\r`�'�)1kV��+��bv(�?���G ��,�4K���{���~���<:+��0<�Z���gĦ�J���$eU ��(OV��+�����Ĝ��o�!��L��X�u�bt���"!ѽ�Ii�����6��9
D��5Ǽev��WӋQ���ߦpb���D�0�q�6�h��l�m���a��b����I�+�"��7�)2
*3Y��X+�c^#�;Aܬp�X���������JO���HE�g����;R�2)��w��Y�zM�0��|��Ђ��rCM�����[w��.������[��A�e.�@i{�Χ~M��R�S �M�b*8�<�XFݘ�����JC�󟰎�O�j\��֨R׸�k0���K�,&�"͚�>�t�|�&�e��W�n�U�F�|k�Ǿ�k��0��9������o���fa�y�h�e��O2�M�����n8��10]�V��2�JB�tr�y:0���s���%��"%�P��7ccȤ曪ּ�5'���肕��s�x����ԗ�D�r;��D�����wl,��R�T$f63U�aM��1������_Um�r��!.���Ӛ�^�3�z!��q��
Wr�nV���o������e,� �z-�y�'&L�y�oUq3��.8�=W�o�zT^�\D1>~��C1Vڶ|$N}���R�V����W��"�"�b('���c����%HP�uQ�5�����^8�ɽu�F�3X��������oX��:,����~ϩ�GQ���W2^��!>6Ln�#�z���44���V������=ܪ,GxX�<�����[H�Xٕ;V�E�\۩&W�Y�RM[_=��[��΢e:��;6��T���ό�=�d�mL��K4��5�l������~f��>X��~������:�ߩ��W��6:�I0�i(y^Yn��R�_�h^&�d�����~�q* �����=�b@������1U���k��k�����}�XKF�ژ�V�E$m�U��-ZBS�P���;r�%��_j���Kop�5[Ї����Vm����:�3� 
������8����"z�\���j��+�_�mR)*c��P���n�R%����le�+|�iQc�L�,���Y�H���0�'�;�@S<d�P;�G��������B��tF��l�.�J�%s��M�ˀ�z����Z��%����9n����[���To2xQh�4�7�����5)�i������g�J(˗D1ALD��dLjd	�<Dž�� �R	l9��D�L�����k��P�fvՆX24���1����;~)\o����GlpF���0s��L�^����8�v�sݐ��:>I =�`�rEg�����|[�S��'��6�������&0�c�(����G�1!w�	���P��Q�����P��t�3���ν�Cr�x�v�il��<���6
&A�T�����M.�9o&L4LO�4��Gj:���]�)�=��C)��Bq�(��}U�?Aڮ�9� 2�+�X�EVh9(�;N���X��g����N#X��CKb^V�}#T�nN�g5�ө*W�H��-�m4���r�|�rGv	��kii��4eMʳ|����ƭb^��k(�\��ǫ>���T0�{�s(]��ئ�/�sk�����O����9F�)�pv�g?���Y��'�`i�� ��aUQ���D�eY�a�j�~���1�c��d��h���&���/�Z��p�]<�M1�~�Lڨ��j�Rp_�pn�z����|~�j��;l'�h&��� Bo���޻�T��ܕ���`K[U彴�=]��g�T�
P��X���nSVp�T�[��[`'xv#�JL�c]_{�'�SpL-7Fa������5�Z2�H�y�A�{0/����~2��7��
͞(���������|����:�E?x��s�1Ț�´������;�~��J��sG�j����#�?���D�D9�~�U�(�*ڂ;�,餗�,ǌ8����N��-Jb��!�@�B��a)g�Z<쬻��{iU��D��3�pK�����=[~q7�t��$	n��xɖ���'��#?=�T�=�������E�:X�/�;���\})�(Jډ�RR���Jt�H��`��4���(�"4�L����KH�h8��{���R�55֖��Ikzm�ɽ��/5Z��BR�Dkrش�1N�g��ؕ$�}�ψ��AP���%��T���OA�3b���A��W-�%<ih,�W�VP.�UvR.�ۇ;�R��ߎ�+j��pe��WYb�lyE�nҷcF20�'�D.�UBz�ޒh+n����I�@kq�[��_�[% s8b�v��r"�Y�i7z���3�����!<��5s+�z�����ǹ*�:={����R�+�F���9�EX�6e�ZS�W\̈"}�k�4�E����D�1�5��a
d�F}p�f�׍p�BS����Z����^���֯>�A��>NUk�ר����,�Z��A��fZ�R�"ܵ����E������{�*���mNQ����߆M%�]h��l2�kY��-u�V�k�2�RLwV�ȧi%�5��>'�#0��=��;�O����$l�b?i�4�����|�_���hóxy��E��u_}ں�fO�-��]�G�5��!]b���[��2���F�����U�Nk��y�D+��t�T1��s0�V 5��1T�������yҍޑ�M�h��aBH���jH	c%O����V�5�J:��2e��V����ڗ%�^�r@��;z���Wo�8�TA�"ы ٷz/���[�X^M�tT�� �I�ǽk2��X]
�����'4�ޙC�!%z��!����PpRf�)�>����J�Q����b5��M��O��D0�����B%�#���9�m"��h졑8>��#�t����ʞ@��6{��Bת$/< G7(%5xmt~�c��>�:;�6t;oļ�?��v���ŚH�����0{	X�h@�H��&�`b��oC�*���E���D9~8��}Z�����{�q:��������
��O�z|�[�6��,)�Y��UYqi�����M�9�R�~�r�E^ɸ'-�
�+�3:W��9���U}��U�8S��2���#T���F��w�1/����W����s}�Y��OZdͦ���rJ�$�jI���C�4
�+��W��K�TF"�@���=�W�+��Vq7ҾUj�����!�#��9א%>Y���w3s����88'��#=��q6��O 7䣇!���sɞ����k�
��L� MO��R�r�ڤW���Y󛶡&�rs���̍zx�e�_Q!��Q� 	���Y��:5HR]cc|R&ER�C$��~@ҖV���9�)�q5�7���������|!1?�;�v"3����$�\b��C����r�j	�)b�d��Bm��y���\�} >,i/���q��bw%�߬���X��o�7���:N/�l"��$X�?M⻷��C�P7!�ɲ1Kݭ(B�Z�� Δ�Y��C����n���ڣ��ȸj9�E�W;�����s��D�/���� 7�z=�PL��OfWѣ�'x0j����|���!]{ҞG�+��������8���3�V8��+@�]�uQ�q�<�l�,s��p�tiU�W'�BL,� ��efA_Vs���W�"��y��@�@�I��Q�ۨ�Tg��q����!&�Wٷ
�A��V!�Ϩ�f˳2��s)�
y��r֝����� �wJM��Տ��e�¼�s�v�x�x�f�z?��;ΰ͠{��,6�ѣ�g��y�O�,���f4ůnf����>L6��D���f`7�#V��b/xڿ��@���c��8o{�+8�J���?*�
5ٹ!�{�oY&;D3q���_eU�&�i�D)�T�^t*�ZR��wq��duD�@ZO�}�%�F��E�B2#���e�j���J��X�Hf蔌A�t���8��S��U�D��̅r���Ř���0�t]9�ѓӸ1P&�A�H�!X��;��_=֪~/�;�E-'N�s2�
i�K-I����8t�#%;$�gގ*=ƋɆ�҅�3�Gn
�ܢןfS0�Pk~0����hu����F{��s��<�ۍg.��K��0����(,�a/��X�0:��@j�)q����Նŋ�P��ן��b*����_�|����1�7�E�:�O�	'��g��Յ(~(?(*+�N.䋪F0
�d�-��[ms��F^��iU^�R��N��SW��S�I�yآ�XXW�OZq��3SQuTZK�VM����-���*���*��N��؀q�\�rO��U��~�"��藇�9�v�#5`N�Ɍ%��l��9'��>�ö�@њ�~;�">W�#z��%HO��#�72S��H"LվD�� ���~��>���̂a��bm<�N���&��:l���r2"_�?�y�S�x UW���1+��ۙ�v��B��������o_*�ȂZ�y�O^�E&�,҆W�F�__�Y�n%��>��"RoiY;��?��5@�1I�4e�Af�@��;��f�R��}��c����ǚ\[���2G�X��$L�rѻ�S>�N�T�(��OE�fÎ������̎3���3R��:N(<x�.o'������48��:N3��z��F���p���������.2;��a^�WHD+�2�aFm�vgϝ���C-��?�k\��IW�-N��%쩺����3c�ʆX÷��� 4���Hed/��5R�xMk��`V�h`ّދ2�ě��B.K.��P*ܘ���E���I��Ѻ\�Z,�&OE�ӯ���@��A��
��g���)[65sN��x!>u�!Nۓ�*�ң��&��_�j�V.g�U_l���.�[~m �(8�=�����$�0/���M;M����y��*-T����?�/�����f�9$�=��J�d\��ּ]�X��*F[8�4{Ap?;x�&�^Y�E��_Zi�s!��gh��v��O5C�<�ʰ߽YfCf��D��
fd�	������״�SA_!g�杏�yE1��.HM��֏_gsXֱZ�A2{�8|��\+C`N緢[�(�:���;�\Q7Y\c��ꅑ���j�{��`Ue)[n�끢B4���o/��W�K���yJ`�iP���!$M�Ra*���\ҍ3A�"���u�}����mt��4���̆%�b��_\2:�%�m9�Zd�g��v�GNo�'�sf�;pf�s�l�n!����̯�K����X��֤�T�#�z�V�Ֆ*8މv�FK&OdRT��
���H��q4��D�+���Yv�Y��m�ү���Y ��r�~(,�h>��NCf�8~���gl����\0y���y_)p!l�  �͑�+�
����2��nL�H��(�1�a��_HQL��q���LwKc�mAYv�Q"RW��*�v�b`�����{������ǚ^!ɑIN����[G����[32ϯ\]z�)�+��s]�^��L��kܢ�Ա�B�s�X� �W��{���f��\;���,j�0xJo�C�(���$+��ʭ�1z�p�����]�
�Nf���V�D�:���IJ{G���m
��"�wJ�FD��̀!f#��V/ �/)pw�{��:����v1㌀�p�λ/�o��M+���b���t�2�p��L�%8]q��w�UEW�;�t��'�-��O|������D���v�p�?��
>�l�N����K~=�m�x�����ۓ�h��S�A�J���@�W��j8ם�zK����U�>-=��9Yw�v�����c�ׄ�]��g_Y'6�}��&
V4� gE'�5IKv������'m��<��Ahp$�t{Z�֠�5 ��/L�f���y�������Pө���p��A*q����ݨ��*��k�O��h���J58^6e%SgDRߦ�0��w=��!��Ģ8��:�5Z�By�<8誅���*?H�7�r�V[�/��Ɯ48������g$#�3�SY��*�O 
q�MR������i�±/q1b�y��ﱪ�/ �X�!�f���ځ緄������3�2V����^���4w0ԬI<���PI��X:���g;4��v�T�C�=����~\#*<s�U"g�-w���h���1S��2��TTm}���Eq	��)f�^��_I�T�r���ߥP������7�Mpҟ%�y*g	��Pt��{�y����/(U-N5a�B7�L�n˲[���2������́�,��x�ᷤ�?�]�A�;R
���]s�v��h���I��\	5%|��=�-�:oZ� a���a��(�)����z���N�'uɊKd�B�h�-�Lx�()�6IA��sj��_�r��.�n�k��;�l������u׵��B&ϛ)v ��Ӑ�lR���-�F���Ht�q٩I��"��-R���%�S�ڝX~(w^��k���؉Go�4~�a�y��V���Z�]�W������3�T2�f[�����v_��󧫟[���M��1n��E�G=P}Ԝ�%~�{���޶V�?y
��
��فk}�u�N�g�T�<^F�7���+��\:M��8�:��2o��RcNZ�ȀYϳ(��h������l��`������b�e�=z*�L� T�<!�e��X�����c�-�LU�L�"N����K~ �w�ڱT��>i�l}�L11��P��.����|�B��/gM};���g�!�qW���^ַ����.�f`����>�?-�M��Ȼ5��L 6�NA˥��P��Bbl����	�+��j,��G�z`�7[E���Ç��rs}*��XB�7�p?R��5�e�/��?}Lq�%�������ը�S	O=J��/aJ�"�VFB�ء�ˮ�d["ni�fm�����9|�E���$��u�?4_C@eTs������_ ݬ�V6����"�G�?��:��D�.��kqp��Y��V݌	��ߣ@��3M�����_0	�`����d���%����95�^K�r�,�-�(���; �T�d���w���Q��R���~G�ƝC�~�>�ھ�O�Sș&�#C����u���@cN�k�݃� �:���˟4S����x|pR2_�Qx�3�O".�[�Vi�,�4��!a�K:���Ϫ�K�#��M `s|wCf��s�{�`R~[����DzN텴t��0�����KdS!+j��0,�+~*�)@�q~���D�&)Ѩ2}_Ң���J��5��@�g�@�6ie�`��J��"�#Q:�Ԯ�(�{��Au���DR-]���7���o8�����F'�:��,��g���±�Z��z�_g�iԫ�L�x�,��'�@����U�=���GX����*�m�7.4#�W�W~-h�x��^�n�J!�/��ѹ�!) ��0q*8��Ӭ�Z��p�N�St)kOul�{,��t�U�P_�)3�ڛI`4����OL=���%=���^���WP�Y�)5�%�n~l֤�MsLN5�y�2�a^#�[�c(76e����Wğ.R5�����v@�	�ا%��ӭ��W$�~)��T���<��i6*��T�Aώ�B��\b�J��X2��P-����=xK�rs���'�5�27a2�Y�B��6�;HS$^/��wX�����^/U�����0s�Y���z˂Z�S��⑴KM �^���ʷp�=�����MH;q,����|=������>B����$�Nv@*.��fPw|qi�e4B�����p����7��VEK�O����]#����7y{���x�bA�WI�413}��2yK@�����۰&�Un���7�A��+���-s
xL˯8�%����H�x���_�cpA���A�Қyu�EN'��&�aC�V���/F�Ķ���l���w���isd�����n�M`���c *1�Rz2^����W��{���XӮ�H_(I����n�������2ö��CKN���G��|Ԥ���2кN�s{����E������7�O^���l���(����!��~�,��3j]�<�2��-�ÔI#.���^ ?��*i\�X��N��
"ފ���>I�id���=�ۗs�u`��N)���j�mjXA�yԥG6I�ű5���a���[>���x�v��E[�U3�-�z%w�P`��S��~+���vbuShqHǵ#R�9�W3��WO]~�3���f�a1�1��k5���_Y�|� FX�氒_W4��yvv����j��2a�G|�L���ը#4�ۜa�"��BM?+%�ɠ���R"���SI|���_;��6�^k��;�o�ݜJq�d������N�g���\T�7�j��2&` I��.��ɜ��`�$I�/W�zi�e�n�s��J���νXU$�!����7��[9��Z��Aq��S;�RZa�)��cM��M��Ĵ�9tL
j���H3Rh���c�f��VO�w�\H� ��Rq�����J(��%učo��g<[ȕ�R5e:�	ġ�ys���+]�_�@�ƨ�/��&��[��B����$/Ng~NSqC�XsX��"��\/a8w$��	l��%���x��Bf^%���<���B��҆�3odaS���iᰙ�F{��f�]�����d�<�{�͠)F?�"����v�T�"qG'�k�¢���s+�x�p^��?өr"8��!���y�.��^)��
���a~�<��Th�3d��u��jF7{|,=m
�|`��{k:-�,�Q��P�V�XX�ўSSd�#(��F"��"��D���)�)�VT�?�_�G�,M}����t\M���42"���peh9�CFu��ʡ�/��]#��8ѷ��������H�:�P�^빃5c�J̈́a������]OZ!�K��5��N��m4����b�;�Zu�A9��k��KB��w�l<���
V%uM��P#�~�>:��%���F��5dgˇ�g�[�7�!(|*��;�Ն�t�5WnFmcs;�����8`FdAV�Y ���R��qgS��B�F쇣��$�e/`S/a֘г+�a���Q�L�݆��
����pA�0{L��n@MqI�	�R�����	�{�	�%�<��-�����e>�6Vܠ*9x��+ʷ_���u&��M����>��qh�c�������D��Oo.��G?d��Tʁ���h��~y%$�E�%Ra�@[�`��~��,������������ԏ�/�c��\����0f6�ȒT�|"�
��i��Ú���EO7Nv��,�X�{����]�?�����jHz#�T~ �� �gGF�e*��i��N�ǥ�*FY1'n]��떹Ҭy%1u[z��т���X�������:�3�Π37^�U$T/��.M�o��S��*)�+�ԗ.��J�7)`3v;`�pS�N�4�<A�h>���3�t��r�@��r���W2e!��f�So�|�/В��Lބ$[|�z�g<�GGf�����K�$�^����n:����Ι�_�YN$�xh�}�#B��h����R�n{��Ц���ߓ!�|'�ăA��Oo����y>�3?g��A��M��x����I���2�y�H��߅�fv�2̂mq����co`�H�-��(V�פ_y����_�v���=}r����M�P��9�ů�����h�/�;��-%�����ouP�:������]�!5�����V�D������z�����8��ק<��g���� ��֘o��A��G��zʥ�s��C�$����<J��i��#�ҷ��ؖi,�+���H
@y9�W�g��z	�/�}�w����"_�몇c	����إ�Ҏ�s�^���E�䨇���[�Փš�v���dз��m����e�FU)�ݬy!��Kf��F�	��Cq}������J�k�y?�3�:s���\:O��1�|�❌��a��?��l�ĺ#���i��w��;��b���M��'��K�ɹnDV*�6�����ܘ4�D+�+�V�:)+��C���"-�P��kz��F�0���Tq��(H��z�|��������Sw�ދ�J�M��)q7m� .�>nwd��<��`k%.�i��ǎÝ��IRpbv3q~����?D!�yH>�5¡��`^#�i����)
�bm��ᯢQ}��3|�D>t�>�AY����O
2[�q��>��5,�h�6��0����L����'J5PE��տ#iLG1�IPd졝�2o?�Z�{B��*�%�#AGC���z����c�]O0�<Qt_M��8������c1�4zf^zW�A�S��l
,![^�����!���S����J�7�a��[& 9�z 99��s ��1B%F�=R�'����G��0�k�'|���>e��OZ{��� �`��h�C&PXi1 �0yuQ}�.Ǝ��k;R�C�ձ�ͰGG)��?[X�����}����u��<���`�{�5�T	��1�.��
"8�}m�w�-�Gd��fU�[��"lU/??rm�9��8_�&�G,Fw�
�v��J�2��,E�Z�E�� Q�X�w��7���Wa�b"ӗt�ϗ�4��U���[z��@���"�-v���|	(lR<s4��Ϋ�m�Q�D��{�.�6���mNT�s�(|���VV����b*�dpZ����Ugza�n�T9KY�q���z�g�H�!W��Lީ��[f<�7�=�6PL����(��c�R� -����M%;����]�tA!�;���xm�{{h�O"j���< �J�i�[}Q�W>Hڸ۲�)�ރ2)�l^��[$H�_wI���aо9�w$��[N���[jgw�2�R�'ش{o�3�Kp(��=�2@E8��Jbki�ࡂy��ts5o�YG��~�+�������1NqL�� ���h�:IDC4�e庐�=��G�ӕ0x���Msl;����f��_����,2��"*�U�+�E�x�1�0���dL�2���%�xѝ&d�n�z������'?u̗+�L��C��Xz�sJ%�6hN�RX����ڰ����rڿ��D"�_K��g�3�Y�6���r��%z(��P��c��,Lo�����ٕ�Oo��Ks��*BpO�*"87a��UK���O`�/jr���&�h.}=�X�cy��<�x#�����P+Q�V��s;]Ȗ`�NԦ��+t����QCq��������-��wa�� �"���~�R���s^e�X�_�w?tfZ�-N ��MXf�qnw}�@��=M<�&�=O<a����Ϋ�)��&L������7j|`]#�'aK0�(M����+t��ʿ�L��2��"�w�OO�J����Z�[��B��'��p+�F��q*Q-��hfř]��b^O��y��Y|΋MpU��l?y�a-dEb�2Zi_0��K����n�]�Q��h	�:-<4&m�D�o@�л��U��X-͖9'^aD�nN��TP�[�ڃ���/����������mtъ @`�f���F���ܮ��ԭ&�ª<b_��&޸!�Ӓj֡7�������qvMuܼ���*mE��F�2x���Z�_	E(�_K	��Wt� +]\8F���hJu�!�R|�B�rnIY�;cW8m��Gx�C�򄭛����f�g���i@�\�_��b4w��.��[>�+�_�0;j׀�fޒ�]����=��f���!�Q:�Q鬊�^��]kNz��ͦ����l,�ϝ��̎����4�ujy��}��Z\��i���"޿��)�b߈SԜ���%�g���	�n��KG$0�g߱�3��b
e� 2>��<�7�K(k.��ZV�F�&l5Q�Odq���l_/�-!i��ˡٝL䝨����S���G���KD�yYLr��I�Q����or�7�H��ף��>N�j���k�F�C�vh��YS�J^@R�r�}�0	��{���v�6f��Hy
̦ǹg��r�L57I�-�Sy~	L�s����u�	l�{@�h`鵾9�+"Hu����� �j�<��tC��֒�Y�%Q�([&�@U=�2#�ꔝF�P�s\���s�"�ͮ�.�������"Q��a���<�Jt�'is���2�e��v^�M*y�v����I���]q��9�1 <��+�S��h�#�s��5fk�S�!�6 �NKI�
�k��8�Z�fa�,�6/i��H��M���u �w�j؛i�s��)|�!L�0��y���~lS���d���������v��QT��X��U{�}�sk�������d��������'��S�h燘4:.�-���O!"�IC6��kІi��LT���.`��M`p��?,�0��G$�h�M@
��u�#܎ �*w���5�3�1a;�Į��D%NY�b�u�0���qQ}÷��ce5� ���eM��,Щg������Rh������ѝ�����ǔ����X{��7f"�z��ol�Ӡ�n82jᢊ�s{��D�~�ʐK;o�lye�C�zɡ%-����H[-)D����ǒ|����m��ľ(E&p,���ߗ9^�kn��F�8r� � ۸�,�JO�&���v��Lӹ&����2��,b�%V�o�^�X�Su$�6�~�y'S����`BU�,�.Ę�h|��e�7�ZE�Q�v��Zq�
7S��W{��|��Q�����/�j�k�������8�����b����8&�`{j8����ӝU�����ә=�H\�<�Gւ	���h
�n}|)sВoίݮ��/�!":n�yʛ��!v	��_�>9qebP:�5��I�\������n�u��*�N*R��b��xMy�M���ಙ�=z�郃N� �1���{��ܑU%��M����+�x˯���Jm����o��Q��s��1�h�}x��ҍ����<�"����Ԣ�ƭqm�9q��S&��S�����tXdߙj�8�j��FI2_��A�T%@����Tvқg�B�d�j!]BXk�ȟ9���&~�~jd3%��FI�i]�O�xgƹ���b�,}KWK�4��^DUU��j��CEߌ}v^��I?�(��4
U,s�?��q�OOzO�jI<�!�}��hxx�D>����۲Vtc~S������X&�c��vO��Y�*��3����"�x�)^~5r�d�붾��/뎝�	�0!��29itҿ*�J��DbU�ȉ\���)$���ä���=Z18�_#}_�<T'��,�q�$I,���w����0�USj.�2]�L���L%:0�=�v�4�{��4	?O7$��$X04p�s��1ɨ��>��������k�A�]w����q�_���dX(��v��I:τ_(�A�:w�3��E��(m�{�ڣDI�s�o �����y��e�ڗ�S��=�4�!���6��!, {�������N�*T>z��.,Y��V�h��
7��>�9��,���a*�6�X�������]/��� ھ�ʇ���2���F����g�e�QK�3�rw4���16)�Cj#x�RyJ/ ��WK�FYE�O��*2�q��v,E����9I�r���[e���ő��0�ʛ,��g)~V2X������n
���9���&i���u����v��q��/SO��>��I
$�~��
7jt�Cr�H���b�JGN&o�t��L�4)J�8���1A��S�Мl�B��#��:�FW7��V���|����'Z�6�H+꫾��=�ׇ��e�@���p�4�YOrjq��\�@Ɩ"Qk�٨��eі�BbM���͙+�2�k��㝇p�կw0��׭u�44PH7���Km�Pzx���C��oG;n�V�Fsp���#��7�.�˳��}��\�ttv7�H\P����0�{�wI�� ��~�����7Q�{K�.h��2*���a#�JrU��Ŀz�~�&0ZY��k��4-��5ў�\?݊�K�*>U�7�v�z�P!����[�8#ƿ��N��4�Ro=��n���}�R7��uA�H�e[�)X�BBL
�N���5������d۔d߆*�v�M��I��#�bZ_�XJ��b�j]e�j��cl�s�oz�� |�_��[o4=������\ق{��Ԕ��	���&��%�@�3������Y�޳F�� `�'��Y��TW
C�3:fY�h�AF��ػt��h0	I�Y��{S������YNh�%s�ڵw�{�6�o{	C��d3[5���h� V���$C�<�$�~�?�;�O@���D����t����+��u��Q�LӐ��a�����:�V��O�1��(^����?��+p��{��K��Y�:ɦ|y�h�OT�B;⛕5�dX����Y��J�3��Ħ�>�ė�.:�q�M�d�f,4w�C���[̗ZC�2����D_��v�����}Ʌ��|�w�_�'�1k\|�zqE�b��HQ�ś�L���cĦ �%�`�N�&�n�X��&;�!��,n�/G�����?����iǕF
��1g1�Mo:e!�!r��Ti�ȑCq<������ϱ0������]Q����<���?nQ姨�a��?��R���v��$��M��R��9:����� �x^��) ���Q��i�_���t�c���ND�,���c�F�uJ�ڋ2���g���\�h��q����'Jĥ�ߏQw���d��@	��<b�[��(1���j� q�"^+��D�Y�T�Ϋ��\�_��>���g`|�i.YEu-�Y�!$�'��Mm������7U}I���j=���QC�՜��	��s:�{��^�KG:Z����+��Pl������rS�v�RVH��5qcV�'�i^�yFdS�Q���vK[؇~���t�%,�>[��Ab�ufs����#��=�e̬���	Ĉe/A{����fX��UvҶ)�����A(=Jd�'mh�$�r�~���TN R��/�E�����-�D�2��X�����T`p�0a5��
�Z@/�$1�>�����$C2=p�B��hc�R�K�:̀�&�O��[>����`%��W���@��or�x�Z�vVXs�OiR��	�{D�b`1�>���$�����r?��7N��ԺU���f���\4H����Q�k|;U[��
x}�4t����)��>��aBF�t�LD�jo2������j�w�Ԙ���63�^O��Zqg�"��kM��`(��A';~�6z�y�4�D����L� � e���%�9&\��+�f�0�j���O�m39���;@!Xn��T~G�}F����T�tO4ܭU?��ҶH�1�=�A�(plؓHi Ly��bVX	R�s�:����Vǆ��tѐ�p�3^W���MD�τ3s��{���/�Ǻn�<�ck���j����G�)���j�>�g&�q��ߢN���7�nQ8�;�� H9U/vZɅ(�D(�n��Pg?�/;1�!o^d��F��[s�378��R�%�l�a:���7�\ �9\Y��'n��жj�������9@a��6����Y뗿���F���B��K��ؓ�x�E��v��U�򮵇���j�{�@ĶL��/>r�]���qhe��5���،,�>_rOu��XNA]�Y
ʲ���I���1X*v�Pw���9��7�����z�@*�*��`Syc�DҹF{��{�:�8�>�M_��<���8�����^������	��{uk�K�ڜ�"]���|xi�k����7�hDhc=G�����e�M��xޏT���;���<IacA �j>�Dc��բ�O��K�PO���j�g��� =d��J���{�Z�Ѻ|�-�����I�<ʇ�3~DNX1ԑi%�)�_$����)�� @!b����ދ,J�$��>�$h�hcmN�}�ʻ'J-�˦��=ʑH�57�"�����B	6�l�N��Ǧl!�Z?���L_�m�Μ�`�boŻ�ۄ�6�**)CJ��Tz^�Wl�l��m-�Q��Pm�3w,b+Z��``f�l�d9���)�|��*n�P8�. 3w��|&���MA�w�ts؉}r�Ԛ�jj3�} ~�b})l��t����,J��%���.���1�ǫ��P���`�����m��ӎu�uKq�׫�����Z������z�u��Q�i�2�;=��P$�f�ƺ���x�M�n�b̔j�7V� �w���ٮׯ�Ae�D����6ua�C��Y�k��S�J�f�{�?�R+��ʡ�]\o�ڮ:b���7I�_���#���?jd3�7�,�@	{�J�tV��:ۭ�C��Vץȝ�pB(5?�r���Y�I`V�VT���ȣ�GoG�Bx��'�3xI<,����5�@L�U���S����O="�k����K����������n��&���}EG���RN�K���v�mJ�BaS�U��'m��T���_{ԇ��]������=�[^(�!sv�4[�7O+iޮ#���@ѕ���'Z��>�0nS੯,�eC�u�r�ץ��B�t�2��/y~�N�	}����ڃU�<��p��&O�8����{<�y�s� ��
��� ���= �a�g6���u�V������4��N�T�;Y_�U�_��#ؙ�!ج^�N��\ ����8�V�N�'jl�z4~ˁ����P�2��&p&5x�PQX��å���9�N�����N��ʆ�S��( �U�r5��(�u\S�&��(���p���n�-���L�&�<�g�d�c���/��,LC��@�Ip���+�;���&o����`�f�|�Ə�p�&f��L��qB旞@Ub�o��_Es �����f�>-��U� �;��u�vLr��\�b��C,�:c%�y.�y��<'���ǅm����4J"��ā�1�X\ܳL���6u�nJ�1�����wol��¬&A�@�Vw�����j�I4�EV����N){a�D۟��%]��P��Ѻ�@(�� 5&�g�bJ	��0a�֮"�o��7�l̽8wZ�JY�.�{�g��6��|�(���C�a�^f�7R�))k~+�3�O�1~��[j���7�\�[�c��P�@'�=V���>��֒& ��g%k�<�r�z�5Zɷ�n��\@F�z_2��8�T��Z��+�!XCn��Ɖ6�+��`��@ޭ~�S��V�lU���W������桁�pg�6{R�����rx~����n��v�5޸)�Q��b�Z�/~aj�c1���U/Ѧ��|�$/Vi�h�O[;�H�gg�� ��L��N���>�h�pb'��s?�TZ��uI��cV9�A�^T�e�7�XX��vIp۰�%��	ݽo��O?k6��9n�(N�w��4NMc�½�~>�j^��d��\��P�;I|��R�c%���e��~uz}�ZѠ~u#k73�+��e�\�ri�Z�2��m�0�!m���c��~��RU�H�h�(ӟJ�-q��n��_2/)��-Sm�i�'�s�X���^�[�c���'���a���>n��]U����X m�M�?�v�h.�f����Kt �9<������m���[{��������[��J�y��:�:D�|>_M��$��x˙w�pP C�IbWQ�&��%�)�:Ih��)c�����fI,Ѯ`�w��}����1���X�р�������_{�7g���w4����n��-�6�r�/wo[��8ھ[�ڋ�ё�[a���!�#<dIЙO-��7��1gvhi�wZ�l��U�Dk�Y�y�w��qB)MzW�����g�b�=�CΚ�=X�R���Nf���Sփ��t�w(f0�9K��È��HnYî"����y��8vKHc1�(�AL�KR�=��-V�'*Q]���9��r�Xg�Z�f��߳<u�Y����I�]�������|$&��9>y�15���G�(2;���<-칇�-�����Y�̣�H࢘ᬒ- ��7���=f���)1��t���Z�zR�p�7�
�ȜV�1�z�}�Q�6܏�"������ ٟ������8�b�57
'g�u�����<>�ș��/)��K��c_p¿U������ѽ��A�O>���`ʵc��RB����f�IP�uX��4A����@Jr8��r�>.xTB)��|KK�]<H���+5g��`�����n-�fT5�ܳ��a�oW��(ѩ�/	��k���F=Ȫ�zEW�X�xi��.G)�3c�Xi!���G����&�5
� nD�^]B�y��_��^���.��S@"眅�4>�43G`I�Ա_�����QopCE_�X칠_�$a�u���&-~}	�de�����;j�)��\�p{7�̖h*�8\�焐}a�JE�?b.)2����Gt�������V .�P���o�����\-�XѶ7t�t�-e�k6��l�5�_�3~ԋ��^�2�0C\���ěY4s�qJ�DJ��,=�R7�<��.�M�Ɗ� ��4�&���y��p��6쁍��30��mNJ|���iw�V��!z�/6�w[�#j��f�
,�`c��h�}wnw���+�[�c;K-7O�J[�vt� $ �����rZ��g�`"	)"_��=�Pz?�#����7���	p��Q�kޏ9�
�C���y%[g�����]����"��CքxR��(�x��bkJ,B� m�^�x�[P�_૶�,��6�&"#�������._����L�tEm�>]5��3��*��Qz;���I�}?r��	�;!~5���gDv� 4$uQJ|�F1��^�g���܋W�Ī���vA%q��cƗ6���o5��ܐ�0��P�_��[�8�Ȁ Tc5	f�v�u��4L�9Xޞ�s{�Ց��h�Nb�M��Z����^���+[u�����s��d��7~gws�i��#�k��Y�������vA[K0��ï!o�ֲ�U@6ŵ4�A����߳5�`WS���&�����sU����n	�A&uH�q}�� �37+��ȶ0.J��NҦ{å@�G2�r��(��<ʢ4[T���_���U_ZX�����0��{O�p�={4P��xq�~�t����"��o�E��rx+�D�u�mAR�2�pZ����p��țի���~��	@Rr�v�op���W��73�*�!o�E��a���!��p��
�Y�]���_Z�QSG�:Џ�f0�����;N�S���Ӽ��@�IuE�����i]<�ϼ�$�����ʥ߬RH'B�[�$�ˬ� 9Ļ
�T'¥ϴ'Zj>��)u�g;=O�c�Kc"��$8�^��I[�vW-���h���T(|g+�H��.�����.���D?8��5m*�),r������ $����B����,�����
�1j��
�i#��E�:?B�?ʧ����_�B<�I�vt�v�e��J� ��6ç'���m��lY�7d#J�c�IS������s̲�1���@��|���7�a5�����hB}���9o�XIf]�-_(q?Bt��m�
��(�Lܽ��F-^ǣ������;�5���g�=93/Cd���
қj��r���6���N��8���A����5Ƀ�'��	S�c%��F�	lg��[������:{�o�ܺP
��,� 5U]����b��� Y��)�d`{𩔄�=�&��������U�s���4CZQO��4��_�܁ܣ��D��fH��:����)�!��=YAmSz�?��(9K �����o�rA3��p�mx��?��yG\���)���x&2�0��4��݁�^�^���^�I��ݮ��_Ӛ�f����ԣ5���!ʽ�/�%�7*�͂I!F�a��!���hx���ٖl^|u�Px�&��|E�&�󊚡�KĞ��~C�j���~?�V.��[�Ю�ct�
��P�#�y� ��T�ԉJ����'�,��wjc�y÷�9�q�Bn�^M���;W�ݼ꩖#J��.U�����<�<�E��+�.g�>A����)7�����\���3W�;73.��e�gh���O'�H`q�|g����,��H��;�%��rW\����f:�h�y�W�d���d^bE�V�q�޶��m�J�D?R[yy�L�",L��9�G^�V�l����wnT�ެ��SCkx�3�551��^��e�Tܟ��ò��ܘʴ������E��*>��,C)��"�k0��OҮ��Ϫp�����5<9�* ʠ�l��C��w��԰�o�2X-��U^�^�A�y]�����:�\��0��4�O��6n�V�w�"	f #g��JV;� ���lIM'��"&f�|k�%Ob���X�=�¼��nu�rJ��%,���J�x�
_b�ι���J��Vm{�4w_���(̂h��P ?Ր���;��*�?慇��>kv��@��D�uÇe
+�a�)}�̕�n�pH����J9"�o\����,mU�jJ���.��ilm� �1���x����
��g���~�$�(�Yv���Z�#RG�J�/?3�t�2�n�xf����F�B�}Dv1�,�*�|�g;�
������e��beh�&8P���U�@K�ҭ�/�Sda�L�K�[%	߆J^K ��+��}0�X��>�3y:^��}�Ǐ+�r2)-X��۱�j�
"Q5g�C�(���G,"��ZI�J��]83q�)���^��!��u���3L�^R���p�=�+Z�B0�^nUk?k��-6�F�$a�w�k�3��匒J*��V�Ɉ�-�6@�I�*���m�'��^�?:Zm�V���b®�r��/��9q�o����hQ��Of\���S|Jᡡ�4��PhR��<�����O�ջ��0�0��Z�@(������oLsY���}��A$����l�68|mk�JP�������AQ#���aZ�3��}�EX�V��+�ͮ�Hd�ݮ]�^]�5��x+Q���P_p�҈�QϟR�؜�c�BZ��ħ���Z�?n��\1z�������26���O?������9"ކ�d�b�ݾ���j_� �<�Ȱo�=�fpq)�ǩu��ܶ�{C��	⁲P�J�M����1�бB� 7y8�r�1ӂ�Ɍ�"�{�1B��!䝤��"т���>�^1��ؕb��JQt)�h<s��k�
A�!�J|$Wu�3�P�I�c	<�^<�R���u	6DŻi�;rv��[Q��5��p]��}$bZ��µX��gĒ� ��+�;��
Ġ2�R�R����NY`���'gF�/���x7ⷢ������3�e�����vw�j�6���]�W�O��H�w�?z��9��qd5�rU ����Ǜ߆��� [���P����|���`���x��}U��TCUҭ$�RwS�r�!�mT*�
����NHS��3
+a�쒌P�����T-��D�l���e��}:�u �4�/Zl�pL�s.\J�>��)}�������03���0C�M���3��0�N��x8��KpT������{T��?7I���/��w��ÁG0�(|��1�N�V���U@���{l���:��l���gW�g�����D���^-;� (pK��1�􎼨dlH���l[ �6�VQ��?��fs�����c8�񪪈I
:��n��붵�C��HQD]6�lM������/3,�����tK�{�;��@x=�k�3�+c�>I��"G/W��@<� Jo��}rq���D����Qb$B� �̤�&0o�!{��r��7��!7ʽ�×��ӗ���L��F*i�ԏO�
@;��TV���>gl!|�c[ �bi�:+��є<Sv]���r[��e�-�x	@�3SL���+�Y�T����ވ^�ש>�٭I	�Ϥ�-��ڪB�K3O���tQE��
��c��)��k����S.�4�\�� {�N�OSr��4T��>k~/'��#���	B]���-�]�BB��y�\��$!L!�˔zL�*�������%E[^�4��ݡ��+/(cU|��!��0�
Z*��Ɔwc�MA�ӟ`el!\��W�����9��z��y?��Q�կ⌂�	��P���Y/���Cv"e�*�[`��ĹT��-j���t�7�x�`I@��L�I�s1��>s�������:?lX�a%�v������$aj���r��^3�mڀ�3n�]�+��]��R�J�����Mt����� �]��U�]�8��|�HE�
�"��?���~�̈́�'}�����z̋��+�����mHV��U/����3#ą��^}t����I
'J����"����*��R,yrsH�ɧ��Kvﵢp~Kv�|I��xku
�OP�D��5�\|���nY,c����.��qi �9B#�S��u#᭡�U�ݶ�l�~}�XW鴂'iE=~/��a��r�+`n�@��v?۷�4Fjx�hk�>�Y	�R��v��by�"����M0����� wP�����]F���u�3mj,��q~)��u�9�#��i�Ɂw}�x�j$��tCU�h�f�
.��Q�`>S+~�7@�A�l:d@���KA!Ƀ��t��X�'^����K|���H�gTD�L�voT L��V3�N��_��)S5���ONLŕz��q��s��D�Әq/\5Rϭnw����0<0�@.���$[)�'XWl�8\�+��وu��6g���Vy4�������M�L`�������̤��A?͆5.&�2L-i�fx����xg����*sH^���5��ym�mf&��׭L9>�Iy_qϙC���V�C(�R�=���Y/��J�qf��#���!8��DS|#%q���k��庻vhf�Mä��D�EZ�ϰ���P��l�Vy[��!ׂ�>�~����^���
��yO���0ʬ��$ئ��{Y�[W���-��>��s� ɡA_�4I�9B
�^r1�z	�3�kG�]�'+Y���">�o`n���_�Cm].�0r����G����Hy�.l���%�++�l�M��AM����8r2W���"c1��j�U]8�x?ʘ�_*6�-v�}��f@�2s�E�-��l�ڭ{�"��n��h�˵�p��O��8�-Î�WW^��vӛ!<�)���o��#5�x��of�s�<�gB`�}`����E�i��Q9���\�}ΩױO^-䏽�^a�<��'Wkq50‎���*5�M���?sX�A�j������	z��4^j$r��W�vOk9�!q�z�Ϛ_{(�k�� ��,��߽/�{�Eg�0��WǾ
r�T�yj.S��K��o��p�ݒ�5�8�bmƮ����� �>���P��5 ��J4Z��|���E�׃��#T����_^�1K��@r|RK�*J����R��y@X���L:���@!��{�t"O�o�������������r+���4J���ԡ�Zy�$r#	�2p{׊�T,.x� mW��i��9�{>n�* �G99&q���+�X4Xؘc���.o�[��%mDH�.X���fR����0'g,+�Po?(`�7x3Tʰ�54I���A�o�s��NF^B܊���:�zoTޠ�������
{x�3�\xY�{�����rY�;e ���f'
�`�q��0U7��c=��e4CiH"?ȊYNAVƉ���|�&E|��',<G(#S��|)~U"�Bc�f/3F{�yeA5�zG��D�Ȏ%m�]�t@74B{zDJ�A�8�Ʈ������_�`�AeP�8*W� �x�)(qQ����o�S� ^��û���{�K�7�e�q�Rs����ƵMk��M��2�#dۗ?I��Ӟ��p�s��$-��QT���|�i�� ��8�y��(�B��O_n�}z�
�e�'�S`�`4�;lcwh�ġ�J�o�rD��C���� �S�s&X���o�'�Ə��X��I7T�4�@(�DP����ꤘdE�y5K�y�]s����g�?op��E<��$�
�su�c��s���^�j�d	k+aZD#��U��hbP�+�'!���z�?K�VD�p����}�l��'w�\��E,b8Z2�t�.s��{���v�P�>�?R!�C8V��'��w/���򋺼d��0�F�0���;�������I~�倳TfK[z-�nnT��铍�� �H���+P�銱�f[�)`�/3��y�Gb�K$����ظ>1�/�*P;� zQ�L��/,�#I\����tnLh8y��NT���5B���cW���I$�T�:��J=�c�	om�u�W���/ �<
�'��/z�n��Т�M���Ѻ
�#=�.�ݓt��aw�sܧ�.�������a_6�� �怏���@��x�k��
��,K�7╳˵��+ B�u��7�D���t~2���EzK=(<��[0EWvM"�>���"m9��0!�Kq�n�g!�٘]����}�5��?�ze��mD��l��n����a�Gp� ���F�q�$�n�^����d���Y�!�CQ{��:����&"BRVZf�\}��CT�W9��n��z����D:w�)I��&�ƿ�Hߛ��ØK<)�,ư�G����R��E��5R�k��}dxh��O�O��>:Ua�+�B��H���}U[�7o��^~詴V�\j�� �ɴ����Ĵ��b��6����p����/������(���F������'`#�������8���ь���y��Ne��)(z���M���.)uB?� ��W8���?�J�h�ԕ�O~|A�#<Ltk3�M:w��e�K[��3�m��Ӿ�!�Ӫ�n��w����Lz�q�@<���s��9��R�^w���>�n�>dfۮ�ǂ�E��������$i��D�.d�'/!�O�P��/Z�tn�/�?j�C��fb��)��#�\�⑱`�X镽���W���9!VE���ss�>�bn�=Y@��ЌЍ���V?�S�*J8Ͻ�_'?�0��X�^k1��A���1����IT�2�s��{��5v�Xs��Rg�뵔G�$�7�=���v��؁��[5�)�����D.S������ӛT�{rjJ�iv�k�<��A ��/G #�~����e��((xb�':}�|ٞkc�����G�<��[s��4=I�<s��
�t�o��|�z�%����@,��Z�1X��\3I���g#8���� ����_U`o���=k�*�����6�0�w6D�k�`�{��E��J�Os*a���\�7��Q�2,?�QT-G����!4=�b���f~op����ƒ_?{;��7�k��:�?/�)���'�|���A��[_\��AK	�n}�XA=���%���(W=��Y�2!ی��G�@/�_)�	�Dj�QA	kO������x!@0���	��S���*V7`*2 IC�~73O	oA��S+&EjU&{v����A�<�tNIa���n����<	i�����^�ϥ�
6�����ԣ���ۭU4�
����#��5��0��d�=a�~��3�ƀ��b�����R�
`}��ʎ�hM�-�\ĞJ��Ŗ(�ޕeW���pN���a4s��-�7Ϲ�t�z�����Vv-*��?yx��Kg�oʒSxW��Ύ&��)W�H`_�]Z���JǏW��v�)�����KdrQ��f�.hyY��?"��y��E흗bp�� #�MV|)��5�)qز�{�q�� ^=bO�������~��E:�=�nG�?@���`���d������o$�,xP�!v���'�Z4�x�.�e�!l�A��P�� �*{������i�8 8��(� ��}���O[[;���G���4�GH�Ḫ��z��5�EE��[�qaR5=��/:1�f=JW�E���c����ԗ�����:|v�2�;�#�/��5���S�\:�#x���͐ӄ�(T�8a�+X���7�1�X^���T�vCp�����Z���0R>��S�����(ў�A��wr���y�j�^�R��]]T���;҇� ��?8x�D)P$T�O�3��&X��]C�[�y7�jR�Ҵ���p^���E+�lkuM��Wݙ��	J�&Zg�D�����_(��_��q���6	p�,A�4#�PM3s�|h����/���ʇ�k��r���9#�&]舱-���a�	���X�A5W�t�*�i���X4 o�=$<�K�Rx�_���"�ۅ?�a�ZR���'[m)k'X�'�(�Th� g=�e��Sm
jL�D`Xf-�I��2��ܟ�H��-���}z���WA�m�N�b�/���p�a#�`�QO�8+�~XP��<�`��ݛ��r�p� XPM�lp�×?k�\��%@~CB�u�'���"
�z�}`��i��!FjU��-��r���a  �C�y�$�eP��~}�9��3�� ���9Y�Z�.��+��5�2@���-�P�轒��蟣]�D,!1��(�P�;(��[Ѽ���x��f��~,W��)����J���gf�����>��)����i��r�N�h�OP���N�{�D�ϙs|�\�
/"�����L$�CG'�s�M�@���p���E-��I���]�Ab`�j����@���#Z`vJ�:ٍ�BL'��[.d�t��"8~�M�����E�o�����%�֏8���
��s:��S]���s߻L%�w��V?��O+V�g��C�%����V|K!&.>���PwN��D)����k!����ɑ;5p��a�: 3 nMޣM�2/��/f�S��L�3�R�bf�;��(����'E3�����Z�L5>�����C�I��/���Ƶ_u��N���H��_���������r 
��p��{���2��?u(Չ�=�)���`���t]`���b����^1�8�[ �i7~�Ź�vK�҅�	��T����y��5�Q����աb�\Qׄ>8�������Sdezz� G��S���&	W��;���E�c�I��d����|L�VUk�R<�m&'n�����\���7�P�4��s�����&w�V�����}: W7��}Z��z���&+�{MIרּnI����GnJ��c���6��,�Nx@�*�_9�T��6��Ty󍅗cQ��30���xXl�7�]̲Q�������]HH;���Y�™����`@0�?P����I,M��_YM'Cl.��FJ�_�𦚵��z3��� kMu���w���e\`�@���S��sLT8�}D�� �i��(�r4O��[(,þS�O�N+z~��(u�W���i��Q<��E&�ӨS�к2��[yȯt�!� �$�]���9�v��@je<�T�m_��]��%niBR��,h��<*�(0�\���j]X�_�Ӯ�BL���0,��R�n/&e���A\�)���$!�|�v�,dǕ��-\Lk�_�`2(����V��xJ�p���1[fݶ�;���da1%�v��`-��j#����tck(��Ղ�h�]�<:���ú."`�+���N�YhU �87;I�$�0:�)�TZ�{�i�S,�b�p�&�7�t���[�T9���"��D͙h������[Q�A��{H�Z��)��d�i�䙃�VDH1���s�ѵ�)��g�p�Z5#7W�]<�
�}aȔ��T��Ư_R��|��6G��^~�q�Ȑ/���g?uo�D��.q���m���sF�W�s�{���`�1�!�_F8[Y\���r�IÛƇ��/us*��⋇ܜ�|`�1�h:(s6Ǽ�8a��j�Ɩ4���XO	�k�+ ��nx�.�B��Z��*M�E�
fһ�u� }/�����C/Z���b7�v{�8X��{#�M�$�Y�KQr���γ+���O��3�%��0]�zu�s^�p��,��"u�X������DN�6v�A�뇎�q�w��K���6���R� ����} tc����?V����|ŗ9}�/�V��roeї2S�� TX1�X_ߠ�?������@��o�%(]�,𯍾��S�}C��?^���!�
E-a�?C�YI��FR�@K�ќ��P�M����n�s2j9Et
z��̯�.�RV�I�qզ�C���Ɩ�>�ߴ4G+��F���lD��4��f�L�;~��?�x�(@�����R��acMo���?Д�f'�G�����L&���w�:BY\������<s���"3�[.�@"�����n���|9��3|�ԃϖ8��J�.�4��jh�J�5g� �Z8W)��5��˜��l:�����Oj?)&���m�м}ɯ���{���O}�D�:����I,*B2��(����{��!r�Jq4ӄA�#���O��&�R��n;AT�a6��C�О����AK%����p�8���y�}�Eڰ�Џ5?~�)��!�h6F�����6��h��N�%��{��'��D5N.���Ծ��5|;˝����*�5͌i�Q��8PT�M�4_��>�`�JS����� ���]%4�4Q��6�*Q�q��gυ�+�j�1�~�o�g��@��	0E�<�Ќ�gɚ�r�N��C=}�[� �ka��u����39tG&?��ԏa�* ��_���J�B�n|ruì���̉�eEI��N��9�q�(�S��1bԈ�� �
�*eꬎ��fز����I�K��_��zH�{��
�3s�?���i�\o��༉d���v�8����4b�����s�1s�5k2	M�I�!]c<z�E|χ3�L���3����mM�*���:`j8:��S����a^�G�\����8j���HM���A�;������&�Ҭc��%���	I>�Y��>��g�I4��7Uu���+�u��P@��c�/��IYF�e�$@v�����6�e�>�c{����vA~�qW#_�UZ굧AC��,�L����RO!�9L-��o3��7���*���R&.���x�O�� �.��k��~"4�S��u�|$*"����o�pS�D�U��VFP��\��Q�ΰ�TR(��8��w'6w�+	�H��7�;��0�l>��y�-#�9ݟ���t�9�q��̊�ٖ�!��!&+ߵ �#;3}��l�J`�N�q�Y^�y���!c4s Cw~��A�^���ݛ#&p�g�"S����T30�/>u�oߊ�:�~c�f�)�+��t��7K)�����Һ���p��Q�q�~$�G��Q
�T���=-jƙB��5���ngyk6А$�V� zf����̒��?���D�@sB�>10@X�0���nΥ���`��Y-�����-h�+ج�MUG�w�M�W�)�b�������Gr�����j�al*�Yg�h�b*��QD�K��k\'��C�=�1���\�_�%�C ��[c�$7�6�>�NĬ��>嶌��aLAGޗ�*�&���xݳZ"4�c������b��]KR(�!�ʕ�F�tHg���aba�maǬB)�����M%���/�����}Z�AR��5�.���q}�s-U��BRHq@�ɀg���0��(�@ӽ��O�l����%RX+�D(��;���t��,�NBD�����O��ka������l+t���/0׏�]Oȴ�ʱ}��m�0����%:#����.1�(

�ld��z���D�^�b��� J�>���~��A�Qx�zy����ņrx�	�yؕ�μZ����X�O�9����u�7�<�k"�Z��J1��?}��nL�m慿Zy/��WTrv��޽:贞&Ҹ{WQ���1�fì�X�i m��8J�#�
ז{����˽�a?��\Cyԕ�3��/�f3ӆ��hY#N���k
'hNu�Н���C�k�J�z����@ms�@d �{v'ZC.��[\�zy�PF�i����W��Ç^G�	vnrKrY��������aJ�����"Ǟ��6$�TY��k�d��ik|U~���z�(�/݂�)s���R`�n�X�brKl�0w�%pn��XH=�(�a��b��Gz�:q97۔(��`���;I�3���Yl�����v�1T�U���^���ke��U�J`�%&����nZV��_��̞�|���D.V�d�c� S �r
T#h�Ġ�����u�z�G�h�hE	�n�'b8sCI�m��M7-���{���ˢa�(*���%�ĬI^m�_�i�3r�|N;X/�����g&�5�N�:�^�i곿�[���=gN�C��
jr3��d�[��B��2S@�B��h��Ǚh�~�4�x:�v�B'�C������a���`�i~��*R���d^ko�S%��P�B>Ε43+�V���E�x�@_�b����1JJC���6�E"q����!�����a�ZF��i�W�]E��!�Z*E⠢V���*Q">}?˵�G�F���Dk�+ta�o�t. �ң9�f1z��%^Q꿟Z�6�$�dD5e�=?"�Kb
i%#�4ڧ���1f�q���Ť�w]��D�e3���\�p��߸��Tl���P8��B��È.�P����`+�I���n�#����v�;��x'F���,Bq|�P�u���¤�6A\W|��!�IL��Y��-4��.�8-+�A�2��uu9ȕ�:�Y�Q�Xui������'�C{�k5J@ 
(4z����L�~;V.1\+$�qt��Y'6_�.���z�XPqN�������'0�]H1Y��s;m ?>��۸fC���L<�E���~���J(xw	��O
=�	�r�
,�ަ�V���1&z6��l�]���`�+º��c��,;�O�D��\�X��M�v^k��h�R�̻�y.��e�#ْ�����b�Qv<��_
�{ͳ0��$�h�4�����7(��;�c_��(�/��溋�{���z�g6�v��-ϸ��\�\M -��wd܅���I��Y��r|u"��p�������d_0��DH�;V��'�Y5(���YXu=�)�yʃ%����/�v@� cZ@��>.��%l{e�Q$lw��}����؅ŗ8�I��ŀ<��F�9�����~$>�B�;n�jr%��ͧb�e��hE�1y��s��R����P���vM$�U�N�w�Rၲ9�y2%���3��;�t��c*@�����4z�S���( �~knbϔ���p�s���­ӛ[�5�5@�0T�n��,�3b7��Gh%Ig!�����=��k���(f�bg� �Mm>��-� �U�&��<��8���/Ly�9I ,�~FR�˫���:6�(�6�R����p݈���VQ��@$��z��u��,<j'ف���}���r�D�$�~�x�6���ݍ�Q	n��F�WRVU�n2zU��Ha�Y���BF���&'?X�#�Ɏ�@^�+]��Y����Т��x�����i�~-��� ]Z��ؔ_:IO	���L�!�U��!aQ���Y���۩_�;x����y T���ԗ���O`� �	�ݗ"�̝�fW"�sV��TC��q+ߐL���fG/d\!He�i}���+Y5T�I�����uW��U*PG�j��s/��/ �R+�[�<tXW�W��Y��.:vߘ��D�E/'`�_+d[�"8H-�R�]j����|U"���k�Ź��N��,6�>�[�3�b���[��}Pem�C �+�^�� ��/�&R���Y���2�˺6=Dqt�*�+?S��j(�51��$)3
�0�?�>���/)w��s�#�N�	�LY�؞��l���]�<+ƨ��~<E���E�����$Y�5�#]5����,�tK�E�
�Oˉ=����Hn�m<�!�z.Fîw�m�UǮ�e��8O�����CK�
�g�� �'����]¥1�٨QI�a�����f`�r}��'Z"�[f G���N�FV��x�Ґl��Fϴ,�(!o�3*�Z��Q氅�"I��]CD��(L�o={d�4O �֜��^ۓ�E���Q:�B�Wg�oD��ϙλ+��sF�]��1wqL���5����Ĵ)�kT�;�,��S�ȱ���ۭ��UR�+;�s��t��VI.l�!�����
��v�C֩�W�8�L-Q� N�2ky}�<É7����%Sw���y����z�֕�"ƽ�ƚ�p�
C��E_�,@=��TnP�I�A +O����प��d�	��?�~`0���aÑ�v��G/N�Q��%��IйY�kIY`���a�ʳ��eJ����H�(�	ɰ�RWl�x�T�;5b��ܻ�
7 �y�3�>�琋̈�o͌�8�}p��ڕp�%c��#A��QRHW�eW�~O���*�Ŗh�<�6�$g�뚛�X.]R��.�V�s(��-�V��+=�T�MT����;�gLW�x�v�I2�8��G0q�����9���#���Ԡ{FB����P��ݠy/���
pT.����H�/�`a�IO�X���q��[>N�A�_��Y���P�P����]�}���ݮ~�����Ȼ�%����7�&�G�&KD}���O�΢E���%��Ǵ�Z�R�;�Vn�1Zײ��`K	<0��$$�XE�ȥ8�/��4cR&&��Q�4_iv���m�1E<\8�~��tz���:]&H=����A���h�'�@�-ف]��4pZ�\��￾`��TǍ����S����!~��#A��:�l��u#<������X�AWs��|��Ld�_7���C�r�١�{���؜�@6&���X���V?x��F��{=@,�mQ�������[�C��h�}�r�ֱ�[	��en���3;K�(ӋU��ڏ����%��@�S'�:��ߊ��i��w�+�f�wҦT�A�7��Eq�(�cYpao)M��5�[[PR0����`";R	y⋈�-D�ě�̝ڻ����j����	k��ml�������
VI�[�C�B~,O�5.��t��BlX�,�H������|��P!SαZ��LK�폹������ݹ}o�ŗ-F���o�)���T:�@]�-��Ev#� ����#V���3~r��:���@9@4��O̚��1�(Ŧ4��(n��VQ�/kJ`�̶)Lg��oxi4�A�̅5-�\3�_�e�Wj9����K(�|��88}[ ��ǔ�9�,�x,߯�&9��i�I1CS���Z�@L�xL��;�TZ�w"�	��sTME��w���|xXLHh�0_�J��ze�����N�j`Ձ���*qs��5��$E?�����:��8{��(�]�`�9�x)���:jX�1J�u���z}C��[���)�k�X[��Sj���%&^��|��}����Е�v�c<�%A�}����4{�h��7�X�/�5���e5B�<�6-�V3If}�&��B�5�/��
��@+�>9q�ؽ�Z(����2��Xx�+=A�O���I��{�Y�N L���R�Oxt��Ça�͐t�ž���i
�&>�fi �5��D�=�U�Sj�-�@�x]��Ϝ���.xEޅ׍�.$��1p_��}�򷏏-�81a�%������:��}?Җ�;���	�j���#����N�˧��z~(���5�w�#�P"|�J�T.�Læ�Y��c�e���󃈟��IRf�ּS:��]�L��)y���菉��uY0�������� >-�g�J���%�EfYr^^Q<e����&R����Rc��N�^A)�6s��Z�������r%���B��t�����*5y-���f~�5�%|F��ጓ{@P����ʯ!��Ō��P�����T�̂��+�/���H|b�G�|�	c�H?-x�5��dWk-���)��K�k&�K���`'���?�n�(='xY�?��(��A{�����q[s'0�X�3�ǩԧ�$�pz���?�5J�|F�7(�Gڧ�R*Π{]�!My+݄��d*�İ�[=��uD�nh^����$@%�7,�y�8<�tJ�!6�L����EϊQ�4��֍u��&�E0tTq�qы�+2�贪xA"�A0���)�s�Y��f����Sd���
������j�n�/��nB��ç(��������z�_߶,���&-	�KV&yܩ.��r��9���ݡ�2���S�X�������ȵg��Kē��D��sa{B??��a���(S����y�n6�lL&rܛ+�	��T*��e����'}�U+B�����˅��23��nw��9!r:irB�~>ϟ�Ҽ��A��!w�⍪43pժ���3���r:=_��ak]t�77�$\�f����Ey�����%�� ��d�{i�5��t/����q!�h���h"x{}��uۿg�����G�.u�v��i�vl$T��!vz�,�<^�6 beT���l���^0V]ZE����8�z�+�C��=�'����(@1Y���Yr����K~�Fs�w>׿*��z��e��]b6ힳ�����m�Q�(�f`VpV4��ڗ,V��N���	nj�Ҭ��r�]���J�~�q�η�x�8 z��G��٩2���8�[��c	��Z�J�^~����q���њ�#E��GtIݫ>�o��
7eλ��0����ԅ<$����#n�w?�a�<�4�8�W�Y�~��ڇc�iu�T"DC?7z�Q���Xl���\���+���L��è��e}T��Q��������Dǵrh���j��eG_�����n�;6�����B[i����d�7zX�c��162��sLv��G��.�XZԩ�E� ��c't���D�e�e��$������i�6�|m}��G���@����)f�o�OCÌ=���]������r�%����N�M��F��}�m�-�K��N�T��MZ�D\	�0ࠝ�~�'��xw$FWn�� MH�)P5�i�����,r���a��D�,(E3z����7Q��P�}0�Ae�p2(R��y�ۖ�(�)�)�Q�� r��~�P)B����"�V�Ė	+՗�5^F�NvU2�l&;��` 8���h=-�!����rᆞh���:�dfF-뱡�m&���+Sl�|p��9�p�������ڌ���Z�����ZhϋPX)���|�m"��E�aʜX�O�Ȇ
|/�����M���x]�Z	=���G�6����`���E�/�[�f�X&�o��{�i�oGD����)�wL�L��h���9oQ�������������-U����+1}���vO <�]uME��� ����p4���Oc�|,�cr�H9W��"�������Up���B��jL:��L@�w��}���AB<����ؐ,�l�=ҋ��?[�t�6�Yn�9	�f�ʛI��<�nL�L��i��6���l���&,��>���V��s�߉y:	�zd�!1ȴ�@��2��Rv�!�Q�K�JZ��j���u�eEY8;:{�L�`��n���g�@b(P���	�)�6f��%?U����t�ɔn��Q�}f��8��}�����õ�`]�	|A�ʚ�}���~�_:0�B�;t�I��f���Y'�c��
�n�Dr宨<{�
@/�cQ�e��Z雠������VG�-�,Լ8K����3=N�?w��}4aݮi|p>�l)���1Ac�n�^*r��g�w�2ErN��r��L��F�8%`0~O�8n�}�y�|��Ri�!��F
����\?QF�t�%�v�Pb!$�Ɲ)�ڳ�Kt�SM(U���.8��iq���$͑���� �qt�W��CLh�%�ն��K��w���1Z��dN2s3�Q��Gr�8�/�b.x��w���k6v���%�MD��YZ����Ӵ��w�P����w�r ��|I��c@=�R煎6q�h�׌�o��3u���G�ɡ������V�$[��f��>˫e�Џ�sq|��w>��&�K��J'9�)'��xb�P������N�\$����w��A�H�Eq*}՛�湧;����3�Y?�͠��+U"�|e �pz������YV�� ����J п��'l}�|���*\R*�9�x�S����~9m�_�����Tj���@o��wp#��ngs���K�s@����3����*n�)�\��*�Ev�=��d��h��!�����{=M6�-'�Κ^Y5��5�O��_�sk0��ID�w_�v���hX˴�1h�"0��֯g"������(�_���8F��% S}�c���Nf��B��r�c��o��+��W�9�[=��%�m���Ȕ-���nDet��~a��	��O��/H�P��W��C<�V�$�K|�1�:���h�k> Z�5/�R�L��H	�,�]�%�{|�����P������߱�{�o\�^6���3�ugx3���H�h���_�S
$�J���H��%��"%[Y���hݤ�.iQ9�
�TX6t�c��.i[���U}l�Ĕ�<u������
����Kw��0#�-�`f�X���I5��q��Z�YL�Q�zь�{�����q���a���#��c|�+#?V3�2�l<�SE~j���xۿ0�0c�W��T-.K>O��I~T��_q��o���([%�Ə��F˕26@�6�޲��thΥ5����DhDG.O�\��kl�k��X��h�oR4w2�~����� p�<=O�6d�� U]��x*ej�����A�{H���j��^I
�O�!F��Ldpu��S���������>���h��񳡿�{�����oD��o5j`���E"�6rIN�'������Hq�y��DF
H�B��������	p��!�KДK9O��SFs�4PX��x9��ѯww�XJ�D|_Q#e�Q#^?ظ�.�FDAXvD`�*�|�=U1ۥ���e�"W����(6	�?cIS�4 �Aeȣ*}@I����OJ3�i-M��!Rϡ3K\�	��'Д�tY�0�M� �d�4��p��A����!?�N4����k�L°]	b7S�Ļ	�w���QʐQ�&mM�=���L�@�<�t���9`�M��Ŗ�dE{8�����JֈI��{��[��2#���'�)�Ѕ�	����a�OU"!����gC�rZ�nw$��
"����z���j�)���M��	^ԃNw��ss�s����ޯ�-=iq�9&�������@�6k�3jX�"�h�dϡˁ
1Ɩ��m�����eQ� ��/6������%�:���-<o�b�i`.G�,�����߈�E�͕�aR-8� �Jj�э���݅O^�YcKˋ��Ǳwm
6�J�fC��� 0�m,��J����"{?~C�9]�`)�y��;
��ޫ��R�1�-\�>����{Z4e$�tVQ~�;R�*�TҰ�'��ї]z�}l�8�)�͇�w�UhL����Tl�j_�G9���~u|����{h�E��|��'���(پ�L�G��]�T��2G�2�íy ޿� ��\�wE���a��_'R`�u>@�S]N���ԘI�^P)� p�{X���I%�t���3柗X$qq�{�Ӯ��f���/o�&�e[j�\�	��(�m�����&!�2Eq�����@˫#����$�zh���ܹZ_{��T�BC�t�-E���|b�t��� Š-�/���G(�.�8�v�{��������e�οDW@��|m�b�	���j��툋|>��K�M���p��^	Y� 1���cu8���d�ŋ	,�&�OW~��(���O+]}3�ϰ�ԍ,^�:�/���
]�������pC���vo�EĢf8z���W�|��(ж~pi��螌M \��	/�{B��q �>���X�]�'*��2ؽ�j�i�*[`��O��QR�܍*\a����<��J�3���N���]d14'gjÈ�kДҔgVu�P3ds�����ɤ����h����k�2P�Gff/��'��RZQ}�8��<�ȧ����9�cIo���̛�-o�仠�n<N�]�G�=G������l�84&؇i%���S�&��.�XW�VU쇾M}�&�}
�.ds��O��$<���ɯ��ۭ2,���6ʯʤ���C��j>�!��ƭ__��?�8,�s�5@�"�Ԁ��<\�^�y������m!&6ś��ʲ���V��fd�����*�(YO`۵�72L���������\�:�2X�=([��U�m��:������������i�ad�5�+�,��N�J�(��8M�g�lf���e�����p��R��g�pV�ŔRqS�o�B��� �DU��6�	���٤��QS唷��$!v�!S�X�H@�1��c��3�Jj��Y�"���lT�Z����L�����)i�K����M���:������c�@C����(Y�d�q����� #��4���1�ǽv��Zϒ�a���⺩�<��.��O�}5[��|ᧆt��EsDҀ^��rʌD���}^��\�7ZDb�!EH0^�C}X.1}��`	U��l�&�a���&��Z�S�,$^\!E�|x)W���6!/A0�`o����F��"��w�V#�DѺ�e� ���h��i�$ �&r�D=��e���mO����[o�3��g��m����q�v�S�5�;����F՚4��1ܬ�Zk��H#�_�nOH��B��G�5W�_��4���9|�D,23����;I���9p^�R����lo���ݑ������2�F� �j����8\��
�e���C�Q���q�����.����F���QXԦp�Ѽ�5�"+k��j�j1D�c��������ßa�#��\��l'*?�۸�%WN)�b�C{>]3۹�X�DV;[��3[֢��sc�9�/�Ze
 ��2T��)��l�Xk�M��/?ԑ�����X=�7�FT���u��;9#T{�2%�:#�al�����	;xF=f�;_Dr[�Z���ݯԠ�F�������K.��?m>���k���j�c�Jʕ@-)q��F"��a�Ԓ$D#bz 
���Yb�RTJԼ�yI�BK�U�������k�7��Nf�)ēi7G�8��b|��7�f�t��E�h\�����B��7CX�P����C_l�H�2��L��ϓ@�P��-d��k�#�3���'V��ıj6����������4#~5�r��\��R.=� ��
��"7y�}��C�Y�e2�Y��NG��m����as�'��2A@��)�:��n��}�D��"<"�9V�ek���Z������i���D#;�:Hi�t�'qY^]�!w�h�/m��<�ȼ�.�V��2���*�bq�
��	t-��Wu�D��5��zP��Ok2~�)S�^��%%�J4�=8Rb���.A�.e��=�8��Q�AЈ��2t�N�9���E��\A@J���-Bx���v[Q�[B�lF's�ݬ��PҌ��&�
��!�Dɻ�y���
���w��R�v$���bY˞���j��|��?���[ �d6��o9�ҊJo����B�4�T/��w�FI����Q�ו��}gGȗ�E/��Hp�*{h'�9t�#*1�ȅ�ahɭ5M&�	�2[�p?'�.I��]��8Z'�Sʖ�ө2|=�2�cE-~�N4ј�E�m��<z�琥3Y` h�C������)��T� @"���&�$���}���㞌��c�6#��=tWo	���n�i�nل����/�8P�l>j�}�>�$�O���"D�R��F�VM�q���y�<,FBYr��5|ן�U�s	�i�J)_CD�<*���xսsib��-����/�_����Z��3����Dg��u��D#��A�JϾ� ���!�c�4�YU��y3���P -��1��`2������=-i��t�~��8Ռ��x��1�J}�ˬv1�Y�
H��|�$*G��R�)^�a�Q�-�l��U�kk_2m��c~�3y<���G���s��A�+P���f���<�#2�5��8mP�ë��ξj@T�z�D�?/�-:�b����U �p�G��,�vL�������o�����6�����&9�X>Q�_H#l�wNQ���.�C�i7�l�e�a���__Z�w���ZԆ���<�s����<Z�GW�c%�/��e&�}� �k��Ƭu�檞�!H�i�[�-+»+.r�j�3� Np蓂��r�=\�@@���."���Y��\!Ӗ�ZH���B=�RD��k�����E7���=p>�����n�ҍrN'��4:�{4�Bt�$>��{�͢cP�-��7�z���%�X�m�'�"�<+p���!�����s/ Q22fR�s%�ۊ�� �ƄdQ�

m�����aJ��Q�ջ�錔���i�S� =�*��+���z)��i�����q�o��ݟw����៩��I�x��5�Hf����?ÀND]��r!Eh:�cf�9����v�J�+o�e	d2�;��I�j?��q��I|K2��/�� ��&^���oQ.+E�F�s�?�J:�����F;ł�ٓ|^�)76+�i{|�E��0�ڤ��`�xN[�tG;������Rx��b��ٗ�*+�*E�k���ǽ�n�IM�;�{0�#��\��_�����\6>�1Ai����u�Y��)w�`|��r�<����q�&�:а>_��)�[+�I@�!��EÆ�{�8=�A�dT�mO0:�z��^���\1�D|ny�KVT��e�nS���0)�S3"�j���*(�p���@c�Pʿ���\����F���_�@�a1���j����y���CԤ�4+.a�v(n}�~�K����2C��9��X�}e��6v�t�(�D�� �vI��'h8f0�9�<��V0�,���Rey�a���"�'Bj����rC�\�л�������W��/�Kwy�j��Թ��c&�&Of���n#D��I�)�k��B_�.zT4Q\�n�����[-�qi`zǸ����~�6�ş$+]Q��r�n7�o�D��s�na������}����Z��i!���z�׀�`��6j���i���9��,��z�P���w���ޖￎ��>�'fxx�h��I�8�.�����
�a4>9�|�]OkM��� �iS�q�*��d� �;����J�/_մ|Vp���7X-�#q_�J�ө�y�L4��yV{qB��)!&u&����`��T?��������D�Ŗ���3��r�7��F��[}m��At�_l�Fh�fb<����P?��}��c��D+�E:Z��p:A�{�+�L���
�� ��)���%`��1��ahp)LG+��x���^*�:D�6R�~�:�|���"�t��n�k�y9��}����͏�1�:v�F������1��7�Y\���5�#�����Jv���{�EX�w0��L2a��(#�� ��?U�7���u�V[-qA!柏�dh��G�@�3ɩǘ�;��0I)x����&�G�(	��)4�X�AvIk�jd�/<�0�sS���KGQ�y_�!�x�%�/�,��� �o�|p�|�c�Ӳ�V�ξ��i��\`;��oo�N������+Ý�;��-/AϠ�`�ٹ1�<�zg�{��oh���(��>d�����M�.�bV?��v�ư^�_��w3��*����(�.f=�����,6:'�J(v�6%��Y��j�����8И����j9�Kzd��U`&��1� Ha�l�~��
��gW�_	�����?�T�X�����(΂cZ�p~�o[
?��qIB��eaW�j�ݳ�l�&��P֤F4�_K�hY�h�)�"���C��-4�O�`���©��π�=���������cv;��]LV���n���ᝐI�#���5��xb䤍	9,�WE����۴"/ P<}�+;Y"���i�F<&)�Z%���ʧB�bǮ����Of|txu��Ǹ��%4�����/��F"L���ǜ$����>�)3�Ż�m�Z��ȅ\XpY���ᰢ�6}Nu	#�����ڬ.������vn֡nZZa����rui�?ۄ�Ysd�n��I �7ȃ��W�=u�JK��a��M4�ff<�3̎�EC����v�\\5�������(ᔶx��X�ٕ�@������Ka:�X�˾�%�I���i�5ɓ}�)��댛����`������"_�����P<IĲn5Z�N=%��8�It�\�ٌ���c���9��1��.6���(������
z��6�'��}��yZ_�����ED?UJ���Dd�G~�y�+�<Cp��V��
�ܻ��M2�e�O�u!}ӧ�/��f�^Lj���<��L��C0@B�v6��=� �0%O���ƃ����D���0.?e�psOW�r��Z�B��=���nF4�dÙ�t�F+z�� 'L�݄�Q'w�Y3�wݏ� ���,���T}�S���p�P?�v"��q�L� [O���O{7���7E)8����#�A����y����z�Z&�4�H�� vir���S�`k��f��nZ�zʼ,\�7TFĴ�Նp�Zw�ċ_�v�v���s_��[�5��L8=]������s�����a1�]\��s���?R��ޭ����]�b�E��rC��׋#�����R[��Ìk��-̚�KD��tx��i��><�s{�y��h���P7�hݚ%����^C6sM��v�����#�gS&߁c�?l��� U����Q扣�L3��`��T!4mqC��]���|�:��YnP̿�c�y?���y�p��0Ѣ��d�Ӆs-�dnx)n(���N��
���mf���!�y87�@E�EK�0��N�.ǘ%�',B�*���(ņ���[����u|+��'/!/�wʹ$�Ф��r�ki�
�X3�}��6��
�Ĭ��#Us�׋�4�����##]�|��M��ǐ�y�5Q��.$��+��@�O�J&!��R2Fx�͗�)� ����o�&�8��s�Ք����"�=�q�V>t�E#nC{6�*�K� p+`�n�������rݯ`w�^�k��֨9n���#���+DՏJ	����)O�|NX/���0����p�YX��)o���[�B���cg���{Q5��T峖��l��Yе�0?Р� ��D��NF�ew��jҲӍ�K��a	>�$L�D}�s�(��#����^����_M�H�!k�� ~�� �(�}��<#��k-c?C��`�I��,a�a�ch]�b8I�/+��AP�P�P���sh�r�H?~�	�)Y�����2��h��y������`�[��/V���j�E�|�w���S�j��c���}��e튜?�ƾ`�w8�N`3�Z��[/l�j�w��}�gPS�Z*a�]�{ H!u�d,�Dޞ.�V���%0�Cw���i [ E������Z����_��R��I�.�W�6?G5�V�fԝZy��)0�t~��ґ0�#y�pkNQ�Yl+%[А/�Ul�x4����s�"�l����J�A;����
A�}aA�עQ��+�&Ű�k2����XC�%�{� u�)�@��!<���%$��5iߑ�z7��&��]_V�¤y�������%U?��a�fs���Nn������V��r��,��w6�w����0
����6���J���._ԪK�I���*��-k!P�S���_�Bg;�Ř�?m�-�\H7-(�c�y�X����%s4�o�ȞU������uG�h߫á"��j���&�Q�-)�sX#�;�д������J��	F�"̑�?�}�C̾�k��;o4�k�ɮ��ڡ�w�L/;���#��$���ڌRD+����o�I�I4�
	��P%&�{���Z~f��T��Q8���v�NBT�萶�6�|x��?ӛ�-}�ћ��X&/7�~n���02E<���slG���j|�Wy=EY�-��m��� ���_�nGΉ=��3gG��+�_)�u�A*��D�e��!'E:�I��b�QJ1�H�|7Ϳw�v��L]�Pa�:�k�'ik�������
)�tȠ�O�gŞ$��Ċe�������[C�F�u�v���rά���Oa�܇�X��˫B��pʘ���6P�n�x8��~\z�(�$�v��f�yQ׏��3�L(���"�&|(7�k.�N���E���������e�Hӷ<RZz�4i<n�Xc�6��F��/% ��z��q�߈C�-Z�틨�~d�;nZo��ݶ�u�]��s��Qp���qyMj��b��ɸ���hi�O��ה`'�{�F�Ij}�����Uk��;{���5S�k��՗_�*����MzA=����6G��0�׻\f��@��]ݲ������ߛ�"��_�G~�>��� ��^X�����H�*d�':"�v2�à������)�T<�a@j������d�q���K=���I���g�oD�1��S.e�;��-3��a���L~�W�6��GC�I2�I������YN�?�XH,CƎWE��l0=�W�� �c����Am1F��hh�3� <7tT/�.���M�g��qj�F( �j��U�c�B������_q�TJ9��:4��	���+�R�pW�^nz%W���Z��u.���g*bM�T��_��gXi���6���S`������&_���%�Ie��ڱ���j�$�;��+��)WT �q����x��Z�{��d�3Dנ�炦@���|��t�b�f��:g!�?FN�Ӗ��%��N���Y�
��׌������%��&�1�Gl�ӿ-uM͈�}���K~g��en���)Q�&�}م�#˂�r�&�/o�?�]�H��c�&&�XMY	�p���@�o�^�M0Z�nJ�I��((jy�FC���ͲT��~���,�i�W`γ��y��d�� ���xs�t�h��]�j��{���h�j�K5z�H`���Wy$pW�NC L�i�(BA�跡�w]����9@Sf3��\D<����5��ʕ0S�/2h@_���9?p_��W�:4�NK�h�AU9]�����C�d�v�:���PH�x�w8�>6�|�G���'Wӝ3�pV��� ӑ/Z�b��#�:��o�܈��qz:<�x�*��&�+-���Au��@c;���QAT���tΟ�9V��r&����e����x���W��F�%Ļ�k�Y�Qd[J�Ͳ�a��^�rt�`k
ᬭXx'5����һ4ǖ?����������5_2�#��Ju��:�����S�:��u���(�pO� Y�H`�G�E��#��b.����;�H��V��Je�G�5������cF��FG���j%��.|�d�����C�W�W>�/��9.E�*�f������ �]��C����j�Z=��q���xm���Ai1����&K�z�*�p �"=<CڬJ�j�L�M�u�!$±6�3��^S
V[,��Yu��;�7Mz�����YH?b }cF�=���eo��l�E�}ߓZnDT�!͕]c瀛��[���L0%�t}!Xtk��G�@o��JK��O���4KY�dpE�X��d�s��Ieg����5s��Fp���܆ʝ�֛���">g|��r�MHɍ�ĕMi���A��ռ�3"��Vм�2I:�;��jp㽶ֶ�w}��Ŷ	�'y��W�1W��R7L��.i�LE9���[��[��_v4ru�;��#�2s�������#���T3=��d|�z�}�O8��VxAj9�f�Js��?�BL�KDq?FH�� ��WHT���r�� $�0�V���Q���-MH0��'���k`���Z�d�	��BlٺK�� ��?͚ـ�ACܸgV���v���״<`]b
�k�~&{H����~w�i��%y��c�g� �b\��T����+ �zo(�$�;?V����_�����}�6?V�_�%l爛�,�S�e���7K�gq|:�62��$�E^l/�\�Q�N7�ևk�0$?�C�;����>{��z�~t=�좡@]����.,S})<�hm�P�CFMLǛ}#t|�u�b}C�_y�jA�Yb����t{��%��$�"�D���mɎ6����G��\Q����팒,ܖt����h���*"��0
wMG��! 2�j�F���"L�O�tk�>U�cqoqy�K[�d{�
��Gu��� ��A��bN��{;{���P�����s̒0TS?
������ES��y�&���5& [��&?pWsa.y`�f*ud��H���3=ǉ�9/�P�������,1,X��#�ւ��K+A��ӂ�ο�-ȋ��]����S�{9�(0y����Xwoz⧔����7a�z��.������L R�ル��f �m�E�rUl�H���T�m�=ks��:)Y��w����|�4�����Xj��W�7ko]�Ԙ>�
$}���q;����vC+�Q@���/; zΟUR���L�"����t5h�N��Ƚ��r$3.7��@@wߚ�\OX��HLQ�%�:QS��t=�9eR��9_�#�G ���w�^Yب8g�r2s����gZ�F+MH�F�����Q����R���3NI��n���M�e��t�l���b�{���������X�y<�t��w�f�,!�a�#ݥ�Š䜋����!>o����d��]�P�X^
�(_?#B���|_�P��{m��HfN����NW�#�}��ԁ��(�xư�!��Y�H����ӖԤ��ޮw\q,iID�ܔ=-m�^�-M�(��F?�MYܠ��:ƯxVg�B�/J!�~b,���rj�X�����~�HHIh1R�|���
� 4���ϊ��c6:��(�^pg���)J���0�e��spĲH�q7
�X_	q
���ȭ7`�_��|%� :Z�=������|�F��R!pPR��x��`��y�;�;Jg�j��0�E������T�Y<(�p��W��(�g�^�$��pC��qk�El���b�l��}�*Z�m	/�wx�1��)B�� *���3R,�m����l������KcE9���a�8�8KY/���Ro�m���+x{2�h)�CM�����/�:��rw��wc��ͽ%�z�)P�M�
ݗ�S�~��˴H>��݈o��Ub����e<��r�-�ǯF~|̥{��&5��Gm%`J�Sv��=����X��bX��#�!��7��V["߆�̪.=.��7��%9:���Nv��B'���M�͉Zȶ/���q�J���Fi����S H:�S�ؒ-���9��xl-��3~���#T�C���U���=��$��3dB5��D�S�i��+�)���I�����l�(:NZ���7�u$��c{҄���2�c'J��e]���m]�ȗ ���R�;�ς��v��kc�VW�������<����W�� |2DUJq74'%X�6�Cn	GF��Ֆ���`/vK3��: �%|�K�It�Z@};�K��~�\�
�OR}���!�AM$m��B7���:��ֿ���7g �Ҧ<Fm��������f��g�#�b��ޛ?�h�И+�ߏ��V��\�Ѓ�12�m^l4V��}�}���/��|��
�I���j9�zu��3~m�z6�T8*Xs�_8r� ���O՜j����Z�gH��u5��?2ZN�rצ���*]���>��иs����O{J��}ZC�1���2���Մ�e-ᇔO�Ar5���Is7#� ��� ��Q%5�H�g�hI+�T�K(��ȹ�V��.n���\T����p�%�����4�4���>fmM3�p�d������A��A�r����E,ɹLJ�G?h�NK>�_����3�%f1�=h9�aK��#4�f�>+�n�����0}�����ԑV;�%���`Ɨҷ��b4�گ���N%>{R����ThQ���6V��GՀz��g ]�"/L_B����F>#�6R&���r��d��R)�߉ĒS�� ,����"�:8�ݨ}kH?�_oh���Eơ#�$	ګ�,,�b��I V(Lػ�a˕��ᜂ��|55k#��9��n5@�� �Yv�
m�z;��H1��-�+�Z��E_�ڤ�$u�M#uVq]n���qS���[
�&�8�A^\��W��daC���fʛ)k'm�e���A�����H���AҼ��HI�E
�Y؛��fa�Q[v3�}5)�"2�|�R��-?���^K�-H�S�ב�P	���c�	.�UN��b�v8����b�&��@lS?�?��*�����Ե�Ctb3��'�ʬ�+���)Av#=�ᾼ�Ҁ
U�P�Z�ȍe	�c"��t�S�T�4�O�5�MB��>u�~���p����S����W��l\��_8¶��!o���`o����|���ɲ��ͪ2��9�;N��̃�}��Iu>-��i�%'�g׹�d�`� ��J����w����|㮌BlIX``��V����ζ�(�,���Aӧ7�]������]X��e�m�sK�71B ���|�Up�,D�Q�R:�F�5�5�gy+�s�>e;ĳD3WVa�2�84U��	f��LZ�-�'i'��	*�u�>���l��S~Q9��]�/�Q�@�is���
+k�w7���#"�j�*�7h2�I燋�=��R��+�<��x�A����p����,��E0�������>L�J>�LEɱj�m�!�bX�$���������:�cY����fnF�J��y��ǝ�X
/�j6?�n��Ķ)NS�vs�}5:�k
��@�Z�;�F�
V�	��?Ϯ�c�k���Ht�|Ʃ���TRG�](��d��EL�w���d0�V���=����*)�O_�H�oc)V�R7��ۤ�r�>/��`�a6�iMq{��R6��ѻ2؅!?�=M��u�$��:N����B+�<�.��AV�T��^�BISk<s�"�����kԷGY����U�t�Q�{Ļ1��:h�pb�	����N�´�wl`�}M#~=
���PΦ���8J�G�b�4��b弄B����Z��o�vh�R��*�.X3�w��X�؎�%ͣU�qk�K]�Z�svN�]e��#�R����"]#�ӳ(��ɦ���BW�S��t�%���h�����ǚ N�C*�v�n$�����=�GL���7�"�Qm��eA,���S@�w^���n��&��"����[��jh�޵�z�l��9w6"\��"�t�����2�uPU��.coL5��4����{��S��O<��7�N=n�i2�(����=+H�w(� _G��`�sM�@ q�`�Y7�mDΪ�a���!���ɡ8z���_�y-{RiH7�y���  �'���X`uA&QgA#�\�Dog^�1��۸3s�걍��#�����/��r�u���`��~m�`+�ڳq:�H��_�<5	�YA+��Ol��z�1�#+�X���-��[3����<
���96��;���:�)�_�D;�iR��A�J�p�~�\��t�;gQ����S��M�G}��BPM�FfS�{ſ�"K���3쓱(:޶A:wv]1��[#�dcM���SmBڙ���T�F��Զ<�}v�_X��|	a�3�e�&�,b�>��f|9v��G;�Q+�4�Rn��V}����K�%�E�zō���e�H�GV��~Y� �L7s��P�_2{��@�T~���lo��W�+�a%��|S�r��H-�u��ի������3���ti��Qڲ.vN)�]�7A�K5�L��)��XVb�1�-ð/�	Y��u_j��3����B���������M
�~��ۢ)TA�b�c����|�A����*���#��1̞���Rܱ���[r��$�t𩄩c�'bzL9Nа�����]>7���rS:���~��#zJr�~#��0���釭XwM�~�L��x�m�MĈ�$/�	7���!}8�A$0�,eOP@��)�vi�?�o1�Az����P�9����F�������Sk<=���~<$�N#�k`�r��A`V��й����"��B~6�C�R>���jf�3+;���.2>�O�bY*�c*%��e��,����u7gȯ���~�X��n9��B��{�A'�2sO
����*�
�*R55�-?`���wy�g��Ŗ���wC��KZ%��g��q���l{^�`�����ͱ��~s��]r�,�S���k��Wg�w���$�)+t�e̘�Yy�~�W��wm�cK�"�j�LVJ�AD`|&��I�r�HCv�cԾx�ͷTʜh��",��l����]�\�9os�jm���!8�uJ�/"��U��1_�Sc�/+�Mh�]k��ޑ�p�7E�U��}����;�s�z���t!�*���+��Ax|m���M#�,�B�V����w7�5ղiD~�[t'�凹�H
3�6X��,OH/���
�����"7�mВ��ҭ1J��;�sϩ�?�nj�ɅfeƆ�����ߦV��Z+��[ǵ�䲦��z��r!8[G�.f�+��:R�2��Z��L�_�^ĳ��,9 <j��n�tj���hQ��@�#,�S��V�����@���m_��i�v@�xh�����u��d_>��E|��s��e�-������7�H�̓��-�#�p�V-Dw�^6�\k�G9��99Uo���:ƴ��n��m��������/�l���c�o5+�4_�?��[���J��/����\
R'����c'6��ʟ e�ߦ}"�u&�^�`��tL%�--�Hǘ������)z�L'��(5�����uD�b��֩R >���lg��;�Α����ȵ�V�Չ���N��9)�t��m�i/��s�J�@	�\�}h�T�{mʰ��*?Dذ���viє�E�e�� V��G�t��"�PⰐ��ɪ��pى�N�W 	U��Ɋ+uT��۲���a0���������̆�����?������r�վD(K�IY�H�ύP�6y�~�+�qO�@�V�kK��c"g����$�o�<�Ro��J�nng��ٚ�.��2��t�6m�L��ʅ��=Jc�Ţ2��Y��b=�;�Wl`�Ko=��BH�"t�VG�5���Ȼ\D���Սs�"�2Ck"sc�1Ut�&�el�3]���˸�2q1K�~V��,7������W��O��b]��Y"	f���r�]�l��!�s=р���^*�[*k�%�FAy\9��Z^u�+�:e"����0����\�w5;N3G{%!T5~��.�����H=�M��U�,���0[�?���h�%S���O)���[�������_G&������bP�eTh;�a"�(#B0^�F��O���	���\lkK,LV�!u�z��v��4\~e>�:�����H�A��-��{r�aw�������"�28�K#Ri�g��?b�/�� )8�J���������lN�{	5��^%����� o�4Z��,4�'�&sʉxNC�pT-p����̒UB$�1ֶ�����y>]��_���!���c�N�h��Jh�[�p_����\�򮆃xF>�Ȉ �8��l���z�"�n�%��b)��̩(�D�C�HYT��Y	�� :�dr�+2bu��5X?�A�-&��|���|�+�����.xe��[/GpN��[I*~u�MUڲ�V�؟��x�<�9�JB�\�_��Gb�B��dH��H0��]�����F�mUj��b�X����d9�����:�8ǻ�������F�ٗ�]�"�Lok���p��[�����=�6@�9A!��g;m8�m��fr��ຳ4�;��*w�I'�	D���V:��2ձ��
i���� ���r$�7ډ�,�{¯�ʦ�.����]�q�4q���KE������L#.27ZZ>���bH�'���/�y���E�x�9~p�X�d�f��\�c������CG��6_Ȝ��Kgm,g�$�15J��S��Ӻ4IAeV����f���^��-b)I{K���V��xA����ީ�4��8nC3ѯ��o���akW^�Q���9#����m|�c�閳~���9:��1�|
Tv6��^�y�T�H���\��v�q���Y�=��J�'i��ol�D/~�2h��P��`��YvM���3�EP���Ů1���)u`)�(W�w�u�
L�}i.�P٩T��I7^]�jz�η�z}PoF�	 5��N�\��
쒾���C<T��~���
9*ϕe�b��B}���'F���;��mA�̘N����n�5�E��2U��e9m�T"N�Q��b >�;�?����M9/�lH��y�sK*Ud_��27��}�E�M�&�@X�&��^��`����9��9A<	R�ײ$�z�q���wgXR�N�+<-N��SuN끴�	l�m�
o�?υ�(���@�$���N��$�7�Ӧ?s�h�xd�l:M���L��~�90�t�R)�bd�S\
%��4*���GEPǈ�7|'~t�D�����.�u\(LF��W �x���W��ũTq:��DZS�rz>UC����[cXDm~Uf�Q�e��f裩���;��� �"]9�L�U���i��iæ��o5<����ngϦؤ1��b)�0f]<���q����"�[Ϻ)V��җ������4�&��,�6]Ј�V�t��:vO�y�-��$&�q���7Ms(5�J�n�|�I&&��`f�����v!	
�<Q�
�E[	+�?��ci%;
W����.nr�v��v��kD��1z�N�Y~���xñ�)�U�[<���ED�G�h��Ac������S���q�E9V��Ł�0J������*��1i�J�â�M�T?��/��Q~@�2�_��p{	��?�O�4�ꔇ�FN���J�ᾟG��05�L@��wÎ���$`w*m�I,�F^��U�@���G��d�Z�,J�#�D#U��Y�������V��IJ�U2��M�O�#������(w�o>���v�¾<��G����x�k��8�v�;Dp�(���*=v0m�R�JH��GD��O_�l\hY�e�d�| ���
�v|���{$[F�:��uCQp^����۩�-��D;QZ*�q��K���2e�����!������;�#�~�Cs*>��g��m�Q�T^���3M �&Ž�]�F�|��ڶl�l?���R,�% ��Ah����'��I�Ls�6�M.�ݓck���cb I�a�[��B4���g�P;����o�H|�@וe�Ȇ��.<j 8|��C)��b�,�>5�e���a��{���m2 �;�| G�tu���u. H���x&xS� 	��n�3&%��G�_�xY����X����A��G��hJJ����g�����r�ʍ|��s��S����X�v,�R~O���j�D)�:��@/�}���6V��7���B���^"C����U�y�u��X�)D/x��g�����R��n̜��v��	�iPz�P��$_�bю|��m��-"�Ӗmh�\��UE� dY��Ͻg�1nJ���>��	��F5����0�;f_�H��}e��^V�W~/]��(�L������'S���H�,�̓^L5��6�<�w&iLռگ�q�=�{��1��|Q9���z�Ч� �8a�)�˸����6ZT���O�[	�����h�s����SE4+Rma��pهVW�+�	4*����r
�N�<�u�J��u�(��@�}݀Sט'��2��wk.}-�-�r}��֛+IM}�u@�4�bO�gp�m	�Lb�eM��Ҩ����q��<<�pw��R����v���ꮥ�@Jh6�-��uPp�.����Cv��@�64� �c@|�aW���5#�}��Y�ap:&�Y��c�ֲ�x,c�����O�6%�b5���sWQf�/�**{f���Bd�w?jφƓ�9m���ܸkǫ�~q|*���֛��2��v�NZ?�r���y
�qe��~�<���Zq��Q��T�7�����}䛻,��$�_�\�W����>1n���ΜT�컞�S��mf��� @q�ȝB� �q����1oѦB����GH{D���ޡ���5��_�K��K�м��oi����[�GH��,�'�<k9����텤����ywd�9��l��g'O�Jw�a}��9H,c^\�D��>^��Z�+Bb��k-D�0a�H�3�����+ ,��E4[�SDƎi�7>�������Lr6J%!k!C�6/wc])3���KQ��p���1�)�a��Ԕt�a%Hl�t��)�yk���L@�fܮIzJ����%ٶz�u�Z�����T�!D�X��Pa�1��3�*��74���%̋ZO<֨�8����h�,�k3,����Þ��[��v�O���&��n')���#����T����o�%�`d�6�7��[#��c8�Z�t3��[�<6wg��i�<�y��"��d,y���!����Sp������0N���qb����E�U��
�l*[�:�����4���2�� �_�S����� �ru�h"�tD�%|Ҵ1�"��5v n�~����n���/���. |UO�Wi	�~3��W�μ��������ϧf���-�C��/�������Ðzk~�X0 ���<�6��e�p_?������M$-�}T�����iw��6�\���g�d+��L��
��zs?���ߎ��?m����j��v�/�ZyW�w��~�+�wE͜�A~�
�`�
m�vz�P.OR�UZGt��M!�<�d����( 7��U����OY��Zﺋ����[bL�����q���.��mkNs��c���SE�홗.�e>�����u}Z�Rk�GW1��ɖ�7�Q�ĬAf��kTF�/��� �:�8�\4���Z�t[/����,pjE��g��s�A�䬎9�6����q7����$��*�0�D�R�P��驿�#�c�����*z=�>���8&������r2�n�ʋ��ǰZ���ۘ~�x6���y.q�v���|�R���e#��d�^�
Y9����ǔ��N�W-2�U�XSj~9��<٪����S�"	�b�ŜY���Zf_hoH��q3�Pnx���4zwǧ':@P��p@w%�V��O����N��U��!���+���BB1~��3vuc�\O<B�����)��0�-J���FwUXΤ���w9���f�p�{�
��a���4��[*����ʒY[S��&IY�8�6�h}4��]�'l#��9��~ P���_����@�0��Y&�F����YX/4�bOqL�Ժ��/�Zc��|�Y$�V�ZЎVŹ�>Ii�ǥp9;�्��x>.MvK�Y�����H�7vg7����hi?�#}��
.Vn�_��bJ��kQe�}�/I�l��S��i^ı�[�޸�"S�����;����(饾۬{ �9ߪ��+>���Yq�t뀹�k���6f�!݆�\?��@�����T��A�����El�Uw��fyOm��_�t�uӫ)&�Ǘ�D|�.��	p���=b(6sh>Գ�ՀE��VpJ�n���(�U2��X�sE��űd�K(�:+���bNh�q�u_�,`�JQ�X�Q�����}�p�Y8�TI�}B���}��#��X.x��/��,Z��i_�؆"�����V�tĩj��9�zWtS65E[.ֵ�ZH�u��T��yI�������}�HZ6��7�n?��Y�k�V��o#[7�ӝ ^ǋ�����u��1ݜ������:<`Jݥ# 
�J7�u2���y��db���'h�lD*����ѪAt?�e�꧝���l~��cQ���*�s�Q+$
\ �d϶L���g�yߑ� �U��g_`�1+0u���Y�&�%@�䣸������Lm�r�U��j�g���#y����>LU�����0f�=�u�\�f�	ۆ���J9g���xuu,ۺ�Hw�P����7��oOA]Qj1��DWl	�Dv�FR�"��xұm�Ha������]��PL�,q��s�c�<��f/ї���L�k�9AD�P옭 \��pq������dx}z�ຮ&.��n��Xw�"H4�u�^�s=9ݕh�Ԡ�����6�~����v�F"%`*�m�>^�cr�ԯq�G_��x�����,_i����r�?��ix[.�=��'���K` �ki|Ͷ(q����쏭6H����ِ	�T�f���|o��&�ɱE��������6��O�w�Cv���7i�;��Hr���2�S�n��!�r�y��:�PM�垮ꨠF�Q�D �ܣ�:nۢ}�C����ޓ�������Z*T���ȴw����B2X7�O(��S��8Ӥ� ���22���c[�	�s�C����Z,5'x.)/�(u���D�J��ͿU
grCq���aS����A��~��Z;[����U�)yR��F�1�<N�b���mMNAx��@���<�f�.�K�6���J�<ώ,}�rO��`�Eq�̍����G��-��y�>V��G�cN���\v'�t�j��o%1Q,Ծ��A��\$퐳c���Ԍ�g#�۬����*�y�/l����$#7��fp�����q���I�~]%�D��L!rf���>MR����g�ܱ��#�籮��qۏ�hXe���+��(%���� �HC��T؄�Wb	�%c�`�h㎻ֲ=�[��a����ě��Qe�������bp���z&#`�1���j�ƘM��H�KoH��� ��1�e��
L���J�2�)_�g)P����y�$7�^��A�*�(�W����+&��58t0����R�o�4��޷�"���\���ұp��)�i"��<=���S�8(������	���"� 1<����3lk.��T����3�`2 O�g�bcC;��0 �@*��s�KӸ)��8��
eE����AĚ�&ߔv�&ר��+�F1Y�%�\ʦ�Am�Ei*�\�i�20-'�}EN|{-s�<�����X�	�J&6�A"�z(`�N�[��E[P�ح0XtO��5b+<�$�4pt�>���l�w+�HQ����V�����l�.���[�gZE�������p�����蝍�2�
gb��_��QT�ix��iV�({�(L�{�V>��53rd$���d�q�$�NW՝�s8�5����Ѭ���Y�j��>
&��2�qUX�?o`���C�;��Ot4�Г K 	�� %���A�G�o���7�!O�B�����Z�pl�s�DՓ����\�r�]�WJ��9%�!ϲ��!UF�R��VO��������L�eg��\��8�^��^QfZ��R�nQ����p�CᄕO�Sy[�n��D
�[�h�C�Z�Mi������|Ǫ���:�)K�z�}���iH���tw~U(�X=��"yp�3d�3���d�:�{�Vua	����8{�p]�g����) 6�	�H����Bi�:�e��<�=uЧ��&��
NP��D�[I4]{��IW�k'��,oG��\'@d�S�l�nC�]������\�om bÞ�	i5�T�ؿ�>e�	�T�(*s(�H2t]�ZQT��d��[�e˹8�-18V���L��5uO�I����K���N��☥I�����˖����N���lafKFǒ�J��灄M�M��/�YĞ�Yױ�n����\�^�\���bj��5�/��C���z�����|ƖAG�7�cM�(WkPU(�F��� �KZ6pn}�Ŏ\�-78u}��AQ\�4��ʛE>����u��뻀�X|o��aJ��U6�u�E޴0���C&����1�.x�ϴZG�e�b��Ƈw
Ꮌ&z��RO%3�+Tɒ)�j�5�Ϡ�v��{N��Pr����������!���+$'��)�M0`�.`ʆQ零�UJ ?fƮ9�\
:�ۓ�z�$4���n)ah�r��i����rIu�o��v���U�-��F�00���i8�i�f�c:S� ��]�r������l�-Y
Fz����@�m>���5���׍�`Q�ǃ����0�O�j� V3$�^�\$fr��ѫ����"�=6I6�!��8]�)��<���t�s�U|f���.�.�RB���{�q��+����X3t�W�`��|TR]l��Tj��A��l9��ٜ=��`lyO�\I��AD�2}(�gpk��?�,U3-�K|�z�EN��X氭��GݓW2=�1�Ć$���jJ��:L��ݚ=ɪ�(��������L�DFR�UO�l��S�ɷ��g��[�oA������h���5�黦d����ӓ��9ٮ+�.����2��oJF�o"4r�M��J U���b�,�H��USGudfЬ����KbW�-BT�)2��y
�&<<����b��Sn�w����ܚ�fn�����H����^ӿ.B�lE���&�5� �U�Z?@���R�O��
]��X��#V ���,1�!M�E ��/.�8�7������K�#�9�_�^��M9=Y���4f{�<G��5���|=$
ޚ��_���gʰ���t$Ẕ���.�	�|�^��B:��z�G�"-�nP���أ͓��	7�������E`b�&��rM���,�:��m 4 �ՂE�Iz�<��뫗c'^y�����p�ľc� NK#�r�+>���e26&�Q��d��Y9R�``�<ԇ��d\��R���LA���J0nD��}�,���������11{�apnh}��{t�-����'��%9k,��N\���<F?��t�<f]|@9H���f�Ҿ�jw������36��{�U�x1Ӈ�I�������ᙤ(}�x�k���1B���
�~�<v7�#h�DZ�
}�i�\��kY�3�i�Cų��С�a4=�\6��x����U�&�_#@�������l]R*��V�\ *`oJV}�-}&�{Na�@U߀�`��s�_5��f������1z��t;^C!�P@�a��z����A��_Rͥ�i���$���S�X��_��6�g ������ d#�#��´���99V��&��hy�BAOy�O��v�W���}���0
��cՕ'k
tˇ5�#�=��xT��/�;	9��@�b���8�	Ê����ྎL!c6x�i� }Ȟ���=Ō��$PG�o#Ď�F�@�#���Y��=1�<��{/�d(��'Tc�C$ܾ�d�\��S��H��=�]���Ȭ��Ł��I������]*gk��+V]U��E��0�P=R�᧵j�J7�?�p��	�(N��)}}H�Z�q7�� Eyg�p�.|�rAQ�U+8������N�,��?i.0�b(�r9:��h*1'�J���dx���z�Ffa��1�<����]`�؝_\������Q���a�S9�����n��jE��|,����8��qoo!�U��۬t��!��r�����B7N��8��AA�x?#�wR�RH�Mο|�xħ��]aV�i����qhT@&�[��X�t9/cs] �?ga:��F�w�?�:�Լ�x����$�/��{��@��w�/f���S�t�⿼[�<��|���ݎ.�L����(�X�tc���a������=����t@}���s֋�=�������Kߌ�] �5��3fW���ܞp��=�ux�-@U
�v�W!���y�t8�6�A�	� ]��&}Y���#�}�_is��J!�0����>q��(,3�NbY�oRj~�mo��\K������s���wK����,_����O[}�������d�e9ut�JA�u$�?��aZ� J�;h磵ב�|�C���W�aݞa� C���~ԇ:E��LƸ���C��J�l�'���t5��NX��Z���Wֶ.Cmce�li��r��'eۓ��[�0F��*��[�4�/���cM�&�I���S��\��\H�1�hw��eђn�h���8.��2P�l����v��W��!D�L�Q��s��n6}!�nT�K���a<�@ǅ��ҡ(��y�u;�G}A~�d�n��d��8�
Q���(ZC<0xc@�1�����H����PbZ%6�Ѕ�z$L�����S鋽��\j���f�~�4���@cܾT�B�Su��v5��YL��H��{���i��ـl+��!��+�����%k�E%�s����h���D��[�/��T�jދl���	ؐ���#�t����ߥ�����0�5U��(+�"�k�J@��<����<�� I���U{�z��Pݴ��{��8�`�1h.�^���ȃ#J��ۦ�X��0��mş}���@�
롵���um-^�A��4��D�w�v2��>�>�n�Bf��Y��=kCZ��5�\�mp��nlߎ�{$V|��a��	��YhMB�PO�2\��p�d<���gb��#�s�*u�Ǵ"��= j���-3�-P��0�c�>���@�m?+\NДt��*�L����X�n���9�<Y��,��9[����+LR��[��GȪڒ�T�o�ZM���-��;LW��	̟܎6F��Ҙ8R:�m��W=s!���<��C�nJ��8f���r�u0�-3~�=�=�,5�EO�u�B�&���:�&������ϣ����(Z�>�fm�"�R�q���R�ӳ��0-���Z�K+������)�s���΁�9$��b�h!��_�FPE9��e�e��@f[��S 5o����I�("�Ҳ͡V���"|�˽�u���ɜ���~&�zB�FX����~�dw�.ofE���C�q�m,�@�!�7�Q>�ng3=���{ ��^o �__�����r�ĸ�����B�a�{�������VGO'�4�ѵ�O	�l=1�SšF�pa
��R�@�ц%gX��k������8�Ӓ*Π�f��5*o��&���I�-��`����t��H�H-�,=�]p��DB������˝2����X��uRXlڵ�[H?�&aJ��"��C�MJ���hKd��f��L�K��K�?݊`��\H��ń_s͸� ?ן��m�h�k;x���u���.U-�mw��2�Ũ3
�4<c�l��;�>���pi� *ˉ��#�#����>P�XI�( �?����qBD�)��CM�RՃ*�MI7MfC�8X{0��=�|a|@vC7���,`�V?;Ɵ�H͢���*M.Lci/\��C����V���p,��1]�l����V$:��WG���eb)^��;�%oW�/��844�Td�/5�3:g4�1�<�X�y��5�yR�{0/.U�[�h���k&o�����p��i��ͻ��Q *����6:'1���4��Gj����憯�TLԵ"Ce|�D���⭟�ArDG/S �ogl818���e��_�3�V Q�y��ӄ���C3�OP����(u����&%�;㺣��}�8׺�u��ؗ��@SQ1��x?w)A�)t���_��G�����W���'�&�ն3I|�0d1;X0��b�e̦�[+�S�D���԰������ޡ��7��d�������΋~��P�����k!:9w���y�g:�w�D�ܣ���������GzЏ(�Le��)�$�K֏��[Mkd�*���H��0[�s�6&()'�Ԇ��sq�L��vpO�����R4��C U�Fil�MP�_�]
}���Q�D�&�UvYV���5�X\\Q+?�$�}�L�wr�M�ʓ��jz�m�eu��1����,asy�]d��Y�\�-_-��?����������_�l�� {n4�`��<�J�S��2H���8Q�]�+1@��ʟ'(%Sm�����ձ;7ɪ��,���2�d��0X^.�q�2�m�"_�����|�F�`� V%�������dPk�/�l�9Bū8������F�c���a��Y#Gtz�
��&7�*s��$3}ٔ�/
��`��j2#5�����{����@�kKм��[`��;p#��g%;'�z����$�<�7	�Ek9�4$�&W$���9�[�KX7'4�� ��.f����6O5K�L���a�Mc,�TF9tە�ϐ���M��;=�*��^�2�m�7�>���t����EK2���O��r{��-�*OZ-��chNj��'?���"IB���阂�"�P�F1+�<W���0Ϫ�����{p�����Ǣ������Br��I9y�qsAP�-�le#3�
����;z���p��[P�k��/�4lxT��&�e�2}R%�)��� Q�,o�C�����-��I���]5'�">���S��l+8����a��Co��u�$n�=Ky}#Јr�#�D@K�*Wut,q��v}IT��fw����2��lM5C>݅\ܮ����r�/��8um]��;٘f�.��7itWVΤV+�EJP���zj�<���&;�hh�g�h'�Լ�[�N֑)�7��ɇ�D��Èؽ����]��e\�aGh��M4(5>E��B�2Y�����o�&D��'V�G��O�ﯡy6������ҵкhf���|�#��V�<���_���D1߭t�B��Kh���L�x،���t�\�r�d���P	���{�٢��3gX݅����D�������#;E��X;7�B%?���V��h��贿���R^�"�R�PZ��
ك�r[�6R���Z��zeG:i��>�Ci��A�t��*������?,�d)9��0O@~�Dr�%����7M�i����ei��(]33�����Y��e�k��`W�i�Ħ��TAo�}0�96��:%��!� L���7*q���T� ���v�U+!���bڶ�m�qн����G �ƕ ����n��� ��
u ux�S��i�gW/X��]V�>����{���UQ�o{���!6t=�J ���_
;��Kh�i���Z�m��g=йB�U�T`6�n�9��-!R����x��n����ќ��x1V�tw�b���t��ʐ�i�.=oe���t�W�~�`��t-��7�_��� ��(f	4�86�QƱ1�&8"�nM��Ч��,���)�P�<��s�'"Gy� 2���>�	w"�`[UyL���^=x��7d�sj�|��+�*l������:�:'��z�c�m�tp�@�)|������J�92:���>0u���W�i��pD{�f�����j�N��E�q^*�-l0i������I�O�j��T���,�����5E�e����� ��ۏ��y��ͧ>���S�F�<���m�V��#���d~��ޫbͤ��~z'kN�z`��2�ٓG0od�p������T��Ĝ��FxmHm�ڨ0tP�z�b�������>*
w��p�1D��G�
y�M����u��x:��n����ь��ֶ���`^/8~וr`I�=�m;���}V����$���{`����}��HHy��"�I��'g�{5l!�e �Nwjm�;*^Сh�w����������6��6:7ѷ�<Y��;�`�%��>�㑌
�6��U%�)@Z���^D�9��VG��)��0���]_�`��Ad�X{nF�|f\�(��)p83a��P��\�ZzY�Qp��qc��+�/"�0G��&e{�ޣ< S/K� ����n'��a���"�8]�|F�,
1ݬ�e�u'Z��t���)¡k^X /_��͎iu�����;��u�^Uf������ZmPG��Ba�q� ߾6'�U19?�!<� ˨+&�g�;8�����4�*�������&�4Жڝo�E�+MM��Mw3�JІ��h\_��0�"H� �[��k\���o�A�ک�dI����pYibeAb�X�,r �?�t-� &��gX���`o�Ҙ��%ӸZPQ�6&�dK����;��ޢG��蟹��y������|m�8�Jc���4��^�״��M�W-m@�IQ�!i��d ��^"���Di)��^��}�ﲽ������p��ڇ��&c:$�c��#�S��)2)����A5",��U-b�x�����<`�H�*~��y�$���k\���!����F
8A��5V�3-AVȄ�dM�]�+[�9F9��b��$ �v{ǭ�Z3r�!��"&�r�4��#4V��L�D��\�w�.f5ƞ.=;�Nq=%�h8X��ȩ���� ֡����q�2�#.r	0��B��I f{O�o��;�D���9B�K�}�$2�hu�Z=K�~x͟��+�G��Z�v_����Z"=���fJ9�,��O�=s�0�Ĭ�`xq��G���$m�+��~�^�(|\ (�X/���4������#�E09מ��m�;(TrPV�Nf]�����B���Na�R��̍���Ҿ�FשI����:MV�d$:�����LN��� �ճ��Fձ>d,���]��i�qZ�e����"?�~���G[7�q�uH��l�h��6h�-�Єl�&��]�}���N'�Gt�'���e��5�ڐ�d�2y�|2W]|��z+�����Լ��I%bT=p�JZqPs���#���t�r�|)s"��*��L<��!>��F��U�Up=�����W�v���-��E�h,�?{B�
+vyM}����l���&�%X�<��!,ONP�� L�W&��?�׿}2ky�t�i��F! s3�6��7����`���ǩtF�����;1���$�v�\a�XQɭ�f���=f"=hʩ�uؿ[�z;�!dyCM)�<4���F�1h���\��9@������ɪ�J1����Jzg��VS�b:�>�T�X%w��Hg���`�c�		֡�q���ޅpU�Z�E$˨�������%�HS/i�s��b������А�Q��+��Y!�׺Ѷ��S5��>�x+�~�RC��[�N�{M]�����Å@>{fd�Q�����LbyD����Ӳ�l�1�Yz |��EJDDgq��y�"��A{�RjR���o$��z\*\K����@�rc������M�o��Fp���k�B)�����������y(t�i0�T�]}$�@��J�����΅i�.���Γ��o�#"b׀0��rh��y�3����xP`3�ʇh핉�`vCV���.@��1�M��$��њ!��4��̏!+��N|��F�(���M�NƠ^�1�Y:���f���7�nx19!Oo,��yH3�ȳ��A$�j]/�9s�i���DI{b:������ⳲoP�hT]�I3F���yL6e1�u��b�ѱ.[���n}n�ϴ��'~�����q�ՠ���V�"l��租`JY�桪)m7�-�v�#~�l&Z�n{5(=��Le<>�9T�7���^s����`�G��������a	�i��t�����QG	|��-᭶<A���2����=�g\T��v��=0�>0y�����L�9���IfrY�z�h��/�"p���$k!�m����j��j�l��Բ^l����Ju�,�?֝�lw�
�V؟�EM���-�i<ֻG���
vSז��8:��>&�2�n���&E�\��E�9�%��0*е�9W�i�{��/����GO$�%��1�N	M]�͊�P&+GX!�b�mDK�n+	q��\-23�#4��>r�������ܟ��=?���B��C�mTߜ���)�]@-Uf9���¨\�쿺��$�B��l^�8��L�0Um����� bB���Gh����m����	��`�&��Rtq\P��9t$nze��U��M�����ǉ�Nڊ� �.�Օ����>e�	���S  r�������j�uvLC�lz�#�6�7ʓ�&i��,�esG ���nv�1���$Ρ��C.8�շ�mX>#����
�C�S��<\N����<��������#K<�����]��~I�:vU��U��3 �����,,i�� �-�/��iJq�3�TwPn06Fk��"���7`:��9
6�u|�>�D��l.�s�t�0��.v�U~w�LI���|��_9Ęe�3
v\Jj�~�M�.�k˱�q��M{��}�.V����@G٫P���Osw���ǅZ�s�O��Z��	����P"i������`0y���]������1��UN�����<��+���W�ö^ڷ�VTs(.�!{ޤN}f8>�	�F'㥠�둑��tW��PԹJĔ�O��r3���ky=�+orp�J51�L82���KթlU� �.���l7�JJ$��__����+�����j�5��+V���qa,��	lq�aWk u��#���<8�u�&ߌ�4�k�R GԀVPk$a����e�6}��?�F��ۍ�B����]c�l�fa�6�Ԓ���raAc^��|s �ӆ�-��e�V5���D�s�2RW�zf�A���3}Aʱ��	��X�I�ȕ��8ۋ��u��L������R�/��z�t����~�͗mn��݊Ċ:�Z�.�9��.4�a�R?�>��` �v�6ꯉ�u����`o6r�Ad��@]\}�_�u�n�O�/H�?��Sf+����x�u>gi���7��s%�r�hM�GS{jV�
��Th���s�a�kU>k���h�*����j��s$�-,�S �rd�M�XS(UQ])��L���}�ad���7\�!�4�qe��.�Go3�Q�[��Ge�v�0h�WIB�D��(�6ؐ�FK� ��B+�$�4�k�|@������F�sS��`k���H@a���j�����:�Jw�O��$����܏�m
���q�dd6n&�CO�</��&��'~�F'Ư���"���
	�nw�݋OR:2��8.|ʅ�V?��1��e��V��i�����<�A�0&$��L+cם{^)��ټg z#I��|%���;��bl�ű�7�{h*^H��\ �����}��KJ+��\�Lȝ���|���D��"qK�L)ׄ�]K>�@��8ʨ����;��X�T��K��K*�����U�f�^Spz��j`�#��g�=�xEk��g��� n�^����erwh�[�]b��?0��R����s/�5�	v�l��Yr]�'�J���y�����<��%�~\�
\�;�u��L�T  fk���n�.�}�f3
�Ҡ�&��_ݧ�~�M�����c� @����boCn� ��R��Y��y�����N��IVe+�)|4r�Bt8�Ga�tl����Z��\��	۠��1cU�Ih��X��IV�$��0}l�P<;�'�lc�9{J���	}�.��f/�I���0�p�NU�sj����F����6߁T���/��A=D��������5��>m�@��N�����O�A�x���R����I��]��i^�� #A��������+r�0�?L);*��%����S�(,��TRg���֝"�$�,���������FZ������f��	y;����4�w�R�{g �z��o��ڝIS�kp�_�J�<L���[BĊ�zC4��Y���!��؈��[�H-���(���9!pa�֞ga�����u{��Ҍ_A��C(v��&kɆ0�ґ#�3��1���6ph=��]���qE��u��!X`3|�1��	��Z�~E����(�����Z��R�'��(`��`�I�������U���a���ctyYp^/�K ���E�/%f�t�H�b��Y!�-TǨW������2}Gn0{���7a��ǩ�V��x�'vs#F��ap载���T�1�e#h>�:���K:��ˬyBS�m���K`.����{ѿ@�^�B��5Y�ޱ�bR��E�d�ҷ��xn�ec�U�\�� C�fh)�y��I��Be˛�� �TS���Z����q���C#]��%�S\�	9_��Ĥm�&��(���u�9�R�jV��[���"����A��,!.J�SUU��,���D!'�i+��A�?���2�)����@(U�N�f���
��А�l,�)`+H���e���K7����Ʒg�H�Y�L��Ղп^��>e�qI�)��t�9{���%����G?I+�u�a�8�/�x�a���=�ǯ��5s�2N����Ȱ�V"����#I��C�U�S�-T�[F�2��,< H��&�x���w��cwxA�*��F�q�����aj	��J�e�Gcy!��qz�W~� BM�#)�{�J���ND�p�k�-��#�����-�F�:�Pɬf�����H	`�v��K�P��YU�y�}����hi	���e�����Oc�X��'!�P�T��DH��D\~�����A����ԋ���b��=�(Pb,�SED	^�6��]�Vmo'j���oT����AɆ����ڐ4�v#��>�%���R7�6���Bjb�@M�=��H������;��7mO�oj���E�?!ЩF��S2���ga����р�2G� 9�q�0<5AjD�����+
�"�:�����|$!�Ѵ!��w�)>���cw�>�8�L�s�y\i�XM��U?�/�1����E�.-^m�p-g���;�ALp����s�����h̃����&�jè������G�	�u1�F2�.����MFe�Ӄ1(H�К@�G�sq��@�0��h<� k�"4�צ���uG���Ѯ�]�\
 p��&P�zr�}���am�B���=�ԃP���\�Z�l�<{r'��ڴw�D�䘵Ħ}^�?1���:)�6�j����T+R�	;ZKƭ'��#3����̝ݯ��7`�a��jU��Q����B��P6x��&j";��oZ]�[vB`5�4E�j}R���5)�n��`����u�,�(/���'��'G��h	hƆ	̃�ʱ�t��_G���na_�8'S�,5�����We��Q�ܘ87q���C�ݱ�|w��2@�������"�����q.R{���
��ll(4�.����|�˅�<���;�P��?�J��l��RE,o7��P���&ߛ�\�JNȝ����%�R��R��7-��	BHqZ��[�������*��gs�dA�RI��5�FCw�X�7dUP������@,��q��T�/G�M��m���CAH���yI���esB,E�ھ���Ʒ�U����S,8N���1��hD�
4���N�:���F�����Q�F���F=�����˷��7Z,dJ�&͠%�F�Z�RI�����o�ɹt��V�	���������Bo��e/�=�I`E7�*C\��C�Hf-I����%AА�o���Ls׾�#}���0��J!D5��1�o��`��/C�AfJ�Ik
�N��\r�@ߊ�Dh4��ƅ�_U������^Ze�������ݏal�Z�H� � ��q�X�Qǣ
���v���b�g0�o=��ÑH��p�Hgx_Do@�4<�#��?onS�Z�$�d��a�q(#0TɌ|����w�{|�8�e��ZS��8�@��
�}�	^�ŝ�0#�ɷ�?x=� JwY�f�G+�.����"CV�M��Ê��v��F�m?�R����jΆ^��Ȫ�I�+��y�l�g��y6��ۙ��ߕ���'|�,����}V� ��^e��t�/-�f��S���l5B�y7�1�z��%���,��ϸ���[� as��E�26�h�����l��y�Ay9n��݂�Jj�&�kk��L��&��x�9�g����f_G��������͇P��.Q��Y(X-[��D�. ��:���<,yV~��f�_�ٸ�F��끟{�qJ;�ae�� �y�8�~wQ+��1���;�g-}D�������;�	G8i�:��ʗ�n��S�����
�#����"��</��n
�<� !5���Cq���L������.�!�b���G} 9�Q�#Z���VgS>m���G;s�Ğ�Y��l���-���:�r��5{̪�@�GvSm�	�d�N1�,�5d�_��s�0�c�Y|��C���!"�X=�$ͪ�0��4��h-�1��ص"����^���z���8�E>���X�I�ҽ�����艶v�#�Տ�/�L�X�d��ej�-�O��&se/`FI%L
ᶞ'��(�S�� ����

��Ҕ*�Hl��!�JP���BX�bh�D E��@��u����8}����M�lVSUk��uA$����kH��;-��M���Pyo'���� �	���ɺ��5ǥc��hLG=\)� պ�\T~<�G�.sw����Xb ��)
H�׵�^mU�| :r��A	�Wˤ�]uȯi�Q��4,�V��4�/&-��a۔��w[�9O�yg�{�$�h��ӆ/˨�Hj�;��p]CH�s/���������N�Be/'}�����$��V.�� ��u�f�m�{[q�q���Nh���V��2���Nz�8�c��Z3���J�x���p�8)�F��~X
�5���u�����&/�K�<  Cm� ��M�0��x]ΓZ��N���]��*�5ܕ��O� �-�!V�X2;��;W��D@F���)V�Uk&��Ԙ���?�A>�S�'��e��
]�!9��2�m�儦��O���\��Ч�B<Y\�r��rs�
~���}��R��ӏe ��ڂq|hG៓G��x0�#">6쾨�\SO<w^'`
M�g����CD�ʴ~T�"n.�
p�4]P!M�;*ɗk\�7��ѽl���C�7�'^�����ksq����]Z�@,C�"���nÇB���o��S�7�C:�+��x�W���CǮ��(���!7c���<p�QM�9�ku5kh#�����X�V�ȍ�Ā\tA��sJ��I�=�Oƅ��Y[��¯�q�YrNL���N�f$�Q��.�!��c�)�ŃG����"j��\#~����m:�]e��J��J�k��0ܱ��@��r��"�	�-�F���7�Bn�o�1�9�q�Z�[
� ��G��Fe�� �:roƠT�.�3 �R���;]Dp~c��L����<4�	XY���G=�	Dm�W���2�S\�L<"��-6���i�f� X��4�)�H�����JOm�Wj3�A�oiq���P��iEc�����6��c���@z�j�w}Bn�x�����P� ���=�:w�/*���A�Կ��QW�	��OH~�������e|��O�"'Ю�n�`ҿ�+z��{���!�ړ��S��n}T]5��/Ky�xU�D͓���c�_�bB]Hܺ`Q���wS8���`6��Գ��ڑ�����:�"ə���x�=f��6iQ{(�j<�O���1Tsx�=[\���H@u��E�칄�mV��+3M�'�Ԫ(Z� *
b���'e>C"��C#U�5n
�ȦO�޲bN���җ��%IP��s�gM<q#A����hŷ����Zb�v̫��7��?Rٙ�y*^Ӯ0�C{��wKg�� �&^]u�ނdv��7���Wc8���?zl���	�����֍������TKH}uX\�J���+	1������9� F�UI����7��?b0�Z���9��s�g�z1hh�� o��_'�w�0��[��~�7��^���\Bc�_]�z7�{��ƈ�p�K���q�;� �T�TA�ڨr���7�\x ��հ~t�N�r�x�h�~Q� ΢�p]���#H�-�V$|��H^ab�h0/5$	� Xu�כ�^��� ����z�R��=�� ��i�o��m�5���g֭-@�N�m�
�������ɰ`��%��M��HZf�K��ZՀ?��n�!^�MI"�>�!N�Eܜ��,��}�r��`�~#����'�������v�7������4�jCR�+�%#��,�4Յ��T~��~��D|@3sH��ݠID��f���[�mg�����\��r9�kJR�i��K����*�*k-a��g%9���?���"�j, ���8R7���i[��o*���N^��Uj.#&��D�ڂ�؊�����Ȧ��i���R)WP�iq8s�&��7�(��StU�Y�g��P@-�#:㟮+௅c�6�)i_��hMv.x"`
�ʨ*�LY|��<��^�+US�!�S���ʮ���S��o��&�:O�(I  D�b�pƩ�E����`�n���� ~�.�>��S�0�_h2��(�~����dJ�E�����
А�j�9KJ��tW�L�(00ju�o&�]�Q#�& L[���>mS�>�a9���st!u�ivi� e򁽒���{���"ڎ�g���N'[�i�n��斺�k���H���_�Ɣiީ,hmZ�ŀe��׭�)����F�)t�߶�Քs�((�z�A�
�Wz%
ږ*�#��k-���Jo���D<���&�H3d�a������gm9�h�gSN}w�R����3M������|c��/�����x x1���.� �� у1+���D�qp��6�����tkD����b������,�A�4 <���H�3OYpHb-'h��NA�P�y Y�u9m���]�������tҚ�#�;Trz0:��[���^L�lv>����fF��~�H�{0�H�Ƥ�������a�2\�V>+/]�<`�Qf�O��!����p��'�8й](��P�����h9`sY���~l�q�����UM�ɀ6��8�ݻ{*G��_����,~� �3�C3���EM����oY3&���'�W9GxF-�8^�^��y��Ǖ��>�<�8g�	� 5�\W������Jp��{��<�B�`9ݯ���~�ܪ[�-�rO�4~�z�n�Ǖ7e�rY%����.�ˁi�O����K;a�� g�w/
c���V�;�x�.Ex~hj�K�j���3�'�1��w���(�Z��2�Lt�����!��n<�kD�Ԕz�-��{�:�{&t�Xp{H	q�_�`��aa�o�)���j�ʔ�N�}��T�6��a��*��:)�&������f|���������>�W����lC1�����~d��o`H���z� YĈL�����|���g������C�6���;?wD{���c�O�|��や� �B�ڎg��Ta���mt�l�>��B}I�E/~��}n����t����E�
�X��9�2Z���}���:�켚!�
�@�>����������X0�7���$y�>ۮ`6�o=t�5w~�F\�]>��1{�q�	�¾H  `YZ��1�}iq,��G���m[.�q�i�0PK�^��&���G�np�N.lR-4�NEuh��dV� yM����(�H�.\�Ev��O��UL��Ȩ{�z�o�y��E�/��iD?����7��S�'9���a`�� j2�y��˗<��Ɖ�
+��L�(5�f��ns��3nC"Rv�t���欯�Y��,�㥜�Z3%����u�sg�Y|�u�CDBy�ws�9
� @ň�ɼ>ʤ��0mт�7ԮYh��|��E�\�� i{�)�Ԛ���2�9�)�B�#q�@�?"i'��u�w����fwk�/ǆ:�����2Z6��8\Tj�g<���$���-V�{�l	j�ۆtj�y���ph�I��4\g>t��<�ktT?9ɭ/�Ԓ�6�7;|���G��8��L:2x�0�s�����j�d�k"��C��z0*c��)�@��/����`��:~P��������E�
ۃ{�Hn�l��V����{�0*���8�E?�q;Lͺ�~�'�ffc��Ь�5 [Ğ�7+����\\��o+�^�׼��������k#��X�E�[9��>%�"�Q�p��b/e�r;��8,4��[nۜNU~��l4ùr/G�%�63�ت�梸 �ø�٦I�c�����.@�f��2:9��ya�����"J�Da_֞�:P�y�B9Z0���$������@��D��λW��ܖ=(�d�T�0����ї%o��A��شM�F��Y��g�5TG��Ȍ��@gv���K �f�T���~I��
+��')`T�r�ս�9je �ʖ�]���=�qy��|�w�9�v�]�$Lq�}�Y"Lp#9s�̟�P؈���:@�w�{�@��2i	�gU)~R�4��N30��v���Q��f��I��G���W��۷?
��:m	#̷��[8B��P׻���^#�����S�����a�����e���h�����@7t	�u@�2�!-Z�!�"�B���+
9F�+I�)���������m����v9O�E�+R���j����n��Gء'ͳ���3�M�Ks�ӁP[s�?��F�2TU�7Հ X�u�2�Sc)Ο i@�Šh��k����?�gC����z�y	֒����;O[�`�Z�W�O���g�p�LI�V�
/�@<Pw)+Q~�B\�X��da�#�ns�UR�� 1͋Q吟�~�a�nxi[�+?>2y�,K=��tgn&��d��>Ro;�� �Y/�`A6��`|�[�HӁ��k����`�P�!���;n� s�[l/�����9�R�³j��~�˄-׆C�H���E#�>���NP�BGU���e���f4fi��-ǩH9�h��U�g�2�6��!&�p2�8�����7�/�,e��N�!��V�}p��l!��~��@|�Y$!�
9���1��ay���<v����R����i����1 3
��_=8#�r��r,O����j��1j&Ipfb/G��-���[�X��e�9�����ZG<���t�{��cWBU�2Vq~q���4b?rvdi�aZ�7#Ͽf�qB}�� ���&�]�_��dqM��˸3���Q'�'�? �����J�GpJf%o��;'f*�=BK��������u��PSV�+����]��ڮ���"��n��h����@�m�+3�<�3��#�a\;����2�nFɭQ��6/`�>7�M��RN��V+���Ϛ寧�+5��鎓)@@,q伫5GC�>]!ʤ��D�Z
��7d���m��<�J�P���3���x2rs�/B|Dس�/K���rI�/�&_�����Ke��.����^�����aQ&�K;�nBMZ�|E���ݜ��̪p����}Ed�	r�ʺnq��-�i�Nw=�� T�q��V��S"��J+�?�Q�lE��!&ZlMWozJ�T��V�~�I���~A�K��<�a�̟���&���y�0z�&�`����G+��^oX��&"�������i�9V���k�94��ZQ�] `�;JK�z��S�H_7:\��z�iHv]C.�]��V�jqć9��ܶg��-�������;L�*��6���w���$�EUJ�7���̨��ș�֭g��}q(i�_�~�xr`�����J����7k�J]�#�Q6S��K��2]���좙*2�A�ܞ�O�� m>6N��2���*���Au���/��P�^��0���<O' E{gd�
�R�@�6�E�v]��2lc->��>�iC�֝���ЌH
]�Mf�$�*��<H䕉���,�f`�ݱ��v�z����U�f�b�BP>�Na� �D�1�|�#ISKnZB�ݏGp�C�lfd���=Z����K"%cR�z��q�FA"'��~$��?�le�ը1��B ��"u�@�^��I��H{h���D�x�����o��a�[�cX�})NQ������meJ���@[�CC�?I�e�L*@�
O�j�#��9�ҭtP�&O�M�\(�Q'y+���t1�\=`A萳��}��ե�ߛ�Y4Z�S�C�[���#��m��E2U.h�0����씆�;ME�>�k!M������*� �EU�|-rSe�%�u9��q��kB��Pb�x7�`d�h��k���D�����Px7����{�^=�y��D����7B	� ��>�����	���x��������r�e�w9� �i��U&���ڊ�}����H�3�������(���5x�,'�r�8N+��D��I>Z�񛵚�;�~��2!�Rf��2u&fq(���>�/g��6k)1s��ghm���w�rc���}ck�����Hp�,�H�,$�V��eo�C����$Wi�ezK��h�i\��y2���a��x����tsٗ�(<AW�TR�CV�q�w%5����!����9}MgI����W�0Fo��-6�R�q֭���Uw.7�-,i����>�Y)�b��w�>�	RC��Y�]�1S\|� #�-9����J�K5��ZR���biqఖ����{�i�\X��$�#�����E+$���ÆQ�D�W!:�>��i����f�u�Q���֭6��/X��/ˎ�ve�:��͍����<�;�Q�js����;�3�!�"��#������D���3�TTP�0pJ�^I�E
(�|Z&�u-s�2��%�hY�'t2�]P�2�5��O<h}Y_	U�di����#cR�%իl(f���3'pI����V�6�@Nmj6��M {<��:a�-,����9�(�E�Tf+�SK��Cia"M���E��)�M̀���&~~0t��/֞c��5���]�/���s��i�Xw΂��*bîU�UU}��D���3��|����E
�7A��^�ԹL�Ac��h`��8����M)��FlPH�� +ωԋ5'Yv����<�XZ��[#[��Ē4C_��[�b6�����wVL�'�&�+%jC2/�ok��̼y��⁑L��*�Q�
���=�zV�@��9Q�ϕk�VIo� �ᜁ:f��O�|�3bwXk�t�4{���y�'��9�<��9W�U�|9U�;��٪x�݈X���5���B9�ѮEI�)��6�ׁ��ٕ3<��������QX�(HNy��F�ogK����kL��_=8
�K	Z$�J/4m|�� 60� :�C]����=��I>(���y[��B��zhv�_��W5J�B����1(�|ʈs?t���u���6�)��⛞?l��T���m�5F���+h툫]��!}��R��A��]'n�9��!��a?�oY<G�.a��(�42p���VlH�Ѓk�P�Wo�馅�Q�j��ij��{m�8��TU�v�:�%Z:W�Е$�z�-RɄ��9ۃv�Q?��:'$R�����X!�[����#��Ï�h$h/KC�+��0�B�h���D�B�8=F�D��F����כ�G:2U>Z�,P�9\��A��\g�������G�ct�&MVx�*����E� �km�7�Ǆ�K%�#'�a�˪��NG�o�u����^e��;w�;׻�����x�o|Y��Fݤt����_���t3��lU��s
9��`}�7�V��EQ ��Sd!�E���?�XJ�)�&i�c��%��B8�|�N��Ó��*�+Sp��^ၟ3��9 @Gqj���Ώ��B6�K� 2�sQ'Ym���R|@��U\�$<B�<���ǅx�s9<	��PЁ��2�c^�������q��EN�t:#�#�~���cn��M:5���!���C�?0�_
IC��ҡ.�F�=�t���р9������0�uH���Z���[QG�j�{���4�TO[�_��u~思����s��X4%��m�t�E���j��E;.m+W�c,��3bA�p��{Kz�X���������D�dwXEo�e���^���f^�_hY��w'ﾪ����T��V@[As�e��A��u��v9��Z�Zݡt�)FDO���f��|�������?�U����F� D9�����KC�x��7�{��s^͟�Db�:~����i�1O�H�%JM}��ʀ�1q���0hTsr����������K�������S�f��1�0�e���ͩb��X`kQ��:��^�3J�X�)����1�A��[���:m&����"��h]P4���N�zٯ��SM�d�v��¸�}a���2e�=�ޛ�9��sL��u
����ڊo�_�Ke�UFS�-���Ҝ���ª��xp�
��{�I_;�0�8�%m���魎դg%����pɫ�
Y���̄_?ɋ�6��B*KQ�U���Vb872A�Ic����U�΅�v���'����)�˷�Oe�5>�py����%Q�ӕ!���5BL�P?�I�&�����})�2hr
���f^���g_�P1x��e�g�釶�2f��Xӻ�w����8͸��"�?�"�e�Hd�d0I�:��sVg��j+����u�R������N�/���h����L�u����u!|���5e��,����`�X$�f��dE�2J9�P��N���qe=�Ti�a�0<\ǔ���k4�A4"�wq6��� ��H�����!c����o%X�߭�D��oZ�MJ	3�=߈���o���5� K�\�n�xW'^Gs����Eܑ0��~Qмr��n�7Oy��*�.O���հK�:� ��9+��"k�����A4�:MF]�>�I_��GZ�|�9����%�����X��s��e:\��=�H�,��ڞȯ��"r���^��`a%&�7�}<���e��s]�ԗ[���x��u�P�P��A�ݨ`"��]�a�ɩĵ��F7�`���#�^�O��{��$��/no�E���	���-u¡T�A��d_����̒�E]�/B���}��J~f������	��O]`�r��_U��e�l���Y]�]ɰ�D��]*�ý�H�EAuEz���:��"��M	X��a�^���	`��9��JiD(����a}e��V	�S��}<7����{e�О�i���y�n�� �ށqd�.]�S�D_��җ*�Y<�G�"���n�6��ۦ�DP}e,�H6m�e�eQ��\Uw�s�u-&�Y7����"V W�_\�ƽVC0e>���4��W�ӛk�6P`�Ǘ(P�*}�ЛӲ{c�Tufu"��9���g!Ԓ/�L���T�[S5���}t=FF�b8"�u}�r[5k�zL���o��Zׇ�n��7�Р-���~sB ���K�/�B�6"y��02J~��[�DQ	`Ŏ�c�dlNr+�Uw���s�(�5"��V*#���}z��9ۻ�]�j�*8v�o���ߝ�m�������+�����q�z�\���\!�����p����6S�1�龾��K�6����>y���v(���K��ʳ �5~Y]�!?�����]��B���bdT�+y�d�'���P�@Ҕ����#�i���J�z?�T^��4�.�FXbu�d���
�?����b�Z�q�f��b��M�J����Y�jN+a��*��/��$�O��#bfN��>�TH��}�Ӹn��*y��O�/�3��|�r3�ɽ���B��HT�`��i���Gi����)x��,^˄���n.��?�8���O@�F�C*`nsH��A�Xm��C��<��M3�����N���Ǜ	ȩ�g�ɍ Vi�gO{��4,m� �`#�*P��T�=����!|,��8W�#B�2��ʳâ�[gi���9]�Bb�7Lt�#���QU�Z_Tta��h��A-�� �cg�i�~�:\89�4�W=�>1�I��@���h����sȧk�𪣆�qR�,�G�~1d��D#w|�8���#<��db�&0�}�4d@�������:����9�:��h	_4orm�2�`�|
�WL|�	�?nT��־ШʍF��_�?�PT��т&�"pK��km�y����W%�Za�;���^�9#���bvۈ����گŘϭ��]��$���cHE`Sr��<c�)�Z4�hF͑�L���%}� �K�
�'�!�|Glf���m�%�~f�4�0�,|9��wL�a&Z���|=�¿��& �;�ol�_�}q0�ɲi������|k��*m���I���<���i��XԽ@����L��at��7�¹�	�i�v@L>i��<�Ѻ�8Wh���_!�C�71-�q6��gʒ�g�cD|���u���r�f�9Gf���E]L)E�fz3��Qd�n�Xן��T�3�� [����"����Ӂ侳�	�F/�#T�,/�Tm̟�9�p/��L./�	��ysxg?�<�
�
#Q���P�r!�bm��mi>ɥ�	A��%���쇓g���>�k~z��&����pJ%w�2�y*3��Ƨv��oa����d��Q��d���_�آ���5i�����������6(�����XJ� P���O��'�j��*��#�d �Wh�$���5��g�2���l|�}ԏ�Tb��/�5��a���E+?)��Z��a�B<�	�
�=(b�~C[1�P�mybǠ�ρc�7&J�[)|s4f驶�wL�w��f$(��(��������i.�4^�Y����/7jh-�#�jy���t=q���hUY�W��G��,�@UʅG\��_���e�0Y�*"/om�!�����N�8�q�>Oچ���S�/��۝l�9�ۀ�tt�%�ҥ��%��,f��Pi�y[x{���S����X�p���: ߔ����p*!�i<cw���da�C��3i��`>[x��Y��1�e|_�{C���4�����}"ym;1�P��
<q�ϩk1��nsܺ�To˦G�0�[�u�>B[�nȸυA�Y�L�DAS<>\<��������:I}�����v^'ԇ�����.v�>HKl�m�*jZJ�&�H�I*��$�t�a�с�T��0�3/���������M ��C�?Tg[��i"
lCK:+yUϱ	�$TpC[��#�N�Ϳ("�q2)��
�w��D2
���3�����7��x�ތm;N�z�yu��G�Eb'_:��_�HZ+�����R�Ƞ,e{e��w8,v�Vi�����	Ή�r0�6�;�6Zfp.Qf�P53,_p���I����夹=��p���J��;6�q�~3T��[2**�kK}��󽰹�Rn��D�E���,�z�`��#ߐeh��Y�_*۫ꬤj�S�'_im����,�?��͝z���(�Ji�YW�O���X~�	�Q����zj���k������y.�r�ÅJa����m\�I���i��b�Bu���AIA9�x�Hd,���xL��Y�ڱ�.�:�V}�(����]��(�_��|E��<���d�ߒ.8Ht�ڗ��z���˟�9�!T�}�(
25g�����/B�H-�o6Y.�x41X���]�?���Zm�!%����t�"�5�F�\tz�4���o�B�
��#$����ũ��k ��xL\Y@�:��Ң���Q����c��RA���!
�9��\��E�����s�sGVv^b�<�-(�%}��I��v<�]%W�i��_�7Ԛ���}(&A6X��$CHb]��bU(�V��;H펱[M�\[ذ%���s��7�N}����bv��P�vB�ʷeB�bw@f�G"O���� ��kۥ��RRO�P!߉�j�&��Y�����m�c�%�~�U�8xCƬ�dMrUؐA̡V�g��Y��x�:� M�q��u}و&$�\�j�l	����J�����:gɒL�m70�*9�����ۥYKA��_n\�<N��O�&H�L�7m�L��q	�W(`�~&CI���	K��`ryA`���L�Φ-��vd�Ņ�����wߵ;}�6�Sz�y��G�Z�(�v&���T�zbٰ��Eu�=�wgO���U��CP��I��Y�_�ɕR +$(t|m��1�>Ëm�Չ)~�7Q��z����-q�}3�#h�ՅiRt��!(Ud.#�Iy��i��M��س���֥!r8�(y��R��,�0t��s�K����s�<in���vw��M~�#x)
�(GK�l�#Pvw�p#������R�3B��M41{� �=��������:�ōh��N�ڽzSg� >�Yv#�����[�����}��8�����z8�����3�"�=ɤι��f�@˚��c�>*��p Sb���!���je<��S��G���QyJ]E��5@q��C�|�+��L5b�;jp�4�}	@��{Sp���b.�%�`~��k�?*���)l�؛s܄QA���v�A���4gCP#���A,� �M�&e���(�D�<�gC;�/�ݗe��'��;~@�r�۷����� w-�]�1J���U��p�������h�J�s�a����L�!�������;	}/k�Gо��Y�q�a�܈���@��kab*�KJsE_\f}�>XŻދěE��$m�T��'��;ߙK����^�3�d���׶�����fB2f��9�I�v����"�]X��h�t���v��s�������.��m�L�2�+I��/W+^�P?���SQ�����8�5Q!�J�_t�	�+
^�)����Ο���������;�'��?b/㰶Rb�n��_���Ğ3 ����^닀T�_u��$+�0߄���J> N������
�^'���Ex���_�`z���W�t�Z~-�#.-�:��?*s���l!�� �WPa��HK/l��&�S�7�A�~G2�z�>(�n�-p�ɪ����g)�$����ߝ����]�����[��x2�_QP��r��hb��&�*�h@��t�f��@�;v1�@l��0���� �	O�؏��u�D���I�A^�� �����<�s�rAD�<����w��hjŹ�Kʝkv����0d��6c�L��,{\��@�1@^.=� 3�ZPÖ&�Φહ�7�fѽH��۽R�"�ї6� Z?��� ���`��B��S5$����ŏ#"�e�kެ]�EF`%�q]��=�����@Hv�&w��7�Ơ�E��<��GTB@�/���00m.!a�vY�5�˓��C���#m����H������ �^q�E���?��_��H��2���[͟�F�N4��e��=N��$'��bh0������;Sz��ps3B��7t[$-IV��#��luP��eZo� �*�B���A�,�����<�:/FG�3S8�л[��	����@�&70�Ͳ�bp/)T6*��N���_.�'��L�ф�3��2���Ɏ� S�,�#�&��0	�!Q���vi�ca���bwi��e;�,ތ�0��r^�
 iq�Sl�׷O�yƭ��pZ/|�z��$�A�?h��\q���mu��;Y��IDX"���Ԟ�qs	����S!��Z6��7����n�.���X��m��ܩ�8����R�;4 .���xF�7�Y�j�ez�2) �T)��483>��Q�����J�̔��buG[����jA���8�נr�hϣx���e]`2�O��[J.ݛ�+Kd�_>�$@FH�:kk}�kK�qi$��d����b�6�M8~(��p��/��N\c��/jP�jRh��ۺP����-����H��KY%w�/(�>�iл�E�^h6��K���k �	��p�4������ײ��XT�bj�b�j����їo���]_�
�/��,�yGJ���Ir�D��*�i�o�Z��
;E(|v��x��塆}MZd:I6����(�s7��F�VxlL��3���g�1��N�����y��a�?�NaB��Y�����
�#��5[�1�4+ש���N�Q�+�]*}����=���jPm��s�Z��M2��9+�I&b��4YǸW���t��ɗ8�)�j� �Kn�t�x�pV���
x���x��4���������je̕-�#QFƊ���~HձF��k����o��J�>X�Я�
F�ٴa6�������~�ZOe�9E�vb�������X��Û|��N??�䛽(oEEr����e�Bt�g i�xm~sk�=��r���mS]���\�� ���:#1UG��6t������(�[�֝�����]�} �}���".��"�ɴ�<�BOC��H�O���0'(,4�S��$v����ö� �-�^{�\�k�ih���~"���Ь U�\�t�Q���0%`�d3m����/��۽ꡃ~:V��\\+VKj�(I�Ɏ`mW+EkxѾ�ƛ��s�$���1�w�B� �^�Xe�:�?U�&b��U_���~�yÃ�����u򓀍�6[��,�it0\V�2Ϗ��?9v:N�wn���R��ߐ�H$��Pm۠Y��rB뱲���]��8�\�/��������pD���N�5S��_�'%&��ܵK0z\�zxS��f�Y:W~�o:#�wC�1�M��v���nU\��?�9%�ٲ��Ҕ�;/D>�����	��9����8(�J���-d����|Y��6B�L�Y�Usz�#�������{jݼ��(g�b��
X�Ϸ&5�ϡWpf�_�=Zõj�R��Z{5�`Ě�.�[��krqi��N8�u/�7T�X��L��&I�2YJׅ��	�X�c��4{F��l��\gi�h��߷0e/�G�'O�M�⨜d�%����.��C96��|��%0>F�f����Aa��F�kw�^G&3�U� $�	_�(��O��ؤ����8#5�17�& ��Q�l��k歱�$�o�׍Q>:~~�E�9���@`�oRk�6���>2z���p�Q@�(j�,���I�|P-�p�ƀ�{/��h�/`�Z�j�<kdW�W��q����q��Sī�ï�Nq���ޏ0����b:���T6�{�7���t�A��:pc���I��gpևF��Z)�<�`\b�8w�KyO��q�@r�1������G�+��d0��`L��%��a�9�ڥw��=���GAӀa:�y\t����͡�p��&;���ԣ^g��f ���:q(���+؁2��i�?�Z!eO�b�yN�"�V����B�v��6�7�>�����V���
�?hô]z���,?�~���/�s�����Ǭ�݉�N���3r.�# \���c�#��px�!���s�-un! uq���3�_�EC4,�K�bH�#W�ں�tK�V��C�C'_o��Wˉ���&����6U���zH0q��<�2����:	(?�3�-����>R��]=�X�����{�M	�1��6����/[>���:�{�`G���w�\:���R�?Sa�f��B����2�Ax�񦁿%-y���HF�g�����D[�]$K�(-��-�Q�=]��
0��Ō�H�lF1�I�.���|��S�2��hcY��9��g�ݙ��?%ԣ�^�0<��p� Y�4���%�����QN��=��id'���[�� �e�jc!*�]r�_m���q�5!����\���gj�*[�c[/���#�Zf��R��5�ȍ7�Ia�M�����������2�Gu���ꏑ��sr o��|���xmK��*�Ohe��n0�Mb�|�x�Ռ���j����!��S���	���ȓ�Y�1p����9�[�������um�s9�6\��-��i#tF��&t�K��3Z���:r/�҆>��=l!�(�'�E�+ձ�G ��Ia��Yc[頧����w����G%�~�~%&���`����F�JC�i�I"���a=��m�_���(�&yt��r6��rvd����)qB1��@e�ꉡx�j1���c��X��G�sل
�ܱޛJt: e�b������{��M9��Y�ã���ۊR���0����x����r$��[�}��룍+nD�
�6�^�����:U��Nǥ39#��`j�z6oL.��hg���\�LGf3R���>NAL�-���O�s����	�]�;�<��p>&1��j&$�������y,9�R`E^n>\�`=d��x�j�c���*5��m���""b�� Ax��T�[0�s:���Ɲ�l��-D�R�~ x���{�.u�(p�u��䀥=�r��� a$ ����xqB �������q�+�hs��8����:`�u�T9̀�\���&X�6t�
���\_��B'p�㗦� 3«��n��F5�{=�xP.���@��J����V�`깔�2��d��ܯ+�ޢ��$( �2�7���:Կ���{� .��B�|���Jt}ѝ��-��� RZG276���aĦ��i��W�L5g��,19�M+e�^����ژ�zQ��haDU���D�Y��_�j跸L>� ,~@<�ldja���]�b�a�<�u�:�KF�l�:tZX��ͪe�H>����'��F�� ��Y^F����ݟ�5�c��b�-eG �����^ ./7V� ��.�+�}(.�b��ҩ��G�/�����aj^���~w�����Ps�
�."�}N�Ēcʦ_�$�b�%7)�2�P�P���5�X��z㾜��%!��:���ݔz�/�1��~:\�H��/
^	J�+����e(I������gQ�u�nݶ�|�Q�7~��G�lP������Ԓ��>�dPچ�1,�BB&-��"Xw�)e�;��۳�� ��� �1��!�A�lz��X4i�D����+�~��{U��t�@<�9@���dh����<�HC)|?�,*|1�i"=>I�W[k�N��7X�]�\뚛�3�]�����.}*y����+��LuP�+�v)M���0���Tv�ܧ[��H�0j�,8�}A��ye��[�l,�f���|�ڳa�l���B���l�衩N����%�ۧH>���^L����7������9�&
��Pp��_�+WF�сL��B��͸x��k.��ZI)(q�$�4�I�?�(��'���}I���0D�@���k��%Nk3XHg�qsN�n��=e:ł~+vU�)�TD{_l�Jy��t�~��E��rG�zr(��OY	+v�϶��Nz�y��3��s������%!>��H���{��u����0�"�	�*T���l�f�xڅ��Ms�˫��B"��S`�J�I7����Ϊ�����bE��t�� ���/���8�3=�ˑ3~�O�O�z�֛���5�A� �X�����j#���ta����E썖����gdb����nB�����kDH�T*I}/q1V���@A��~���lA�i͔���_@�Y����!�Fn�bP�C�x���βT�>йq�Pԅs^9kViYJ	�Zz��Ϊ�Q������E폀�,#��x������4�˰�~�e�`t���hj1?��1������6ӟ���.�˺H��&�ԓ_ 938?��G>��s���g	���놕�+���\�2UK�t�?�ngO�>�Du��y��(k�c:@��eq�ӎԣ���\|���ς�pB\PZK�BID��[�����_<�*x!=/CTl>���i�->M:]�U��	�5�-֛���B9H|��y/|}0x�sH�3�Ż=��{�7z�|��j�C�v������:�_��ԉ�P�*�k��H��$0�#�:�*��8��������}�^�x0Wޣi�RK�W$�J�}[�UEd�{l�,��dt���28�G����b�I�uH���X'L97�f>8�u��j�wYB&*4�\� �qԈ<N+y��(Oa,R�:���A���v/�����n�Y�keR�����#����}���/&ʅ!g�x�}<�C��G��9�a��+�t��V��q�@��x<���g��L�.c��=���;uqJ Q05.D{�j���G<�;�����mG�&�j|xݽ8ڋ��h/6<N[���?K�5 ��b�P��P��������R�܎��Td���zc�	XvA�ܠ���>�3:�8.Qr�C0�K���f*�&����p;�L�@`��0�C� �35�ؐw:g�I<�%��+��3�h *M��C?����	c֝��C�G'o�VQߑ�:�M?hOFTT�� v��e�r�_R�e�̇0��݉WV���+~}�rf�p�ܤO�}/ݽ���1O���V 0�(��!f��n���]f���cA�� ������FO�����/FA��O���
 G�9�i�;�8�'�Ɲ֘��m՚UF�ۍ.^,��	���k>_�Yd��|"x��ex�XQ
x�Ϡ��n.f		�|�o�� w���_������G����X��p���W�	Il�W���PR$L��Cǭ����o\<��q�*C�>>
{5+]a#43u���J4�!�d�J���I-/f����w[��v�����͓;$/ut��� ,�X3m�hH���W�biҸ�	��� �a�}5�ɸ������E���C�K��D�}4��C�-�5�*�{��Q��և��w^��ʾ��B~%��
a�v���$�� (@r�	8eS��a�#,y�P����`ꚙ1��# ����sWQ��y*5��n���X�@,-�4$�����Y]
�z�6#������f�i�Q~���赼�K�b0�)�L�	��2�ھ�=L($�w��D�?�'	����C�{��1��w)���e�:�`��VBN�+5�(�\����?��ڜh Q�!ɠ��i�hu�\WbM��N�gy��Z�~���=��H#]�8� 
�U�{��m ��^G�
��P��5��p��m`@Z�5J`�Q92�OG�V@�7���?�pt����Q?m\G�ʷ�)�pGv�?£�k}�������T�!+�x���]�#|=�f;i��N�,0�qo��t$�jF������f@���ȆDc-g�R����%�ɼ<�z8�*��sި�<W�E��Jto�����|�f/�A�/"�#�m[I��>�w0��P��8��Q���KQC{��,����{��������W��iy���-��h� ������U+�3�G��$�j����k��Iwm�<�rEfS�oQ�L�}�o�;���/+�1D	B�S�H��-[Ny�iSn��q��k���B0'��+K���t^���*E[�! �ĸkXR����%��`_��lv3G��՘h F* \����vB���6����+�ЦP�vZ����y�o�i Ϥ@s�H�� �;�w��_3�Ʋ�YF|'�)P��WAi� qD�̵g�����E�N&.�_-���[��:�;	�d&N�X�ލ�XC_��)�x�.�AU_�YM���EO���q����\��N�[��>�H���kw�%��?ۭO=���D����˼?�T&ή��Ry���#�%eB��6�Cu&+��+������!��K��i#m՟.{c~��G�7�I�V���M�mEyh��+����y��0-��iad��E�G���P�M���!UT>kh=V�g���N�Z�ܓ"�:��?PC��t���x �݋ơ,1��R���kn�V*�M�M�@�v��㣋 r��G���@O�5x��g����# �"9vE������&^���+�S1�h��%�\9\���Ѿ�C�|���t�u���6�>�*|�p2Fw� �����3�7�����n��~��07���k�z:���>H�_C'�"����Wp͏ȳ���P���5��i�5}�f�.��M��b����;x#=-�QP���ڊ�X��m���h����C2PN�&�j"�,f�S��-6I��<����2���8`cJ>��W������pw��c�K���c�(j��ZA��b��8r��OVX�ޠL^!�[�?|��ch9��'����Q|��oQR���7�%��{xR]]#�^�`���İE�S?�.�cS�>����?.V�ԇ�Vp:P/)X6����h�U���.c�f`sL&>�ctW��A��o�Q�zZ���^����&7��b�cV;����0d���� J����i��I��Нyv-	Y�j����x��,��SY-m?Eb3��&����� bl�S���fa��H������4t�6�gn��B/{��#Kz�X�(��r�mm��)�pBrW����*�j_���B��H�-pL�Q �J�'��e�������>k&��1[��S�lȑ��v�#�V�/,/Ŭ�?j��9��Ƽ�g3��_v�מ�a��1�72���B�l9��uA囗�1���R_;ܠ�� \a��"yZP��r���>I����a݃w��O�Q`=�,xR28�����G93��EF��4������P�'���MD�"�F5<��Z�vT"O�;<��d�T��"gC���b��(7�l�{�kg�6�T��~��e�����1G{
&��g�+R��We�u0l����D�Γ�_q��\#7�-�Ɩ�H�����DW��C���J�����$�����An�P	��$ּ��^���8�\�Rǅ��A�sg����C��<IOKA=��A�us췯=�r���4���n;0�Ȍ)�as�'�i[.�LD5^�4�"%�J�hd���-ǁ?�xR`o�?��I<�}��梼4�߮)*R�����z� ����/����C�vO�̔]�NؕWd�,�L�2�)7lK]$��f�w(5N�MV���$r^0�f#ն��YE
�L	[�I��!��V�� Bz�?��5�2� �e���I�̝B\Y��b�5|��u8�g� #@*�D�`�oL�:�T�]�5V�셝q���8U�k���m�q*�(kLS��$��+��_���̏�>Aޑ�+�و�'jVa��+ ���r"���4���%��:�FF��4�r�mb��i��R �P��"mP����G��-��1L��V�o�LX�Y3�>��5�Ѥm�Q/��C�M�w
0fu��h	�H��G�s�)U�H�)��k2y���跻o�>�	�ʫv&����e��7��#gx�"e�G��#lJVX$`����t��=?-�J!&�o���t�mԬ�j!�e>؃��n�/naF��
u�Y �_��n�$��+���.����a�M�c�
`/�W��K2 �L�*d�SX�NAY�'<�uj:y���YI�bT^��ߊ�D?���� 'R8�TqC�DH�p쳘aq�߼1�Da�7��\���A�8^R��K��i|��t��y�&*�>�ԐI�CfU vIg��^��Y�{��������Iu��	cˠ:<!�5�}���Y��B�������](qg5���!���aJ���p�cｫ�=*�9]'&�f�@?�.a<1�%���yw��|��u��cI,�7:�_J�jo����
r�/5�Z��2ZR��i4��+�5�� KV��}"(��RL�p����ޛ�'=TP�ifNw>ol_���Z�ΦY�����kp+��rN*�!�C5٣2�mí3�Kr��G���!kGW�=
�7��|n�|Q<�!,���$�؀o_�5�:o쥙�mfm3���{�7`��1��W~�X��% ���B�E�AH�9���a��Z�wI@�����d�VX��QaN�kcu���&B�N�
X�-U��gAB�$������\�zn�P�/E���=r�����&�Kɳ�����5w]J'��\�wc�,9��#>7j�&Ϻ�-lՔڑX�f\uՔ{�8�	V�#�3A^����s�`�RZ/H��^;���'};�r���b�:��z�h�T��K��z�������+C�����#�uxG}��z�����M�Hf8l�޳�K<��xv�$3f��t͝��؈��L�X*E�G�t�eEN"9�A�)��^k�s\�����CJC!�̙׫�$TrR�G�>��xjg7���!Z��:tYʸj�[T��Ӷ����N��Ù,3?^VO�``͖WW��a��C;�[�&0���1��YOU�:���x���&� P��8z3s	�i��r��L	R�G^	o,}�2�\��B��Z,3^o$� ��Eh]�%����O�+�����=�������AޛZ����h2+i�'(y��0��ԭ��J��V~J��Lh�)=/��N��?���T�B��d���W�dB���@���G��5��C����Mg�ߡ>TFC�H�⿗�{dφ짮���:�%�+�?E���{Q���_�ǆ2��X?���<�YK2�O��N���n�mNP��.��xy�<��S������kÆ	��YÿX]֚�[����i��JG�K�$ [0�`��y#	�0Q|�c��Q.r0��Ί/<�tgT�Z�f�8b��$�>ү���О����Q�b{i���A�HMo�Gf��l������]ʿ6�3ȵ)t�XC�F\@L/�5`�1�!��<|�� ��nv���"���U�#�<ʵ�b�]h���oJZCީfQ�^�!��tr��ΚCr�rȵ���K^�$�*��t�+��Q�.f"�{SI¹�N���J�ܪ�4;} O��O��`Eq8�J������QQ݅�lK*������P	}��������h9�s�1��+Xs�L�*���"����4��cI�)Oq�-��kC��,��������{w� $C5;�:<l������兄�Ay{6A�-j���#��G8M�6O���1���0
Hn}�ظ4����O�Tf�xFִ��`�z���-O�֔&ȁs��5!�F��]4��Tn�����u�]�,xnX�#��z��r��݅Non^��Fz�©��^�M�2k�;�T�Ȧ����S��'6���l� F�D���,�Ȑu���}�zg�4��ʩ��ն�lt�.�(�h���p��+��b;fl�A�[<U�P���ޓG�K��-����#�fZ�kp��{�;�5��d5z�)cF3��p�c�e���
�g27q@��1�*VK}���Mj�.�]zx6�W2��߻y�9�<j�ќ�����Ӭ�TF�i�Q��3�z� �w$��5� E�D
��>"&FF�����k"\��@�t<�凩�:����z���+z<�Wq�ZZS��@����k+|W���v��x=@6g������K�ʕ��2n�}�o�^0������}�^����K��S��O[�tb`9���N��"ϯR��v����?��a�>�?�z�jE#�61����PG���]
�!�R�C���0���{���S�	k>��,�����:Uu)��t@�+k��LGj��u_�����AM&ɻSP�U��t�T������0qȅ��܆]g=�z��n�X�P�"�d#2���0�Z�R9��N'0Ҍ?�W��;r���:���;�w�t���@M�Pm����)&4����P�g��m��6�� �a3U�/����$��+rͿ�5��?[�l��B����櫉�*�2�d���#
g��P���)z�Ѳ��r?d�+�@����$S�?�N�z��('=�-�~�S�@`'�$i��3-�VK:�G��g�c.��Z|�x�<,C��Zn�����v_���9���:�� ��ͭ�Y*���6L��y}D����l�hl���,�����Z~�/��7[V������#�ހԮ'���J^�b\�#��k�FQ*��ೱ�������IL<�L2ϑ�\�	�0w��LX]�����I��6kn��R�ɾ�q��pk�a֥^a��2��w��߃Q���x�HS�]C���{g�G�β���D4io����=GQ��7O��;y)}p;��Hf�M����C>�B�O�a{fLCY�
w3;���9;���֓^�	��d
C�2��;s�<�ݚ�돊�C8�c~�d��gF�6�'�.O)9<$u�]m�dQ2��{C�~�[3���^��$�P��~0H�ъC�Str����\��4�xYON{ٵ�Ŭ���T������	U��n���)!�L)�P�����
��� ��݁b�"��p�w�MS��2����x
E&ܒK&��c��[&�>ǀè�P-��Y���՝�[:��r�~V�h��AnM-x��&L̖[������ m��2�ǉH���%\��ue���'��_0�:M�F��XA���Ҷ�/�?Ƿ��U4�[��ʖ[��]�f*bb�_�-VY�����Ҷ�g8���yV��[z/��Q�@�`��{?��������zj�i3�#��3X�������x:�+�X���L�H�~`�&�N+
�3���_\�qٷs�a�Н����D��^�Ν��qz��7�7���EJ�9=I�i4`�"	�.a�+����*)�7X��Q9fK��T�<����$�����c�O�I��c���F���4�1����]�ѐoWpM��O�`��!ֻD_��{f��;��A�\�'$D�l�)5�f��gv��$��w�D���<����6��I�Ԙ��v�*_��~������	Y^U>��!�y�#��|�&�ذ��/������@V��v�&Dt��L�8��-.$�Es��H�>�m�Y��?�T�����Z�VTu#�7�"��;�ӂ��?��ً�*�G��Į�1��qhT.	_�A�<0+;�I��i�z8yO�f�1@���k��>VRʧ���I1|rk���(��ĶU^@�K"���0�/��M1M�Xu|�fD:�86t��&=��79KB����~W�X�����P����iOvN��5��W*���J�`�������=u	��ɻ�:�0�4�'-]��A�"Am%�_�OW��>�?8�cH�܀|��m��N�H�J�*L�DG�7L�U�%���8he�I� ���N�Ƈ�����C�nY���9�o`��pCv�#�g��!38�BϤ $h�u����+���<�α�	
�l�/��; �HOǋԇ�E���u\����[U��i[�]���ؼ3��+���:%Pz;�
�k�j��^�I�`Ԧ�#�8~2 �Lp\8�،�Sh�)��;ea�
?�f�r�� �_�m���nɡD��p��R�|U^�/}j.��P�g~��m��yA#�rИ`[gvY���e�-�9c��(�H.�Tuȷ�oJ@D���f�T�������Ä}q��O��d(b���$�:�{@�մ/��qٿ��[F]��J&�d�ِ捆ܛ-eZ���ѿ��]�ا%Ou����O��C�Bݳ��Z͊6s �Plh}a�B��E�b������i�dFE��)Y�5	���jm����K�9�{��;}��j�(fHr,%�������q�]�L���v�)��p%5~!�7w�CDqA���D�[=h��0qYDV�oB`�6[i���S� ��t�ʪ������ƥYp��ޓ��$�����)!�o�Ȣk�n̀װ9`%.⡘®��Bxp���V�v�0�tZ�#^m�{H���M���%b�i6S�jΝ���8;�(���zA�p^g`!v��m����<[���O +
�������wFr $���g�E�x����w���2�(��K���2�Ď|s9M��������
����4z�堇�^B�6��jP�������b�`9&x ��vmC*��W��6�[(\�����Śf�lt�D���z�U���r�����.�3�)���v�/I��Y���p/�/��]��=��#�r�f. ��}�4	�Q����r1xE�v�Id��]�:����$$X�|�?����7I�4���n���t��x)����Cōh(����~�UV�o�)NΊD��,KꩳT�@?��x�Խ���:������M~�r��X2SD1����w�����j!8y���9�Փl �y�A�_$^!����@Q�:6�
Z0x���ѼM���#��G�"u�/���>I�_�>���+qG�D�e��U�uX���SЭ1�s�k�*��ii����4V�	:��ji�8e߸��"�.�U;J�L�[���ŝIU���3���:<$�t�	�q�E~�ŏ�=z���F�ŵ��9W(����v���E�������%*�jt�%��xA��E�4HW���j���r/�7�R���_�h�p��'ѡ���9�3�%�:F0��O�*P��2�:�"��U����0���@ ��suz��)A�R���{�)��s�Hy��O��@��r�� �E��F}�y�vS������Zs�6�2yt���:�I�N�Ym���[�k��ZF��rr�������!��$c!!V��
-"�Ejf�zp���}�4�e���ج���k�/�J^��N�:!�}���������C�-u��B���C�7z{h_�憔�qܪ�Sm�R��!�]��<_@I�y��kՖO2��v<ԩL������Ę��"/_��݂���$R�uĘ�lZ���z� ax��(�a܂����m�{A�9����B4�p@��gC�-�G_>NE�I@ǒ�Hr�&s�7�-�<f��x6B ��s:�_�i��E�z�����'~{�I��?���6�k�xo��	~�L܈���Y,gn@3^�"� ��p�>�Y�z�%G������A�G�&�i����W�?h0��d^fWB�-f����rI�^����d�o�7�.C�<�2�_{�����\�gu 5rI�Ў�n�JNTk���YC�?
U�N��%��S���q����<���P�o�db%�w5K�o�s���9���'ք�A�_y�6Q�|gs�'�a�|�f�7�L��1�v��e������Q�Tr$�Y���K�Wq׊ء}L"�F/�B9������ץ�)4z���l&�2�Ui�
g���t��5�$2|ڃ��~R)��,,��Wެ직�lr!&r�����U�V�&�&,�u�}�l)�[��"!)
������=	I����Sq�y��.ӫ��q#yT4�K��g�{�81��EP��&���݊��G�Mcm2{��g[L�^=#eu�A�8/�Ў>k�S�����ؘXW�qo�����Z]�ƀ�8��批���s���B7�Y�
}+�^d
Dl���e�S<��k�k�N�M�\$���=��O��0�mwjdgA琀u��� ��V����+q&��C��_�L�V�;�wظOs��y���;�ꢧ�3j�|�~ei�����/~���t'����V�2c����e"ב�Ϻ%�g��/�[�ohP3�+���d�[�] {���o��%0ϼy?8�6F�:3�E[B-3�v���G��%��y�䱋�&�{�$a������,�h�6���-]N_�1@Ez~�?���5�C��AC��ސ��f��|�������x��<�<ۿ5�%b���a@$%,�ї�ĝd�K��S��"'��F>�������<� aWbo��U�����RE��>c���EH/U.�����-`Mӈo������������r��S�0���2�qP����5�.��^�#����j�ﱖv���J�.��ѱ�t��R$�����Y0c�N��˄�V�l�34�`_�hY�B��}p��l;���V�"]�������yw���gt�R�,�$��i��U�Ş�)^s�i5@����wv�N��}v�&E��I�����a�����������Aɧ�R�I�=N�$d?G���9�4~��)S�'��8��;�An��gz4�`�ڈ�_�����*ͮ����$�c,p�i�>9�ʭ$�a"q3��G�<�f�Ȩ/kwK��6=,h���u��a�pv�����0Iw	�{��M[%���󂡈�ˁ U���LY3����o��:F_So���^X�|w���{M�k��DAqh�q�}��uV��,�~�K�Gh��ܽ��G�K4r�R,���4i0B"M���E��+��_�-�ۛ��gx��p��$+jcI
����	�C��LQ"�u�h�R쌿S�W��'�d�(&�Da�L���3��]4@��M���\r�q	L͒&o☾x^���k���]��M�!Ze:&�Fk��5��eZUo��)HZ�0�E��PJ 'XVi�-v�t^V�s��	4"��GշD�KVX������Y�K�qw�65쐔��O�b{�&PHv�=������
l�� 'a�
h\�=�ō�]mJ488�m�t�����V���M�_��?�L��+T7@�`G�0(AزF$_[��ɲ�/?�9��*��t����)�\��"$��e-^�#vH$x�.�p�\�vw|&n�f`Xp����WO"��������������R�}�L�T��w;۵�z�㜔*���o:�8������{����Q]A�����v,�b�Z�ڄ��ܼ5˺��I,>����Lf|����3En���`�5�5GT���ݴf�c����)�1���/�V'\�p`�ͱ�i�g�3`oHƤ8��d��KO��
l~Z���2g	)�tNX1w���,`�6X��2��6�E�,a%���{E3w˽�`�ե�<
��͹b��c��G9�-�L@.u������O���?����6�d�����|XX�Gӯ �{�@��s�~���S�c���K6���2��1�M�%�h�!���E���1�����X����7P��}_/=�XB�p�Ўb-����ўر��y�Qə��۠�����<�<����B�p�߲/u#}ϡk���4�Yq���?ИN2�ţI',��~��إ�_nY9�+�A��覶���h�R�a{���&��������7�����3?�$�rn0�lc�~h�K~���SF�+��P�[�O�C~EՆ���7�ҲSF��o��$"g{i�!�v��u��#�C��Q�O�S�@����V��y#t�y�����W�X����x�}6r�w����G<dx��,��褲��i�����lb�î�z�>aHtZ,��Q���=���ئ_����.�E���X`�Mls�Qd@��&�����l����#��WX������>��Zٵ�QD/�ѵ�xEj��X���]��s^|'O��$mZ��x�h�0��+��5B��O8�'&PZH1%~�^?��ݵI��s�%1�!��`�C^x�?;.�"�O�b��5��I�=���m�
��xE!�#�,�����J�ο�ͼ��%#�c0I?,{���6�[Ҿ6��}��~)ܴ,P���Y4���鐺�y/>�����ы	t6O��s����q`ɸ�\�n�7A%� �9§JV��q�ss��G�񜭮�˕��/� �E��Bq��)��pޮF�����2�W�|C�v0 ~�����E��4:v�Lߊ��0�jTu�.��)ܑK�0J톌yΨ�\%n���)FpMY�,��H��EDl7��E�:t7���+N=�kȁmQ�J|q�?O9ӽ��:�C��w=gY蠞�>�$�⸕4�.����϶{�����}�O�vkpV���.W7	צĸ8_�p>0>q�wqqFos��|��I�Rl@y�w1����nfGW&��LF�*��V�M�ې5R�㙆�/7�rQ���Y$	`�'�P?#7�FO���К�b808���Cb(����{�y��h(T,XV���ft,�o���5���>���aO %�	*٭�-�s������];�j ��s��!��Y�0_��q�M�)��hY�i۫��}$n
�Zz����ՠTuH�+u�1���l�p�\�=[�78N-At��� c��3ī;�dod�H�N�-����YW��TL������zD�k	`����S��gFE��+�ϯRжAo\.�o�]J^c+R7���)������{R2��φ�u5쌯 ��ڷ8{ٕXN��*p�5���U0���-g���E��������81\�NCt�#��������9g��#�#p��%;f���n��Ë��S��P����V,3=�v?ke3��E�l	c�bWo��HT�A�����a7QA�n��<��˶�>�pu��0dvLl$L��H��A���	 b�\|����� �V	�RȄ���30��@?E�nj2}$(�I��PaE�z|���UC	%�Y��ݴnA�&Y�aZK��p�-��&��I��mLO>-��m,J �@��3����ꧭe�CZ��jm��؀Z����d���� �����9�D&j��lAg%S٧����c�|ո�i
��-�h��`� u����i���U$i�&�D��p���쳛m���J���,�K� [�h�1n���t�4��/i#�9��D�2�By;�G�����%_*��N�S^=�<ysL��It��v%<k��'D���0��rbL�W_��v��xĮ\&��FBG��&cO�h�1�4�4\�o'��g2��V��|,V"��r��C��.9�K��|���
�Q5�H�;���
M��đv'��љ�C����)�==�pH'�^S����ؘ#���������ۥ��(�����}��GrYSX�k�֍�����ah��Bi��3���=�*�G�gyYe���m;������m��|��q���y$�w^!+s��j/����K�EI~W��X�L�3B�vD�a���|�d�u���3�C��8�6T��K�Ј�� U4�?~w-�!���	�`*�C�"[��� ��y.�x+�����f��^�n�Э?t`�9� x���:�i7E��������f#$�-Y�����pST��Ӌ>�_�V��q��_Љ�و�'<߁���o�����
����L�Yo^P���l���"-�R^�$XL�a7�XCP3�Jŏ��z{�W��uǒ{�Ĥ%����<�/_�ؐ�w�i��G󰺌W�g�V	�	�t������KȦp8�U�\������T뜽Y�Neޮ���+��9��
[�y@|In"K�J,UQK(F�\����h!����R^N}�a�"���hj�F| �`��RO�ooX=E�J[`R�Wǘ��E6S�ΚPԄ�q-���:�)*}�N$;�~kς��|XCN�-���h�;�������ZXK ���������5�n|(�w5���7U�]v$��9�Ԟ։�6����5�'g��2�oA:�߶�������䓝m�ّ7�	��4N�����3��������%+�o�9�
�[��C�2��*4�SB.%���ɘX��!5�����:(6��V���h?ۮ\@� ��������:=-!�n�&���@U���v~�T<��8|�\IF����mO�I�xMڠ.��q�1S�.;UA���*;���?N|��;�����ڻ���]m�ĺJ.)ZA��6�J�ɀ��}��,��8���Bk\�3$�D1����ִ��u�ː��9���@�Q��
�x�A�Bg�{[��F�B]r�t�����aq
?H�G����vՕ#
�j��Z��İGr�x9 �V"�N�4���l6�@,�愁��W������wrhi��Y�M�*:��`a�_�E^ll��y<q>p:v�����;��5,����\f�!��Ւ�j�91S؍Dп�j�𨮏����09��:_�P���������s�)�P2I��k<:�wu�W�y����Ԏ�p��'��o��A�Ĳe���p���;b�p��p�(��w:� h��# ��t����ENxH��;�$G��c3%��o��G���Df��,�צ���?t�1n��a�w�a��D�慔��Tql
(5(^+B�<ͣgT��W,��$���2��"����ZR_��B���pߗ+H/�Y�E��S�r�+"�6�L;P��Z�Ǭ��ú�n�� �d3�&Rj8��~���j�LiC����W8�D����?&_�/�"A����� �CZ�}���)tː�yW�� �G�G��j�9��-�a�W�ؽ��Ӎ2��Cc�� �v�?lj��ȀO��)~�A�;�;�	��,N��U�����ϑY��3dD�p��P����-�D�n��M63]G���uv�.��G���H�bY�0�T��*]���p!�[��^N+l�a�(�F \��QL�▜U���|b#X�z,�F[�dg��˕%�=����;)��y�&%���1����:�Wq�V�e��oj5��h��7F��U��:/�ٚ�X��쩿̭ˇ��u>��U���#�B"%�n�cq�y�w�+6�6��Jw�d�0.��w�����˖�2���'�Zݺ��/���{y���Z'M8�E���Ld>C��Cw�-͏-�v���=~���j�6ɳ6��4��?�qۮ`~�ztK�n�@4 ? �2V���RJ���%��]z�	�KbF�y��Mw�;��e�Qt����\%Yx�%+���9+��ޯ1��h�qY�R_��ґ!�%+��9��B�t@7F?��/[��K��㐚�y�Y���P;�ܢ������l�б���n�f.r���%�����QJ�I�3O"�����J<?K[�����wn���f*��gF��e��
^`������"���3�T�L�G5��[@����������C.ׅĴ �~X���㗫i|�������d�k����S���h��q���Y ���4��`1IUd�S�?��Uc�.9V�H�i�t;�u��[0�h> 0*]s��n*k��)X�����=Uٯ��8�&����ʁ>�k������kkr	��9Y��,�������υ�����$��b+�	�I��Du�y�`N.q��Mo(C���<�p%��?|�!�5�bJ�NI�UT�xg/�䠅��1-�7���Ŷ�#�]��
Wr��jв�p']n$��3�y7�k�D���)��6���H�1���6� �!yZ����Y�+|j��
�y�V��˃^6d���QhOj�閥��o���S�݁��7SL��r����e}�x�ڭV�l'�F��k����']��R#���)�hj2%�4�W���&���J��3�3�4jaa�$Ƙ���Z���D�l���u-��ד�i���Df_���������t�R4��h �+�#������2�F
���hM�>kV<���G��O����X��$��a2�����$�8Qܗ�X��F��Π�m�������L�5]�,�>0݉��\�ho���l���m�,���)�Ӿ��B�<[da�%��("��Ϊ���9�������M�g[ϲ�P�>o����2����cz��|W��b�u6����>�6T�QE�>ך~��}��St�5y����}����>�<�eg݂�{��(�rК-q=`����0��I,-�)�T0�cڒ�x���#n�@p�{,�w��&>i�'L�*�e��W��f�y�"�Z[u����}��+pkz:��)j����`��;ĝ��W���>Oq��M�Pc��V&������^����X�*㚐�n�ّ]����r���t\�G�/@k��� �$���3"�g=��.;ň�*��c������I�6<�Iǥ}�G$���,Zm���;]4S#�[%Jߥ7_�c��77Ƅ��[��;�����(� �2�O"��Tu.F!&��h	��O�Q�v���f\%��s^�˖�{>�6������u�D-�ђ�:��KO�]e���#!xR5Y�XYi�t���\��|H�P@��r�8�R���6�:��g���{1�bk6x�B4��N"��Z	�YN��-�tںȄ�����@,�b��nL�R,��"f��<���Q��X���Z��^{�M��� �)&�x����0;s��(<~:�6��=�8Xyo�l)�{Q�\�=k��C��@�h�1���h�PΏ��F&������k��Fc��s|A����{��M)|5��sخ���8� 9��[�X���M>�
銰[�Sۨ�l����� ��F*6RMw�a]Kh�,#��2١���D��o��bm��5~걩�L��wyflG��]."D���b�r�A�Tn5��i:�Q��Ktĸ�'
�ꃛ=o�}3W
!�[�It"�sL���c�&�L�Lq���̠Q\𐜒� j���o��_�2sQ�z�%������*��%zh�r���?V��SaY���88k�Q.W7K��]��J��r��י��H� ������Hu:X@�����]}�vm̙]���ǀ�Q#=����І�V��\�����z=	h �x2c���BN�1��Cv:Z��i�u�����Y�A�]5�ZyT���(?ixo��ͦ�X^�5&�A�4�;pw�15t`o�;B���U��(�������`*b�u��h땲���R��N�o��ܹ6�YE/�Ǐ�W�O�DPF�]QI�=����"mпq�אE�#��}Cj��6݇Jff�q��O�> ����7^�0��}�zo~0М�ό���оȸ%��=1,� k��m���~�[�h<��,b)]~���Mv�ujGw�:�x۹q1�����ƛ]���j��/ݘ�FN�f��_v6WM �f)7$��S&��aq):�W�ϕ<�P��f�[�S3$���x�)G���yr�sq����8�e:�_)�6+r�$-,*=���R:+9笤�W�rQ�Q�����Aa�i%���N6�3�M|���gb�[$r�?0�o�W��,��穑������+�gHʞ��Bbg�a 5��}�$o�n-O`�S+�8�ʤ*KVW��l�"��������N%�k9�� �pk�v?���QzՓ���H53AYś�X�3j���������O���m0����0'�[��VAu�<��t�ŷ���w��B��ͪ*��;!�M�ZX#�Tk#eA�$�u�w'�Am?$�[v ��x�����F#@��]������|м��9�\+���5�ug9M�EmO��w�yC��5ε�s��{)C�Z0���iܗ���_�j�ף`�_ʚ�A�b��m7_Hcsf6��͝\Pq�ښ��3�lM
"p�ý��o�r$ϴ$��Q�Q�;�[���+�2Yzzn���^�d�Gn�=}koB�R�q�`8��J��:P��}bz߹�����w3�iИ��`k�Ko��v��O����p�y����ۮF�z�.�-�L����׫~#�!��Ū���?�<�̀:"��iw����u��N��쟤[]�_H����šs
��~+V��PM\�TIn�A�^�l��XW�K�E7bo��"]���]����̃�Ȁ6PU��G���oO������D��OI.ژ���A�dD�w;��6n� ���}�*����
6s5	7��4�1ϴ�F�g�1�V��"��b-_����0�k7�g#g}����3��鉫��8�\��-�?�;R�X������K&,�E� ���0<X"�K�ȫ2�};/*N��M��h-�o�m̬^뗟�}�v�� ���&�v�i��I���v�l�W��v#n`H���o��1C��/���(Q�lt�۬V�3�jZ����X&J2W^�D�N��x�<��G�w�x��i1�5c���4��5��gs,׈�5�CS�K���
�]��é}`�l�u�;��X�=�򠊢B1׀�"�.5	�yR.��ι=��(����~Ѵ
X+�=\K>�|-�V'�*kSP�0[�p�'.x�PN�_z���'�6uVf��4��X'��r�/l���R��ù�eG��XR=x8~��2�J�`ݖ�򱶞�56����IH/���G�_��#��;��JzP��
+#����4��q�vא2*?Vu԰�I�8�e/��pI��U��9�u	�Q� gC�Q�G�1m���X�V>�S�����`Z]����GD�eIv�D��K�$�ҷ���V4��޳'�#ʜ�0R�.�Q>�Љ���V]6SN]��Չ�
�$�SI~r��?��(��"�=+	x��s�[�5
_��%1t��ZL������7���SB�"����D3F-�$�-�U�4�/�[��vq�0jي����Z�,�P��^,=�ri���mtV�liN�pؑ{���X1��>�TE�?]�k������ 5�s�hܔ�w���@YC0��H� �Z���S�ֈh�
AO\@q��Ƚ5�v�������aRÈ�U�;���Ư�㠚&0�e�:�N9pi�{נ�?7~�g@�H�]c�wIu�10i�����E�Y�����"�G�\5uTEp�R�$Z �d]���޹E�����Z9ב���)G�1���A#"���K�#��P�+cҚ��F�&�t�j2��H'��qI��+��%�)�1��yJK�-	��ɛ����8;�[5=O �z8_��%�M��6�sF���b�+O��.n�'1D�F��pm��F�����I��K{X��� ٸ�<é�Ϛ�`�j	����5ZM�	�.�e
D~Ĵ<�Ȭ	��Ǜ�K����Y_n�K�)�sjNў��V��Z�}/P���+�tR�<uQ�m�t֪�?T6��O��s>���_Be����y�_��m.����ɆKBzc%�2'�X>��
<�2\�s��$�Y�T8��
�\zZ��Nm�߹~"|�^z8�&�%=�6�>e�����~~<�.���Qπ�r��׶����VɌ��S�1{��c�,�n (z�e��8:�3��D�ǡ�}�h�����`�
?�T��zSP���¶N�'7��9&E"i������J%��T`��rK^oK����B�����:=.���z�S	W��L���5w\M��FW�윝�.R߶ӽ�$��Jw}b�gT^�&Β��Zr;��ɢ�+����ۣp��A�B�d�*�k�����h��:'��A��y
xT*0�v��}h\p6�y�T*��C=�~z���8?,�M�D���mqc��0�˽�۶닧a),LH�!홝�έeD3�0����'�*i�h��?��	|���',�o��Xf�� ��8�
1�o�a�-
U��f�@��l��f�|�	k�d��r,_Uћ&d�c��ܾ�E�A�/>���,L��6"��nMY�c'�&�H��8d��h,�L-)5}2��j��	�)o��.t �"��֗��_Y1-�*���#T6�~��St�p'�	?>�s�s���B�_�O!�Cڟ��Y���Z�q��a6A��xy�v*��jw86@Ab歇7S[����^�ڥZ��*l���c1�9;WQO6G.������֢`��G�V��S��D�����6qd�<^ j��/�6�96��+�I���3i�����n�����E
|���X��'Wc�Ju��e&�rA$����n/�&ܯ#�:|��Y�i��Ȝ/��ﻅ��B`_A0X�Be���]|ɵ�+�[��%Bc�U������������ނ�G�]zH�����W�]=,�ʱtYҲ���짲I�\P�JѸ�K� �&Y�[���j�\�'�
��/�/���k����(�����v\O������GѲ��B��ͨ�e�Bˡ[F�t�)�9�i��h�����(q4�F��\�V�*F쪀Dа�iy�Z�B�O�b�OJڵ.i�����8%��T���1q���4ޔ�'�g\_�ZV��,������e�E2�.T*>hɃ{D����i��'x�Em��z��k�os�J�:�J���{xp]���M^�خ��Q Й�����R��V�CB`�!�P����*s��V���������3��������Z�6�._�)+�p�4܍Zr�^֍�l+�V:���M[�ҍ5���RT�y�H���Ɲ�Fj�';2/>}Ӣ�cC��>��Q���Y���� �gӣ��X�(I`6�t��)�C����;�E�=C\���{�as�)XKYܕ���F�_5������)�
��H;ԉ�<�[��n�m�y��.�QdGb)e��@�q�D�f����|m�^.@�!��=����k��b2�{���m������
�s�2T�q#����7�
A�P�����B�YŤ���&��j�߬�\`���ը���ZS}!L��H(��	�`�5�}�c�㳗h73!��ٹl+r%2[M ��ף7��0��!�T.5\���[�#:��yR�装�Sk$��д��d�k�=d(e�Ox�s�`sȽ��d�j�]n��k��* �s���rѧX�	>�m���W�=��1�����v�褀�K�A$+	��ο$��S�!����R
6(�~�V�"��8�z�	��g��_�� e��T!��5�f�V�z�J��XU���\ͪ
Db��y8s�P	q���
Ν�eHt7;�V���F� r�\�T:u2��r`�bή�3���M^��)��p:�^��҇��z��~�;��8�>F�?y��娓V��b�j�`T�+_7���H.8��̦+����ي;�&,�'�Z���{�?U�xf�%ÂĨ��/���-̣��9(�i͒#}��Lc�& �"�VC�{���ɼ���uբ �^��[��~�7M�"�7\�3(��p�� � ~�-�_��7�{���b����k}JԲ-7�Gk1���dZ��X���4�]y��L{�"��WE'�˒��P)a����h��\����]n�n�fw�[��U�Ӈ���1U̢��s�9��V�5A[��y�F,��켔ɦ��3���<R�l�usߠ�:E-H�����]|��"J�Q�ȑ���n;D|N�t\Ce-��VmQ�����,���b��oa8��$3�$V�7��p���Cor�Q�(lS��3�i3~l��f��d�.���v%�9����
�F;�~Қ��	ǁ�� ��*��IJ=��/�WQ,D��~LF2��7��2*��5�ؓ��Ⱥ���Vb�3vFi
�$�r?�F�|Q����K̻������#`��Р�yΒK򌁇9�@����f���wG'�����o�x��}VjkR��$m��_w��,6ף=�;_�t�C�[�x�T1Z����ƭa��_�5*�(���
�3�6�ҏ�͖���Y�y�)Rp�����ļ����Y"�$R`�(v�&(��
m.�L7L�3��Qt�0;��8�uħ����h�O�|	&�H�IB�9�}EriV��K*]�-�!/%{*0K;�qr�ywi5�Џ��PV�:�1V�`�;��n�c�ҥ����
.?�)q�~�QQ���8�5CJ��ĥ�4�P��Xy�NQ�V��B����4B��a�y34g"����K�Ӽ���#�U�oĕ�����r�����( �0���+�r��k�:���o��:�;"��j7�#�r�Gf� .G�它�Q����Nj�m�VIgFg>��]q��D1�����p��d�Z��Q;�a�{�B����0���HM�׺�:T��]99��DwF�ugT>9��t�nъ���#B=pVO���lU��u��o%�|gH����1���\w.�F���
�(�z���si54���"��a�J(��y ��:c�T+��o�����)�C�_����j�n٣�O�s��!z������Ic�)&D�Y���_���6[�4m)>Ж�����^4�k��l�		0s��;-��ފ���;�CK#����S"�r|���Uv�8聣����� ��-qi�^�ʦ��#�QEQ�#a6��Vأ@�v�����ZG�M'�I_)�O9���%�l�=y]PI{�WO��V�J�٘��t�#o� �=^h��0�|����
��C��]@�3/����z	�	�ՎW\W7S��|ļt\�^m*~���3���T@ `��(#	)�Ϛ�ˎA��Y�y?�OϺ���3�R���f�UO7#���"T���^�Rti������E�A!����8�ZJ'��T ��� �RP?�/��c�LҜ�_�=@�N����,J��$�nym{^LG	��;h�ֳ̥�#��HT��V�]�Y�Ov�4E�I)�r��3��������lQ���;P���tg��Z�
GJ��Ch0=����C��4/}�GA���Sd��t7����}W:Ӥ���� s-����-�
�.uC����l1]K�Js���t��c�#^���t�����|1j	����o�Q�n������$�����Тc���0z:�;��	N$FN�����Mw"��4�4�B6�p�(7�t�/q���
}� 1��5=t�6��6�\`��0�������1�ȓ����?WQpBSh��Bi�3���J�h�腮��׼mv a������l����:�$F&7�Ƀߚ�H!���������~?Lo7B�ɭ?�S�i�h�����RZ�"f�	��w�PD�?�[pw����s�I,I�������!�؞�I���e�8�&v��_uK���0+'mn���cM��a�"��H����9�բL�E��
3r�7Ӆ����8�msD~}z񇩘6�ri^�G�^VE��j�}s��l��a�
��5�A�˵��P��N�Wl%���F%���q��5�Fp� �&����Ef�e:Fl"Z�?J��hi��Sҥ?R�}�!Z6�P��q9��Z���"�e��F�D��j��ǲ��"��YG�Ĝ˨����-d�B;�S�8)��4���c�KqE�Wf.�Y⧳@஦q	�D*��v
8�A����)�K)6���LkZ��3 ����=�K��1ׅL���*tI�ꐬ]��4 t�R���M����à���+xfƾ�o`:X���'Z� ���z��g�ޓ>�ʵTI�Q����Bb+�|F�)��pHr5�(Fnny׎�x��z���ݣ�e�����,����~�G�U�c����|-����ɦ!�c�A�"k'OW#�ޚ	�%菂'�	,x/��dd���J�N�`����ʸ*Sտd�J0�R�8]jRΥ�uJ�u㐳����ڷ�Oڽ����:CP�٫*�����5b�6�R:�~`�v����oA~y��h�[�O���\J �#R�PQ���q���(�%uoCGխ�	8��,����_�q1V��U�V��<�h�oO�l��A$�>�p`�欖j�3��Qw�(�ڰ�@�A�w�/�G]=�7��-���  ����Jn�s!2Ys�'�$I�&�^�b"s�3A7Į���T`"H�"��1uy�Z��P/I�v!JQSc�{N]��;�Tݏ2��Os��j^f��w�}ž�C���(�#�6KKj�V���im���I�QK���k�(����i� "��D�Vs%0���+�S`(���'PF�m)����uS\V��N�i���#�爓��%]��}rU�`C(
%��%�iڑ�6ϼ�DQ��q��F����{9]i��^L�]Xߙ?�GF��bI��V��7ۃ�z�f��b�NLG���$��q�R�F䏗��Tךٰ;�0_^����SIK-f R�)�/�cT+����Pu�dL�-�=�����ɬ�[��AƸ�*z�K7�c(D,�V߅�+,��j���Pm?H^�fK�JD�S�7,�i�|"qu�1Jfx�ŷB�<Um�1�����%�^�'VH7 R�K�y�2cc���5��]wC���/�kJ�S��Z����Ty�;	�o
�#���x}�J'
�p�ZSa��.Ox������s5�n����z��km8�(��:�)�p�}.Yso��:h�w��{�D����B�n��2���cB[[E�4�d��*8�D��K	h����lcR.o�tk�د�E���IT|�V�u�j�eH��/�.r*p�5�HOL��;���Z�k�~H;{~�:^���KD��ؙ�B��D%$��T����91�&��7����hFI��"`���mŌ*�R��q��O����p˦�6�f�}�v7E�/]'�"��PJ���Ulc��*��.Q�;�*�={���m��c<�=-�@����g	1tdt^� ǑD�!��X���`=�_�"=H�B���L��m[�����S�'��m�E�����eg�PW+�2�\���c�
2�Nڏcʨ�a}6)k� >f�I#?��g���������v�~�V�5��R�,p�1s�`"�L%�	�������z�-�39�����^���gi��C��H,����?�>?7�8�V`h)�^	� �O�A�ɚ��ի �d���6и�ޡ�T0��%̯������)4?'@8c�A?鿑��tlLǁ�o�^���b稌��J���Na�	�,y����egE�S�4ĜTR��V2���O�CڔDɒy9�0MD1[�~E湧�a~�Ys��.O�⼴{!o� xśz��\f}K9F��S�+��?�-_)��;��[�"�@˻�@�L|������^
���Rn�ֲ�s���L:ޢl䭇>6j�xΩ��r�x��Bz�/Vl�d�I���7�����NM�V>��џx5�#��8��<���-�9���������A�[_���u�^�D��fOO�6�)=���Gc*i#f�G�5�}�����^B/��.�f0E�C�&];d*.66�r*J�S4��P�՚�o�$�zG�aR7�u��
�}t���N����gG����xk❨y�uL�i���hHb�"�T砜�=8����*P�mau���:Cx��`��8������n�3�e�432����J��� ۣ��ү��w��~8]����-�$%��O�����8[��)��a4��]%��M���Z�q��!u���/8$1�Rdһ�^�����4��X��G�7���H�@�$�n*=#F����9Vap�!�Js��ǵ�Y�ߩ�q 7/��O*��x�F# ���ʽ�$E�$��n�!���R#dPp&8~��V��3	һ��"0�r
rѷ�����Z�y!p���h�'�"�2=d�1/mȈ,�b�{w�%n��2DTobp�r�ˡR �Ż��¿��:k���������z�8*�:g�O������m��5T)���L�f�[F��ƕ�]�_������rKJ���DF��@��q-�x[�(�����o�%M�3E�"��SpJ�`X\���S���w��3�豢m��k�vh��H��	������W�F亁ͶR�K�?a/��J?CbWM��|��.ύ��=�kz��?�_�PK����Z.�h�;�����|�f.���1����}�@@*�Ay�~A��s���غ#���5Y0.�v��A�%��6F��5��fV�)Bۧ��]�G��G6��?!	����+��Uj[�_P.�����M�0�	'���U��q�6����=����x���
��e��9E�������]	�{��n���K6͵k�Ě4����`�m����h�k���1�/�=ӊ��J��g5�r]g��h��2�$��ע�� ~R������tǞ��>�!�l��
��z��k�F�K�f5��YL���8��aU֤6�>Wm�O�ǜ�-uGQ�>-,��#��,�#uB�!�q��X�EX{o9��d�plܹ�QN�"K�I7�P �[f�lȱNs^f7ϵE%	��蘻�q���$ ?��V�R0��у4k��=E�$}z)l�i�a'k�)N��ϗ��s�V^�����l�Fݭ�rUw�Pډ1�TH��,�y�M��	����f
����n8	�9�
�-�H �ڱt7��XЋ/>��q��, �=T�z��.y��9�^:��Tz_�qN��Le��ЄP����D�]ع�۱�|���Z��`VA��uiڌ	E?E�S]�����h�C��ĆL�9�����tUjp5�<Q���x���Q���	lV�p���^��$��<j�؎{�cE3]Z���s�����Z�H9$��41{��>�2)�`Đ��9�3tSQ��� ���(8����_��u��ZqIkM/��$�K������᥆����qW�'E�����[��V,; �~q���H��m<��?�CɃ(i����Ҝp��z�$��ĕ\�j�J�
�A�Jv��Z��B�d� �_eRe�t�{d*�t&�V�2ăAHr'��{,sU��+ݖ�b�Sx�<9�C��-ŝetz�%3b\��z��Jv�q���E�t�䅠N�{�h�g�o2�k?�����2���J$�.�Xɢ ,���=&�R��y�"�`����±߾ʟ��R�B#T�N}[��	~��A)]�e(�Iu�;��J�kA�q�h�oѯ���t^GZTꔏM��olZ�����ME����uH5����ȏwp�U꽡��H�qs�}�!|4 $҄�j{��K7��{Q��.�Xit��& �4@U��uK�(���i���.x+�1B�'���:���iQ�W<}��R�j� x:�C q�R/�i0�R�*k��M�&H�s����D�T4A��Ʈ�)j\�Z@�q��<�J_�xￒ}lҌХ?Z�s6�4�R����?mh��M3a��+L^�֟޵�'�-�3�Ss W��2��md��P�Bl͇M�V�v�J_�g�Y��I\8��y��E����\�#�~�r�?|��\��ޜ� r��G�+Ѧ���v�G��m,��1�z�2�~
-���ByИ�QJ�Z�#�s(�$c�|Z���'R�}9����u[��5(*0�i�|�
�P�dB���o	Z�O�&.|<R���P���_����M3�m+f!�1�Q������Z.�ۛZ���V��T�
������K�����������?a;��Kkv�
�x�֑�N7��ai��O8]Q�����#��b��*|�O�c/��4�#��i�v�����Ȯ�AV1�ݓ�\��8 �Z�Z����H�v��d:ʼ=p��pPD����	5�"�H�q��a��d��O~ZJ�!��J4pK�>�<�a$O���8 2�S����}ċ�֨���v�ey`g�n�S{�:�Q��jw�Cv�J�x7c;W-Ӽ��Ԓ�Ds����OO4�e��``��(�S�o���5!�>��B��s1n�n�ɕ�FN͵�I�{�:O�Ň�0��u?Qr���u}u�y�_Qx�t�z���yT�u��P$��n��3.�b�c��I���a 8ꛬ��2�7��d�A�BOVQ�C�6�U?␲ߥ��3�S�+	��!�pH��P	�	D�~L���A�F���o2]X�$��-l��ѤO��*���1���i,��n�RU�N�$���1�U��L�t'P�; ���N8=���A��2=7�o�&�8��f�u��0�Ko���mFx�n50�!���b���B�)1\
U�M�VKDB�vȀV�A�l-��G��)�=yK�+��Vp�RǍK��nݎ菌�pYɅ;ج&M�!����_@�aam�9�R���k�1`'^��]t!��n$>?
O��)���ͻ���2�7�ɯ^2�;�(�� i-i��_`d��0���T.�Gf�Ob/A������=�پa9;�e�Mp+���0�K�+��C~UQA����'̜�f�Ќ�׏7��n�����@����M+���߁=b��Ri'8��q%A���0#]|��� _�Ac,�Y�4c9���m)��3%�"Gy��M�0����Q�����<��O�zτ�����9�'�{h���L���~UN�ݴ�jyNڔR�F�"��_ٿ�E�BkD�U;�n��i�m}�*Z;}�@�kĲ�6_�G}f�@n�pv��_$9�7��M��X`uɨLh�l��qͶ�¼�й�i8܋*q�������_��:��&�*~���P�uG�y��LƲ;�@���嚄�����0E��/`�E�9|� �������4��P<�����X �T��I��aνG������	F�Eo��7#g�7ۢ�/��~7����c��A�N���zTW-�W��m��Z��<�^��F�����
7&�T�ԁ�;g�:�]�;IT�@��rR�py?3"��t��<�I�=�d���ެ}=�U�k��n�n�8�b(-fIi�'V��/����/aː&��Q���!���y���YϿ��V��@.��>��~y�wC"rI��j���B, �{o�AA�ɪ��>aF�9�������5�"�R��:�-ڱ��l�[b)�_3�2WW��R����lP ��K�:���rK)�˼�t3���sv�4�8p�W�M�u.&�Ot����p�ň:�L"c�"�Lh �m'WJ����0�}�P�Tv��D?�8�1񂌬�t�V�[ڨ�T$oy�GP�<��ߊ��b`??�[�R���\P��LUk�[��$l��i�)�&eoB�An?�#r����}�)�p��d�5Ij}u���l1QD���f�k�}n~=�_#{n|Х��׾����F�ef��A�d�=�u�o���V^���у�`�F�4���_�A���Z�$�殝�I�5W-�P��T
`o��,�ȫ�fs��� ����+Z~>C�|C��G/[� ?���Y�<S�|��ț�L��;r_�_��F�/. ���Q>H��(g�E.AKl�N��Q�|�@�-�[��uAo�Ǽj��Ʉ�f&�6����쒷��$l�����*��'@Q �~c�\^�)��`6�k���S��@1-!H���E=gk!`�(�h<2)��#�3���2��1���,���L!��_�����Jq'��vs		�(�t�1�^�J�����.l�*g"����*$Lq,��aFC��㪕���2GF)�k|��t �~������0�`h��Z�H��B)7Z?�64sJ�o����WX��p�=0�Rt�U�nn�}��rP;uoz�/6:����E���-UGu���+X8�!��9���#CufhX�)��}�Q�퀣���<o�.QQƃ��$��yME�s{u��K���/�4:���MvTYc�iA钎exP}"�&�|v�Q���?
��r�l�Ҩ���jv�V>�ĝ�#�����x���'{sY|pR8A����:S=�J�\G���-s�2��2��=���>�'Of��Ӭ:KkꫡA��y�Zn�F���+"Fu�(�+�~ۦY��oN�D�0�.�yw���Aq�]Q1�@^�_�O!6�B��*�ٟ��c�/�Ɉxnz ;�t7��\A>:]\}�*��k�S��������O,Pϙ����0��2��2�P?��e������8��m�(��Ϋ/{	�)�fq��)�����/8y�g�p��OS���a9�)�����$j��4q��'��e����,�n����`6����նW�=���������ñ����Z嚺��.f@�+�=��N@`c[�"�y@Y6�66U��.�"Ѹ5�0�¸�K�V2�)��c�8�r�T��c���$�B�*Y+�6��,�cڌ��������1��D�S�l֤$Ɂ�eT!������ ì:�cR��iJ�t29¬�M]�.����)Cr%���~xã�X�I���=N����Vzـ�~��;�����6Fjm�6C|	�����<xg#ُ�
������z�H���ڭ�B܏W��:����K�K��Gǣ�e��L�s�@���(�Ghz������e+�$"����)��U�8/����m|/<֜5��ϮaL}��=�@�����pz�����q�0�}���y`'W�]��q��?DQ_�v�#7�˟�u��!a�� �80�'bS�*S�����ղ�x�=�yN��~�q7j��Up�OH,.�2�&f�,n�G��ԧ&5A<V�Sh�B׀7�M�@ѮcnR�u"��f?�����k�����S���(Νܑ�J�KN@�H%ȥ�G���⁝���J>l�����y�)���nt��X(�8@H�@�1pk�C'�����m��h���J3�� ������>���x��g�.���������lH���eF�׼2w��+BA8%KoxR����O�DU'���@Ir�=�j9~�� �r9����sd�����ُ%�S?�%�&���S]	�<�ծ��S��L6�Vb�糒g�ʁ���G��б� �N���R�h�fI�ٚGl�aʳ'��[��^�����̀)50��*���ǝe����y�l��J�1�Yf�B�Kɣ���l4n���^y�q���c"S�.}�2�J;w&�[�
֟��&&׮��T8T�x�!y){����A+)պ�+�%�JS��ߟ�~�H�	&�`�� Ϙw�t�A�$!�þ��$�S`zvZ�1���h��^�D��WS���mN
���QP��Q��H���u	�~��1=n~u�(��F�:_q��;4�vG��#Z�
�P�;<l����^_',[��>ƥ��4�jN]9�w	�L�3a���X2#U/��wD6f獲�g��u�W�����FIVp��j�5��=�Cb:���3B�$j�v:�3NA�;ALB�׺��6���
�$&�>�:Sq�e-ˢ��N�ı�g�R�%�rd�a@��8rz���;݇l�ėh�ac�����`X�E�}��%�"&�L:)�8���lf�>^��[!$�o�09�w�LZ��O����9�ǭ����|`cE o���Mp��>?��L��Hiӂq��%�f)n���w��ء�=^�/�G�y��"�g��嵲zy��5�w��wQ�F�����K�1Q��ǫ�7��'��m/�Mn^]P����g)�6L�q���C�$�g�scg)d���9:����}����~�%*~z��`��c���J*7W���6t�qG/k4*�����P�hڛ�����B%SC�wP̻o��a[�E�辟m��%d�$^K�ND�M�.�k2��p=}�0�:-�>-}W`�s#T�8_~)���A%�H���=�<Hf���
��4\���ڽq���[�d�\��Z�\��;7{�3��;�8`���Pg�_���-���~82@1~��}#3����%�b�oͺ��Qmf��X�����D���h��T	�@��K�����Q�觴uuZ]8�����ʼ��zh�����es�鍔�..�)��5d�����i��"y�@gr�x�B8��7��'�5-��WtoŶ���u(���t���nz���H�����{��S�GxrH��Ĩ}rB+�l�L���X��BY*p���T8ͅc{W��M8�9���(C�-���w�y�t��6�=|�$�現���v�"��wM�k�TUXz���U����Aw�)�I,�Me��Ӥ�%����o��f7ZvG+ߎ�y�x��x�Q�ό��?���E)�?���b9Έ�Ӝ��o��T�U���ԉW��WX���ߜ#e�b	q�_Ua��rά
T��C��پ��*ꋈ�Vȿ<�U�Bo:8
��G����9g��I.���oox��u�"�����듒�Ү��J�w�vh4���ˬɘ��9r���&C��~����C�k_|cBb�{��gGX��xmu�dM��S堻>�xoI������^���\���<Ψ;p���I(����c9N���q��U�X�G䢃XN\���Zv��H%UW�V�a�A�P��j|vb�����������Ki/���ƹX����<#A�]��"o�5�a4l���M^����RGJ��r�U��!����c@V���D���y�e���e1�hɞ�_&�$$�R=z����1^6=��}�*3�a2V���Ǹ&������|~��dh����JD����٘?&�O ��ߩ�x�y{M�T_�A���p&��ZzoG�����wkd��a
Q�S��чz�!fbRm��Ɇs�p#�qi4����Y��ι�ECY{�.2��L_K�b�������>�,�<��ʩ�?v0��qP���(d���k�U
҈��=N�fպ�vew�(gگ�xH<��kfR�L��"wVA�u��u��ˆ�:8�w�r$r��ԉ@8B�X�p?�ݑ��k$�>�<���ATG�*��'�t�y'r�=�)D�r�@>8�\������a�ШvB��	)�L�f�\c�$�)+m�-�������pӢ�!	�nW<�L��%�p�@�A㶜���xr��'~��[���#�dO�0Vw��C
�x��g�Щȁ���bK�; X�A }.\��$4�F��g��n+��~�j	��I�-��%���^�Y.d^�3�|�vy!v8#*o�%W�K7\�K�F�bn���$�\�C�I�/Z5���2�#�x���@��ȼ��C?��MD\������	ԶY����/���)h��ζP�v!",�Yp�t�q=��oޅ���v��1/�>���=���fz��3`�aza��'����(�l"��C4ĸ�Gn�*�,�X����.ם�n��&�5ƈ2�NB$K�%�H��AKk<���JhF�~���	4��)d@�T�U=҈��/�;^!/��' �-3dPϗ&1",C�8� Hkn���1��o�&�GP�ʮ�) I��F	��m6�$��I�n������&z��Cu�4|�Y�<��pu\��%U��ȱ�#+�R5�T�ќ�[2�9� ~�	7%�@�Js~!�	�ذ�"����g]�W�8�}�"c�&BY�K������,v%����c'��������VC� ����@�PT���s<��������5�f���h�V2O`M�j�gAɕrU�X��i���&�,��.r)�|1ᲊ�<�6���Z �)��l����\�Z�z���fla�;olp��4+�~j����'���L��B�)<��J��;�����k�����f�s�z�b�s��A�\k���3�aW�}�b��35��bj�?��8�;:�$�r������j�x�k�a0��%\	baoY
}������{PԤ,"���n�S^pQ�Z�iYU�~ �{���|�9:�������Τ(�+�0o(��>�ߥ�vy|�uۧ���l�?K{���C^&�L��aa�T�1�H?�=�׉�&�_��ΫAm�T��յ�j��^b�g��L�Q��z�L�����&O�6^ȚP�������XK�����>=/�@�� �l�kvK�ܓp�3�!DE��(-D�q��0W���3x�_�N�2C���K�CY�V䢲T ���1���xK�IEE�߻�@*��f�v��荼��(�B65����Ryn�b�=�/Y*+�2���檈׍wBV�ϖ��<�n� �e�	�f�D=�&��8N9q,/���@�?����G��͊�7KF��ye�Mn�J���RpY[lUì��O����њ.o�~S�ze��/�H<�.�P��\�^��x_�����M�/u��ȴ�5>H��������h��%��������M�!�h(?����)��u+�N�A���gq�$7y�rc���?����2a�=���I��lu���*N�mr��~4@�N����!�e�>FCi�gqNG	b
-��.y��Q�Yz����f�6��/��`u�0xH��){T���I� �<��M���Ka���NYN[m���C B���x�<b�����wk#lOa��J-E�33m����r�IZ��4�G���xݐ��9�ӐPJ~�w4I�Qy�۩�?��"�P{���hA�鷅�F��!�g��Q˛��g{Kt]��MJӹ���	��Sa�;�?��'ɰٰT�\%�����C�dnai��P$�>D爟RH��e���,N�� �!�_�_آ���c�;���e=� Q�9 ����;G��z�t���zx���$'$���4��AR���w���]�Q�O��z�~]}���Eٟ�h� �4$� 9^Q���������3~��S���O�(mфM(��N$�2ߴ�>�m;ôU -Ѷᤫ1�I�n��MK����0�ր�z��&C�Ѓ�D��r��V!�u��V��`P�-7U�MsNW�R#['DyS��ƃ��j�"�vψ�c�@���?n��� � O]h��sf��c:/J������唉؊�
g�`jD�7d�n[g��y�"�&p���z�Ld�d��`���Q�@e2�����2~�������y�I*5"^�yc	v������1i{0 J\�.�]#��W����w�U?�����QK�m�݇�m}t¤�z�t���?�S�����3�w
$ޏ���%��6@�L���M���Z�T��i������|�omCy[	)�`�`���a#�{�����K�����1K����K8�19q��m������,�Y���ɀ(6�u�ȶ}2>4��ϋ���'�d�ϔ���M݈->�	S��h�k'Pv�(��ƭ�
<������]��p`���L�*�/ǿ�^�́�)��t���>]UA¼' �7���2���<��ٝeq�S��vD�����?B�נ�3~�V(���07js�_�w�v~t�6�@��Q��7��yX�� C���2ڵ� 4�T��d8l-Y�(�K��2N����|�Xf�17��r+bb�0�߬��&%���(j���T����i�I��!x�$m_����H��ܸ�׹��j�io[�G�����e��$r��
0�sP ��AՄ[��s����b�p��=��[A^2�I���8�Bń&�i3�HJ�!T��]a��^�mI��R��f2Zx5���%�*z$���dw�fmTVQѹt��n�O&�`�~0��tw�{KDp0[����.M�d��es?�C�gN�M��d�պT�]�߈q!���LƎ��8qG����c�gM[�\�m1)h�_��%���nv.q�Cv������\ nNF$�%NT�J2������%!Z��pKd�}���+���~��(�]�(1� �B�[�$���caS�� D��?�
3�Е=n�p���o�]r����^0yl�o��x�$�s�Q��c���*�$�����:���/S!�@�0��-��R!�6���|k�ci��U�I��2 j؃j�\��3��k�nԽ1w�]�"�£�����Ƙ~�hk�ڱf�nе�-���*��i��n�	#6ķ��|��e�/qb͆�j��ey��w���kE������z�I���$~zW��R�Iz���ۣKΫC��q{��X|�I�z]�a}Ř�w��s�� +��r@˿_G��%A=�����>L��8�K�1nBw��L�u�M��p�RO�5���4%�O�(��1U�E�s�j�
LN�
L3��_���@�k(�ѿ�9�-��,;l3pyoOc�A�C�X�+��W��]��m�>��f��E;�n�E|7�2s���k3�l7S���Cx����.�I�ɜM�;���1w:4~ى~����V~���?�G5�z��R���$W;�C\]��zu��T���n�����'���<�[o3Ƌ��n��� 4k˶�|g�M��\!uT�BNy!5���U���cp)�aQ������j�,=k����=����(j��Eb����1�ϋ~�D5J�֥>��>��^�f����N�E(M~(?b������~+-Y�a�qm?�a@��I�"���L�k�gIu����˓�h��&�������y:�]Ac��v�e0:S��,�?�:D�Z��G����@��\d:�6A_G�J�r¬3J�MW��8ϟ�$u{'���Vʱ}tN��g5,Ӏ&�8���Z�Q��#�k��Ղ�u��gM���	]	�py��9<=�J���ʻ�z��R~�4���˞\»Q�M�۞8X���3����W�z㻙���<b%�詁��j��������5f��8;��@�eǠ����s��Kz�a�ԨyPW����g��wA}��s�7����PW�m���Ӓ��W�Ӿ�jm?$��0�UD��2�*&����b�3�}��z�\� V���&�2N��@��f�;0 )I"6� ��ߕa9�f�e�72T&٬ʨn����d��"�͗���$@W]��fC����cI�DvӤAUZ�Ʒ (5��H���x��u�J)-��ꮤE�AYj�l���$��� �;�y�ç�N��#N��њ�$����K2�M1����C������cIcb,����T_��}˹��C�'����M���&a�9 (�F�Ws!J���h��eY�D�C:z��$�ڧx��G�0n�]0����Y�^ 3£@����%�Ÿ�Q+p��IG���W`��w�xNA�G�z 6p��A����j��{�7+��(Bq�@�`(v֨�n�����w��d�u�,U���,�"���Q�}�؋��S%|�߂��ah�y&80�,Go�Y�2��	�
i-�0���9���y�h�4)�P�����"�e^���|�c���V�zL�ch'��5�����(�*�b��M�ɉ�>9�v���nAs����*^k�������ń<�h��1$6��L[�o�xr�m���j�	}��6�;Ebr$Kj�b<�� c�D��)/Q���C��[��^425�L7�T����ӎ��
sҖO�1�{SZ3�������P�����3�/Q�1�bB?�f��G���՟�8nB�ڇq̕詷-�d�p�dI0�FW�r#~V9�í�o�1)�w��Ý�PU}�e謂T�ӿZ�6� ����� 
��C�BF�g��5F��-M��<�R�>����q��ɝ��˅��Eem�@�u�b�R�k��B�}d��z#5T��4�wh��R+���Xh�~�7�����L���GUAЉ��+_-T�sK>��n��A'�� h&�B��*�%��oVs2_���S	��侲P1�M��s�&�:a��:��1�A3����,[T��h7�);�L���{����m�N��n�OI`���?�06�EV���b��<��i~��%���m^#�'>K��J ,.ߥ�c�z�*[?��w���j2ԡ�9��e*b��7.a>]��*.rkCU��>�b�Y�"k\�#�!�<X���&O�-!��:j2��o4c����K����1�l�ϣS�\�.RA�\6tR2�f8�ePv=ف`F�u¦$�6E(#�eO����}'�&@���Ӊ�{��E1$hQ�����"�7�M��2&k��c�q=���河����8�X�f��P�����
#G���������D`�C��mv��"�X�XK�^��$�e��0͑�x �WUl2:5S�t�U�I���(4O])J�#�`�^�%p�A���8j�"G!����
>H��0�o��P�j���3��N��3��%�r3SA޲�9cDBh}D�����I$('��º5��ꓞⅸ/'B�(eA3�?=���Ӝ��c�C�:<�xl�+��g���>Ww����¹C��1��-�@7^��h�[ث����	�Ik��3�=ءl�E�����"��*�3��V
����&h.�|�7�j_�d���infӖ���II��ܹ�4o'zкP:{ ��0 2��p�ᰶX���DrW��{��J.�j�=E�H�P���I	m�@M�ӌ��ە�2
�<�B�X�K�y`�2�q�Qi��R���˒�JZ�O? ����d�{��P̄}�a�#"�&r��k��^C!r�RW'�<IJO~	�Kʇ��
k�c�;<��T���E��J�X�9��Q�m�;�rD#��ms�@�����A���#!���sƄ.��˔�X��;��[G^r��6m��7��34=J�8t���{��7��K�4�C�ҶN��*J��X����~F��ύ�[��	�]m���PV�2k1�F ��2��ζ��� !<a�>����Z=��nIs1*��![9S�r�w�Ld����KX	�r��L��n/�TA�]L�}(n�wY��؞�S�ֱ�Y=r�C=���@���f-~�E9gv2���nW���ɷ%���C�avF)K�-�׽����V�2���: ս�(�c]	�9ۣ�K,{j�h$lH���4EZ0P�өfg�v��)H}���٣1p~�6������Q�_�NC`�4Ll�F��2��������6�I��G������Ǘ�!a4Tq�=�.��!�5��p�&��l�+��{��d������}B]~Jg5��(�2����|X�����?��\O�fڛ'N4��z�Vx�]c��~�)��]�����mA��	{c������=�r1�j�f�n��g|��g���R���,2B���2b�� ��Z_����ޗЇG�Yt���|�Fi�	��H�អ.�����']پd`�4|�K_X�e��
��<'7Y1\��������HW
.nC˂\h/o��iW�7�����}����E�K�?AO��j���{�/�;�"�n凤�����;#?.tX�׻"a�񻸶	O�K\�^��;��O����#
��S�mm�myV I8�Y�^�Y�g�N�����ˤ��n��c2[�Ţ�oѯ3�MfF��b>V̦��_Sk��C�Ow�>~F�#s}��wJ�575�{��v�J�v̂���̔+đ���+�gs�l�}k�o�zbK+����a�H�4�k����Y��cu�҂�Y,����tb�����A��rQOh\��G7����QZ~�m�$�\�"{�Q�1�� ���A�L���*��x��
 �('����G.lN�Ӛ�G�~M6 0^��}��kU�P��R���z���ZϤ��hvSҎ*��8杵�w��z9���N��Fe�HrXUO!1<�`�J'�4۫�ag�GM�w��2��7I]0l���!��8M?T�,���E\��{S:�)�r{n��1l��zG��"!��%u�������q���S^�����.O��O�����T��O}�	�qF��H�mƫ$�)�K�Κ��<:[|S�ߪ��r_���<]؃���r���m!�8gE=3OМ=�]�b���"k��b{���E�ĒǮJ�(P�>��M���;�v��H��pPL@qTO�Bu��+������%�hm�u�Zo��=���o���4�f�R��`�O4n�3%-�'%�f��#	>ʃ� �-���?��{���du�G"����l�6���\�vB�"-F'�|��D�&� .&����@7PT���z�Qj����Ty�$��b�c����*���}\!�����R�4cQ�7bh��~�l�����Iy��Ut�<j8H^���O���GX�3���,��uM\1I�l�yVD��D#s��z�A��:ɔ��d��9����׾�H�[lEӟ������n�������@8ȝ^`�am1��䦺B neY��;��^\h,tj�d�a���:�盪��`��u ���S���4���s�=	x�#�^+lc���g��-ls5T���9i駻.k�>��_#@]��(nC8������νR���g{0�k_8C��X�-`۬��f#���a�l��n�ǽ�۶�Il����Ӏ��_���hL�a���n� #���)U�!MuU[�|t�����PX�O�b�%��V��7�ɟ/'�U����q�-R-c�@TmB�54��B0����� q���
[�]� �F�[��O�+����Pܿ}�0�fvd]�c^�*�#_�-�RWj����v\E|��\pK����S}`c3T��㐬�+��.�w����o�%�{��y6�h��%lM7�� �-�I{TG�~q�E��J`iʾ���η�ѭr�"��wIM�]��P�\���VJ�4%�q���t#�X�	Uw���t)i�����Qں�v�g�3ș�"9C;S�]"��C ��.�������,��P{ؿ˭�A��wkm�B����,}폕+�~�= Ī�^��k�։�a�|���LJCæ>������,ؖ���*�&���C�.���{s�s�eQl<���"U�&��HSG��z^^a:��6��=CJIpbaU������'�^}�lҽM��H�i�
�YD�,q�U�4�áz*��'�	#�$`ͩ�&?��1���6N�q�sR��ķ��7���u�&J=�ӿ��h���oFo��D���#�?��w�	r>1� ���4 ��[[�B-v%�i+��6�d��A��՛���>�J��m�!��uc�@b
LQ���΀A��:��k�	�ף��8#�W"�.��^mH؃���Bu�dg�ˢ�{	��\%I�,+I�!��b6b�+��B籮�FŞ�>�y���4.�%<�&ڠ���OO��?}{D^���`<b�;�Q�[FQօ�?*��`���)�y^�l������l�'jKo��`vq��V?��^U�4�����&bw�V�D�E��YVۃv��}4Tʸ�����>�a�-Z	ut�����s��F��#gV=�#"�T����g0&�%P���1F�`�lj�rm�4`\3��י��Җ�0ߢS_��I��|./� �	�_%�>�N� �w����\��I���ew\�����`�"�l�^��:iۯWԚL��k�q���4�������e���S<@:��C��Ń����n�@I��ȹN�z�`j�)M|x3��8
M1@��l�B0N�{�֠h�0�F�5FV�a�!��N�Bh�>�١���8��j)�wz�A�[o)ž�D�_��|��z�B��'i��������OR)���6��@���/2��y쩀�²
_��i�����Q�	��/6���'�;�Z'�?�O�C�������=��iob$+<{IU��n��'�+�Oqd����C�7ǡh�V���"�e[�s�E��¯�|&�('���쁦��Ia?���y�
r����	��
Ur�L�8Y�!C�*U���S1>u��9�s:�Ӵ�B�k�3�X��1�ԫQ�aY�˶�9ٶ�d��0�}b%�c�P�:�^������	�=aw>��(l6��:���e���ٯ����#U�e���-$O9�;R��oCK��:�$��QW�V^t�U�T�.�d�p��@w�/�D�̚Į΅��:�!L��sZ��4({pW����B�v3�p?�(�ܐ)E�Wx��qУl}N��[�a�T�ϙ�ńU$*7(��ǟv��H,0\�g��O}r�O�o=:�g%�]{�c`�����������ġĺ4�!��#l]��	�RU�]��i�W��8����;5a�v��'ȗ0�2�Qf`8
Ү��_�8�_�K.�Ɉ�s��ԡ[�j�_$�4�����I�!���u5�x-'{O��h*�v����;�����t����D�Z}h|���_����+��kR
:n\fg��w��05��=�A����!/.�4ꪡ
��PΫG�C	���cBM��������u����I9AF�Dי�~�k����Gg��e�([.W�I�8b�;3~r�d'�
���#����\�� �8��d�}=�s����ȣj�r�~^�W�~y��<��C�}�@ZLX#�͸���
PxW��u����<��!���!���ݰ��*�`�M:k����}���*��I),�X���$ٚ�B-�o��"U�m�g	���OU�L'���w$nZc D��/Rڒ.n����,E�ce�s��I��]�-� ��pg��7.��B"�F�#;ߢ�����S�I!U<�L20�)���� xA��,#c�����,���j���l��$O'�A��l�K�
�*����Ţl�ŧa��r����3�i�>^�c���(��r�]p	��g.N�0��A�|�O�G���Ɇ�$z	�3B����k ��n&�ڟ\���Xd,�R��LXȹa���O-|[,J�($�߄���6���Wh!r�d#I$>��p�̄ѻ�ݱ���z�sS�\GV��u4w{���H�z@٢9|&���R
���\e{y�=W����� �i�`�(�j�?T����3�#�ޞ�B��[���@t�b�@��e��Y�����+x�R?��2<�?�;]�^��>|�ܫV;T!�){������ǔ7�:-0�SDJ��	\
�ԜN�)ٰO��	�y�ܓ,2
gI�ӱ��75�s���/��T��]'GӁi1AI����[��&~��'��� s.�ڿ�z��t	h��ʑ7v��Qˏ�X�6�m���ו�jeC�)[�vGb��Yׂ ��!�fSbc�D7�gȰ�8��9__�d'dp�@uc�� 2���Qm(���ҿ�G��i:�%5�8R6ŉo�����{V�!��az�[��r�,'Q9>���[���f"��e�p��S�\-��u��]�|��a��چ^�I���v�O���"���2"ヶ�����;���0cչ�M^�O���RVy�Ӡ��F��[��3�xL��|�9�p�+u���>��x�B%���Nk%j;:�f |�S�f)��Q��N����,�V��2!|�qv�`t	>����Yz:D��b1�#<�ĤH ��IU]9�_:x?��d����h�����[�#�[�r����*@ E@K��ωZq��W�|mi��CPv�\e��B�X�H�ן蠅�ߩFhw��-F�jr����o�[]��PI5��3mP���y��Mxͅ�a(K��F۠|8��a��e��j� ᨡ�7�[Ŝ21}��J3�����FSK1ѥ�RxVA���q�Ď"����Lmv�{���8 ��W��VC��X�{��4�6�+V�3~����y��1TL�5�/�m���������[��rA|��[`1y s����=i%�[��ٯC��}��������F�5� r����0�����,��)��n��J��ט��|Q����;�Z���x�+�o�����A�"(O�W�$��7���}_�yX�6fW�^��B3�U h���z�"h{�9P����V e�>3I�n�����q����AF��ν��NMm�}��_D�Ȇ�fߐ��&��[<����_TA� �ͮ��6�h�H�6�ǻ�p4�t腉��R��l�m}�|v�]��ُ�7+*�whO��i��;Ui\�,:HT�y��X��������2���;���,>��e�d׈�sp��bZ�郁O;W��/�&o	H�t.t���7F&��0�$���"������8�;�ԟ�hY4��?�ʆ{���\��S[2��O��*.W%���L��!���NQ�UP0���W��M��]]��Gw����(�J��%[W������ n22���LY��c��gLM����H�s!��:�7�h�xŬ����^V�O2T.�DxQԵ�M�xF�5�e��W��c�x�(���u��P�'Z��z�5�ex�
HgD��������_�ӀY.u��+�@���ۉ_o�����aʹG6M��ZG9���n�����= ��6����/�m������/��P����qC�.g�F-%��r�,/Q��R����v@i>��������	1�Q� ۥ�aR��Lc���\�M�F���c��$�99R��+����0��T}3��Ŀъ��^����	�W���)/�Nj�:�`x U1�sw���)o���w�q��$qP��(w�� �j���u&���K��7�7�Q�l�����B|)zZ������w��Y�rI���ʢ�6��חv���E|����/"�b0�bP_;P��w0�	7ϷZ�P;&�D�ľ�R�dSh�q(w�RB�R`�|����޷Z��[���w 1o2�t^"��W��=�A�l
�XX3��r�,
O�.�֤�H@o�P[�UAM��'�� 	Lf��;���o�;A�.�:���0�`�F�r�>q��7ߖ���M�s���O��SÜ<����vs��#]�¼�xd��D9��9�����c�O���y��N؂��V�O��8�C�'"Iy�K�H�i����ZFD�m��C	�x���Fș��u@M�C����*��У�s
I,�`Y"���� 6�K��n���ңA|��X~ -�����/�a>��RI�99B=��������,����ߐS=��DL��U�C���Ѱ�r�i3�7�"�ă)�؃N^K��v]����s!��[��P"�L=�7[���:� d�Z8��T���x%��H	������h4 �]D���u	h+�"|=j�UT9Y2S�9��9��g��)�?�K�dX��/�}b�[�@�BU��/���xWv�i�M_�ǰI��#��\ݬ����+z��~y��>ü0;}��4�91Y��O���q�Dx��X��1axSfT?��ab����i�'>�Y��#W��γ��]Z~o����f�p�ά�S䥊��)��ݾ|�<xD��FIc�Т��m��E�b�YVi������Œ�K,e���#c��S�I��p���e�ӭ�c�acT�|����8J�4'j��-�+I!������Ǖlԁf�'7_mPӐ��Q	��Y�G��F����9�CX)�:���sZ
�w� M��<�~:@ʫ�-L�?� U�a����T�(F�^x�y,�F4�rwC�b�;:s׋�Q/k��$C��d-ԯC�SSx���p���9���Gf��K�0�2�.���`O���j��������p�5�&���9DW�zAͷ���23�ޓ0%�b�����Z�=��U��gW��VNN�eVj'x
�����:;%ܛ0�i�\%��Qc���`��1"����􆵣���/��q�K�8E���G&ek`��;��-ԩ�Ua�ꛊ�zW�4�w[1��B$���_����Ol���C��� ���^I�	ƍs
V�șa=+��
2�S�v|�m�ۆ<Z��GP�����2�w��@�`��)����e�s��7���)h��e�)�������E� ����#�&�t���'fd.l�2�� �@0j�Kjwވ��͓A����<����_G!��܅nD j�,l��W��v9Z@`)�z���j�	P�;t��P��4�RVX�:}��mQ��2|�ՠU���l�-�5�58Ȟ8�յ�P�KZf'?ʟ�j*��cE�g�0�{Q��B��>c���I���x���Gq_�"� �e�a^Tan�J��\����ymw�-NRf�<�r�C�q�ļ�y���|����}��͑�������R:��1��d>� ^�x�@3~�����Z�e�� )��m8���^or�[��C�	�,y��['d_�ᑓAvT��c�`����o.vE�#[��i���f����Y���z��F�t�xC�vc����(o�l=H��N�싌Uj�$����۱?p�P�`Pl�ᨪ6Q���~ݞ���{�����g��~�>'O�7��ウY�2�P��@DV�θ�I��y�g��qT[nv��w�����(�8?$�v`��$A��T���HM^8��T��Q5�y6�\�¤�9;B��eu1!��7�"e���M�r�j���wn��,jA
�k�bݺ|w���R�MM��^R�	�� .�M�G%��ܱ�ʫ���M�V5�ݤ�(Ks�IR<�7��ʄr�@��=z���Ȳ���EQ��G ߨ��`�s�_�i6N�eѩ�*� ٌ&�����h�=���mnwe�N�|b��,ꐦ���͞b	d�Ѵ|tDu��X��x%������tE��_��������I{�����IB�~5#��h|HQA�N?�w�W�Rj%�b���,h�ئ'ݩ�=��Sa �u�u�ֺ�b=�f�	T6���0K�X�H�x��m}`��Dc��{=��ˌ���h�t^��Z�`f�԰��̒�m
�
�FZ���M�%Z:$�>%���i�m�����\����/�T���Sv��2u2=�/LS!E (��t��xw��^T����8�˿"�Ƚ(w�]���#���w]Trf�K�7��]�l����~l<�n4��g/�������ka��޶���#��vL�Ad]s��6M�:6u��)�9���j�F%��h�����9�	a�����Q��]X��B���;{O���r��J���;��,�>َ)U�U�7�0ek�i�!�$����P��tѳ2^���_�����H��~ٝ�f|^ܐQ��D�em�z����������!�BI+o{x��~�Q�`�D��`U{4��_��.o�����DO&)EA��J Wv�?(%28K�L��*H�K�!i��t����+������@��C��ǒw4��u�x0�j�A����}������q3Jt>ax��1s�3�M��謏���?�c�Grl���\KəK��BG���+��#�d��J����*LŎXa�}�C���<G�g� �X�6��`~݌��s�2@Z����\���}�Q���z���f�>k�1'�&&⮋{�t�2���|f�"�S���r���FlE<fyk <�BuS�>�D�l���ؿ��`�$�(ZWL��27=�|���M�!~� �=�el1%�x$�ʭ�#�ꂫ�D��8�یg���sb����|�mZ�2�7��m��8�E~˿b#yG���둈aO�_�x^ܴ����[p�׽���d��[��ST0Y�oY��c�{�O���ϕ��D,9� ;s�������@�V�#+����k_Z�/��%."�g��.4fv^c>�H <ұ�?�S�@p��]�,c�L�Z��`�KM�,9�Q&F%y�Q�.���`E��@AoD)4}�uϛ��l~'<-�/7�;�q�oFe����t��G��(�m�����?b5 �c����?A���]�.Mo�V��2dӞ�IZ[+.T��t�r����H�)�*�z��<B�䪚���z�b|Bm��um=�η��b���4<�3��g�����n� }�D��"�j��TY�^	��𮇚5W��H�d�N��#<O7��Ugc�<���4��Rg������
��_�.=�>ylQ��~6�����1%S���1�J�s.z�^�Ϟ�rC��^�"HE�)���M1�� ��Z�q���J9ñ��>�T�[f��O夙������/�xeDl�C�3�����"k*���(wjZ1,��^G2v�:[~����1�9%��v��/�H��u�茰F_Ts�������L�|�����z.di��)�n/�@NO_䒙� <����~�7ڛ��q�c�l5-y)�1EH��~��}��̉�s�p��W٥qI��Ņȵ��	�S"[��D\� vg"�:�4�����M�������fx$�:��p;d�H���_���_�Sz���x*4��SfF^w{G,R�v^0A�*c�'�U#1����+��΂� �z�h��e�t�(�����+m,H�[��F���S
'�ș̂V�/C��
��A%�Vf4eQ^I����8R���'��`@�^Dơn�>�f�Zw�����7f�JY�қ��c�	������i:!�ޠ�|n>���{7�A��$� 6xXW2���.�tN��дaJ�e�+��3Y:�T.�nLr͞�d۽{�+�4�{}��\^%\����[��p���l�wW��[�"�:b�o�16���	!딝S@{��&�Buw�,�C����_}#�<��-��9�܅Ԥo�_���e\�l�J)�H"8�����@�V�Q�%-"�����N�ϙ��p���9D�I|W��T_��?n;r9艝2C�+p$�n���
q�bS���F�����'�d�v/���-խF�0病p:�8v��8dлY��pM�ġ�J��
��]z�#YK`G�P�l6o�ij�o�z�%��#�m����N��y�ly�Q��,�[B�U+,L���d�kze�,Pu� �Q�����s�wΘ������1�&r�:?��h�&��80��r��S�� H���h�>�n��2u/w��YX0�i�k��݂�D���փ��~�!-, I� �%(s��jn�!��{Wl�1��d�JB���#�{��f��o4�������p���4Y�n;���*�x7�{� �*j��;�	qr^_:U��W^�9�O?5�&�e[��׶ ~����9B�uX��\��N0;n]ݭ	=Rq�[JV8p�.U�|XaK�q�XTzQ��C��G~���r�pN��-�T��iNq|$�6W�1�/��E�\����T�D�2�������hQ�icT�d�&��s⒂-��]50@������ۧ��'���j���zbjn��Z�Tt�:y�dG@Q����a+��aEݛG�eՇ酜����T����iK:F,��c�sq�=J`8{d�a��X�-m�9��cT���A��u���9��T��n6�V,���}}2� $�u?%�<�������4S2�ƏY���R�U�??ԈX�[řt�̪��U����7��U�PR�c�RDEc��W�a��vi[����0���b3�<��lX+��R���������"ǻ9��ZQ>U�Q/ք%Й���o���[��!|�ud��Eo�(����&��(�K ��������PiY�y�|��h�6	n_k
�٣}����=�X=�;���搚��0��;$��9�yxb<���L%��죌)l��H4��RLb�mE�p��&��O��!�rj��=SF�'
R�R������ڇߒ:������Ge�%n3q��Č8��{��h��?�j[�Xq�o}�0�9���K�VxD�\��eyB7�G0 .Ћ����0b&�-����Bׂ2��"iĿj`%D&]��j$� l�2 s��k�C�HhW�U���1�e�v��s���k��y��u���Q�xd�v�)��������!`����u�!N���q��f���$���8;oa�tϑd���j�@�(2,Z���-�ǣ���w�Ɏkà��m��� hH����W����s!�BP���K�ɨ���z�$-�����-�N�8�Ty7m~��X�5	�i�'�F� 
�����6�56e�{w/[~�>����c.{���`HB8}ۆOz�:IY�\���v{e�	�BY�1�Q��2�]y��+�Q�4�?e�?f�8&g9V��}�����go��r�@��_I��q����w�,M7X����.񀝒`ivi1H���I,t>W[\����k���$7������45�lKK/�z��zXzo��`�[�-U٤8���� �P�0Kf�Z>�:�<�;s?ǋ�.$������?n�2���Λ61��S�H���L�0�NOmYf��Z! ػk�#�>8ż��¨`\��>��@��0��2�0dd����"]�O5T�֧{TXK!4�o�2�b�bh7���f�ќ+mL�O�/$)�5=ͮq�6c̸���ͳׅ��K�k
$�j&.�6��fH����1;�W�5�(�P��C���xVY%������f��t:7��0��(�BNY���Xay>��w����O�~����t}�XJ�z|��;>B�ܣ+�\�A�f
�L��s�����g�і�iIM�VY���]t�o��#O�k�Vo;�b�ϊ|8U�gģ��(�s����Vpc�"'٘�!%Ե�����y_���J�����I��8�զw�RE�B��s�X@-,�o��f��Q1�����D(ݑ�к�y��٦���l��ȏ��g�=ў�d��Gv�1������lFK�F�.��i�B��TG^t<_F}WN.��ej����3z����=�U[��ڽ+Ž��D�D��L4h�&��p�w�p�ʖ*�%5��\x3t���o�3��KK!�[��^� �U�[\i�6�V­b�e<����v;*@��5�ľr!̈́a�6�xpv��O']h,��7N��!���k�R�=is�#IT���F)8j�lq�^����������ap��:� 鷮�6߃��a\����o>'9�1XMJ�O�>A	E�v��+?i`�Y�3�ˮ���@�E��W��[�`�Fh�dw�P^<eDؚ��`+�S�9m�ӕ�)1h�~�g��?����*�>mM�b_N�A:�&ߡ�,���'|U���=N�Ά��W��Եr��1� q̍J��r�\��Ӎ��j�J�'<�
�`ʠ��^����4n�_�y�T7���@�|!���������7������MX�����a�vMEc&2�O�f�vq,��L��ŀ(Þ�M��,֒Hw�㦈 ��~���W������q�*�79��I�37����N��N�`��]R���Z�<��^�ު�ӯpb?�������)��2�sG��v�����R�M u���E2Ap��y��������oI'�4�>!i�	�y܌\��n#i�i!��z�E���u�qk"/����P�����y�:1���B�GYeX[�p�����$�_�k?6�I8'�Ju;U���~�$;�|}h?�k�ޮ%��by1���N��5��փ�B �-b'b��h�i��V[�ﴀL�Ş�I�$YIz:��0޼�/�c�fS�,���%�%�|B���54�?�t"��
��"��Ɗ
��vDq����9_y!L�[�� ����Rܦe�+LZP���.y'�� #C˵�~������[��������,O��UY95�����˦,��?��FN����N�Qe�(4 �o�v�#�6���Bc�o�jR�+ģz�ы�x������?"�2.8�츓�����A��B�x��ݬ��e��G󹴿9W�]�0t����)/,Sn����B�,j#>�G[1*s��UFV��!b��P�C�~��Tc>m<�<>*�z���n��ʎͪ��y3P � \a�17&�!����H�f׈=��`����6�ȿ�����	�]}��[�z�L>O�����d}�;Nx���Q��{�c������`��^`�҇�V�E��7oPa݂����,KP�`#��3��X�jo���E������1wcÃ���������j��VJ*3��KT����iѹ�hZ�c��.��K?���#;�w[#��&)]���e)��:O�E�㎴��Pf��R��c�Mת���9�Ў��~���&>�B��cY���ÛŦ*�;P�	|s��5	0�['���ɩ�ŋ�H�ٱTI�e{����ps;�T�̬��gm~�]]+�ԴF:K\е�Z$���,�`���6��l.L���J.`�w��m��F�x6~�c�ϝ��s"[��HZ��dƿ/W�@�ġ����i�J'Ƶ8�`�b��8R�\�O���3���{�D��{�K)9���y
G�?�20` ���>C��1���J�������'D5}7u���8Cɍ]2���N&.���l��0c"ʴ1�8t\���p�����}{�&�g"\�w������}����A�c<�R�h.����֢&����-AW�?��.S���?t���~B�a��3�3މ[s���`���*�]�QHחK��h���\��Q�)U��O\CɖV���i�n>�cₓL�ip,"U �?v�|d��S�`�"Kr�v��4�eat8�t��yfK8A:a ���X��\�옜}C�U�]X�xa��Vmһ��r�8�9�3pR���Dc�R�Ӗ�v��i�)ȧ�V�����/�,n0c�
��[�۱�o"�͍E*4��I�$�ut9���t?
-�9���z�{��-2�~(n��y@J��F��B�u���&�ih���l�k����淀d||�&�bO�ɥz@�x�;���H��uW\3S ���M���������#R�y�41$�5�8՛��	Ƽ 1���\֫G��KOSm/��`a��E��D XW��T�%՟\�^��	�,��
�NhWy��+&Eh;!�&q����:�Ʋ%�qOV�`��d��%�JG��O3d�*&�|{��E:���Q�a.x��Y�h�����7�C�DS�{6�̲TIv�W�X!�"�����4�hLt4*Q|���!�(��X�[+�^x*W����#{c	-�3P@r�'��۱�����Jt=J�p� ?���`8������q��h�t�F*F�Q���@Ws-}C��X��	z<%1�oW!�1tq:��JK;��Y�6���$@��^CM�����bV���������h�m�U/���ୀ�Z�y�;�}E��-{-m#si
�ʓh��r��
�<k�4���T��az׫k�އ���ε6��9N���,�~�8i�OJO�Ů�n���������o�x t�}c%N��g,�9����Kz�8J3�� ��P�Z��.�w� ����C�-�^��~�T�WS�ȭ�	i�+� ���!WttV���6���w%�XWW��x�t��(d��t[��j��'���H,����`mleU��c�V��l��T�ء�L�9�� P�	S���L�	!*m��R��R�X�@���y%��P��+S���.zI���UCo��e�,�g�l����3�n����c!Vt"����?E�N^٩@���H(L�&B���@	k���a�	��nk��Ӂ
���C�e2=$��M�f^BlL�1qh�W=���t�[�%�2�|�P�i��@�+�l("@m�+<8��$����q��ΑG�:Q(>:TUD�c�5Z!�am�\ �yBj<�����}�U <�#����9��4/���+78K2�z�~�g�bX	,�Y�K��ՠ�W���q��eQ��#���k�F"0ȯZM�qay���u�yO���mVN�H4��vΝ�g$�����refh�w�F��"4�פg>�_�.翊��ꗵ|4T�T UV�7�&"ᄶC,���V�f�軤��]��ӵ����Aa��OV���W�9�ӟ��o�����YL>jGL��W!D�6|�A8&9T=��5wg9�EI�C|yI[�1#�.��x�k�7턗$\CKu��d������f�H����v�UDw�$R���<��C�P�P��w[�(�ܙ�*����E��YR�"e9�^��(��cga��cf���f?��뭳�3C@�X�As�n;&̷:��Q���0�úQ[O��4��J�T�(��)D���P?����Ï�X����Sy�1[ܠr�2X{T���-Pi	1�i����R]$A�:�Yc%�z"c� �9+�-�lR�Fu�.)�'��
�v��u��A`ް挠�|Icw��6���9[�F�Cڽ[�g�$vx�ۦ
6�k�m��@] ��m���8�	q� m�c����(�͠!C��r8����6	ׁ�!�L��q�_R�
�LI�8��ߙ'6|*j�����!���nY��<���r�"�e�n�������d����9��U��5�z��nA��.򺎔��<6Au��1)T$����"N�9�AVg���T(ıIk�
����bc[dv�3AB@x�:�V��i�9��u�}��ucth3`��G_b�l�Һ�z�|$nM� :z����7��L�EV�q���%�bb�a���!����'8k�ƀ����V���}J�C	?u� �}��	�(@G����<��"�|Ԃ0a�6���u�s��߁ju���
���6�@�$�	�Խإi4\�7n ��o��
]K��A��@���E���vuǯ��L2�;M�ߡ�	O��y��֨?���?6�.~�X�X\�B�`یWq��6G�o5nN	B��E�%�;tg���5,����E�@��ة����SJ���$PmI���\�н!UQ7�)�C���J�����R����j�c
�7���j�lZZ�o�	��M��x���~�� �RQ���`a�q��o+-����fX�e�t�U�#���
cB�3_�>F ��V�`���޶� 2�>^b�6�N�}�{�ƵD�C�Q���~>D[
g�j*�]�8�#�o=v�殫52.R�4���z���P��r,�/�n'>��Š��N��f	��f��O�b�&�+ڭ��pa�*"y���ݗ(�4���޴��r7GS��\̩%�
�.�$$���2� �sт3?،P�N�B�P��f3���N�b���۾)���R(�Z������'�g7w�:���h�6_���0\�]�S~LE�H�ѧ�����ä��s�]hȫ*[�F�x�G\ӹ��<=�:��t����32g��>?�<'���͕���+�HP/N�#��=���Ż��r��<�x���[T;��P0�0��0�а»̞��ѾVq��Ə���Dî�&�,yp�WoA�4�q*��A��jYTG]�zV"�k#���g�W���5@��^Y����w\'7�:����Ɔ��2ߝ��y�Td����i�4P��G�9������n�Q�{��KE�%p�`XxH8�
�w�a1!dp)�H\�}!���u��_��7�,�������`�kM�ʧ��<��^�s�y!�$����3�}A,2u�xE�T�O�S�]	�]Y���I��T�_o�� �K�>� _$ٔkh�H�$�'P�?�U�J}u��0z
4 �'�����,���k!�� ޚ�@Ơ�π��4�ـ1�>k��4��	�8�w��^�(��so���ML�a� {#M����6V�ɦ�"��U����@��
:��*����˅������y�6fZR/%���V#'��t�0��_� �ޢ�I�RL��j�#@ B {}$�L�K�����\L��hz�ʾB����Uf��� �d�40u�h��D���U�(�\ˏʼO�ۈ��+�J��#������لݘ�gw��D�'�Ӵ.�״6.�>��6}��`�lv	�;�/��*N{��9`�WK�C�/�pwW�߅Jwއ�V%��m-��uc�����׻�h�_��Y4��&�e)L6j��[;QO��}DU�CF�����C�����@���*��L��^���!��U�r�-n�c�� f��N��EA���0_E���:;]���L�tgG&ъzs|��G�v�篇���ǆ�e�>��@�׷�P4�P�7��QhW"�Rz�����>_�
��9��.���P���Xp������/�]�@�i�R>�-����6s����<��{�T"CG�I�G�<t�&E�sz
Ɖ�Z�J*��̀E��~ɗ���Q26��n�7��o��4���nų�s�0�-8Wd�+p���Lu@UtŮ�F�3�CZ��$9[�EQc�@}=ŖJ��¹&���1m,T�%1���o/���ȒN�Y)d�)�.�xG�iR��D� \գ�� �.s"�m/�Eګ�KR��'�2Ua�bmj�]׏#���F�3��S[� a��>QV�X����=��K&%�bd&����̚(xm谗���-g����Vf�E�a9;�k��q��'��̕�k/D����_�2�H��j�*Д%Vg������f�)�2�1y0�;��������,M;RV���/X��nYw��k�+�kV8���,hԬ�N�%>�(����b3�?�D_+�jn��/.��w��]�Ŀ���^ΰ��I���ux�!B�o-���0�"*�_�,��8��4\6@40:�9mQa��@i���W���`Q�u�#X�g��Im�m�^��z�����t�P�:��[�P=n I��&p���ʓ�s��_��J@*�����`�����B���T���'-n����X}r�E��S���?�gN�	��I������.�#���ŗ���X���'Ń��;t
i)х��@����Өqs�M2�Ú+xQ��.~$`��S��^�^sHH�S��a�����[�w�tU��2Ը�8�4ϗ�� ��_h2Y�B�Bh>�2Ka�1��ș���-�s�3��٪Yhv=�l��f�����K@ N�Z����8��7T��D�Z�lz�/ڞ͇��]Ķ�aB��F�^U���� �"	�Q���B��8z��
��1�f����ݏv�:Z��L+�j�.��� �}�iLA���^�J��N��O��	cz�g�r.%n:���!��W\TvD������ˌTb��zt 2�2p������FѰ�U��Aua5�����ϔt���	��L]^�$���¹6��i����u�_L,��I�nرT�V�o˰r���`�e�f���@*``ϱ�wU4�ޖ#��W���F�$:��Q��+z��Ũ}V�-��+u�A�dB[1�ܿ"c/mF�E�Xn��]?���>�ӏܳ#ؚ�M���E�����增i���	�3	���TjA	�PѷAtД�"���k'�:�H(q2�h�XNnV4+����\�o�^�� |3��������Jo
憮�R5�V#@� x$f�q��m	0�zUϐ�Ǻ��[t��i�L��}x!�7����+��}'`]̍k��{	�&�*�����Է}!�;2�����K	!�����!�τ�S��|��n�pr�d�Zj���Kz�)��'�'V��z�@�M`�vUL&�!k�f��^/��V$�>��t7m�$��ßL��$�c�WO�֯G⫴�LNB�~x���ȱ�41��s��:�/:C  	zpH3J�i .����p��~��"�~���0{u^���H�}>s<���R�i��K�N`E���r�?3Oyz����L0Q �֋�����#N�Q���´2y�Bwނ�����BUs�[�-(�����iFL��p=ƴ�[̹׳�3��}sĶk��z�ݜI��Ȗ��󦔢�WO����B�ݖ7�&)(%���m+� :V�{����ȍZL��vf���PϚ�Kw���/�'=2�AAK��j~�G Im$�=W�i����nG���^i9s���L��Q'�}��Φ@
?yLǎ����U�P���W��T�
���' j�]G`n<��u/�0_���'�:�#@x_���'��h���H������_���Fƈ�z��s�[�K�%��bu�p�i�	6
#ώb,TxTg??Y�Wb��&�X���,Ԝi�%&\zJ��b?��g��kF}�l��2a�m�A��5�l)��]�Nȵ"ZJ1�v͟9�(8�@Vi��s���q-{}mJ�1����Dl����:�y�5@���u@��Z2HS  �����~@J�͍H����#E�9�z���Q����3���/m�X�W�(K�ct�)��;�g�q�py�#D��N��p-�I撢�`;�m�X+-� ��c�}�d�/�<� �P�1$��b�A��
$�pS_����w�eS�n������u��� �S�k�跬��_�����I�t���4��0�Z8w6ןYD�o,?����3�};���ͧ�`�P�5q?�G,l�Ҡ�ab�1�P,��N�����1��3j�ju��p�b�o�g>9%G5	}g�'�J0RRvs�Hz�D12�O��?�Љ��h��'h��EC�����x�(�}�����{�W���7W��W)ª'C y��@x�(�&�:�!0���E%��d(P������,/�E-+�p��3���s8�B��(a���u��J����-Y��SX���it�9�[����vx`�4up�UcP/^WK�!���B'>_=�TH$�d���o�tt R������u��i��E�Ϛ���{�����dإ��΂���a�\��U�%q�q�~l���^�׳�A��F3��)/�S�!��^v�洅����S��˲e�QA4i�<7���\�Jk��\C�A��x����P�)�`��G<]�Ş��&J[2����uy��S�U��A�-�����7WxR��U��;�X;s��>Cwq�մ�-��v�����K�|�t�"> �)痃�o��fvV{�بC�4|+�qX-w^�͔N��)�i�~M�N6�f�3-�u�(�I�scڅ����J�
1��Ha��n?aw�9z/T��<1��Wg��2�hR|9���_���y�u��}�$��3g~'$
��4�|��o�&Y�T|2v��l��nh�ɡxK��T��x��9	O��Ƭ�K�.�7m|+�R����z�8�O�z,���0�.���}b9�rԓ=Ʈ����_PXgG]Q�D��>������օET�}������ğNk�4�닙!��G�
����[/�4�X���Y#0���#�^���G�tut�I���d"�g-&�'&(��;�T5S�wg;YJhn� �В;J���L��&>
q�����w8��a�~1@Qv��^��?.Z�����/Id�5!��Nä��S��ji6ɦ�%��}���_�w
�(�n.��>vrk�{��g(�ΠQ ��_�2�aE�|ՂM,�a�� �?�C�!�1�����!~�tKʴ��'{\����H�8R[?��:Se����}�����`�ћ�m��d�!��hcH��ӽ�r�}+덩�.�m��r�n�Y �bc������񶳟�W��q�؊��b ����p����l��+ L��$�ϸ�zYʀ�e��'|���~�C��������J�*.1�^!Z;�����m)�m˭EU��)���DR�U���i����I� �T7[�*�)��\�����<�W}�5�E2�F�<([;�ˡ�:�ö{b��f�@���@���U�u��iO�4~bl@r�<�b�Ӫ��7�Y_=�d���A?�}%Z�4�O����/s���7�#���T1�E^ey)l�R")��Ƨ�Y���[`1����������}jB���d�[�y��m֦z� 	hC��k�d�,z�Kϭ�@�B�f\V<���j!�@GCʼ�$�P�:H]3z����v��ƕHbK;����O���V��q�a$;����T1�Ue�Js�����ͧt�K��� ��#5���l�\�q���@���D�*��dpN�I0Y'���ѝ�.�0�j�(�O��Z�[�&L氂�Z�� ۀDY��ٽ�M�����񡅫/=�*m�'�øK982�hf]�D��˵8HF,������ 6.�A��^������fiW��F��0 �3���4&:��_:z��~�,_�W�*�	����n^͂�Ni����6����;��|�7Ps(kR��;�Ӛ�;���Z�đ�O^�KT1K�c^��΍[�bU=�{����Z�_������j�/s�w���J�;-���i�Ԭ�`|w��W=5��Mqn��2Ju���o�ۡ@`�jZ����W��ϡY��,��qs�# ��2����!:��*Q���d�iaV��3��vK�xM�v�:�l�kEa$)�Z�xӯc*n�F�*ỷz�65'��;=��̾��7�����q�cB���	��rd�G�9L;��_[��z�񎇹"�=�ӳ�Hh)�>��8��qɯ�����S9����	t����l)�*����a�G=�+D�0Ñ�/i�dp�fQ�t��}u���{8׻A�p%�(�q�6O�sF��c��f��U.pZ��&� \TɥE�D�� �fAUP֥(z��z��U2!e�1r���>�<|ƫ�P{�kA�����ckT~xZϝ����jW�U~�ц�IԿ�_w��bR2��b�/��C��U�i��<c��S�@
u�]%����_��������4�H�8o*.o,O�
�	���i�BTsF���vЮ��B��V���Z]�7,��`�d�zz��)�B6�,����HAD���QU2�����k� @?������V�G��#�O��B��[�	��:��&�M|�;mWk���U� ���=1����k��:!���G�gX[-��XH"��7�4�����>A��Y���sՄ�� L5r��+��k]�9�?���1g�������k�cO3����5��S��h?k\r�D��W2�vFk�Mnwb1�ʺk_���6����n�^�Ά�8�D�7"�0�5(Sn:�����q��6��&`�O��o�a��Z7M������z_=�/��V�b�����V5���8�Q�_M$�8�L�T3�fu���E[�P���ifo����0� ��y��`k"�i,ԡF��`�7� A�ռ�0�UC�l��8��Pr20�~�M.$h��JL�M��"Os!p�8��-�D�˘#Z��؈R�y�[h�R�"���	��iK�*r	S�+�9nl�L�g�g�zT�-%�>c�Օ%T�oo�-��<���T��bM0��|����YB����p��a~�q���� ]I�6��N����l[m����1~�'=wc���Xf��{(q��Ų	w�ژV��5
O�@9}��ćY�!�
0g���%/c��~�ΏC�צJ{�O�i��Sӛܗ���"�D��&���q8%�i�,А�Y�UW�'��Ǟ.l���C����EV0�l��J�]}X��Wm�+��u9+�*���9lpߤ�2�=V�n�I#�
�=m� c3���4��%���]�&���%�$s���+�	�E,gl"ʪn@�W[(�= ���C�M��zR��u���%=ݰ�I> �
O��V�C��w���t�Nˆ�4�O6�OԼ�1|G-YZ��*����k�@G$l� ��l�dE���&� ���	���ӈ�$�Y��iA��Ur�I�>���=�[�C�t���g��`?Ǫ��֙.�&����N�%aj��d��;�FWp�ʞzZvXF�w�2�~ի��$��I災;�E���Y��t�/j.�_��?r����k?�϶lc��N��5Aa�@82�4
�a:8�&��,���}�ۑk?�3�/���~�t�t�/bʞW�ef�Z��K�����"�ĥ�R{[y��,,�/~�u��BT%yb����o`��ǅ@�9���t�v�����̞�w����W��R�z7��Ӆ���Ԩ�Q�6/Bf�����|6�D�y�k[f�����.�~E`���f�\5ܨ���:9e��r�mP���,�r�	^�Ms󷥬�~��% �م1��w!�%O�����i�}�E8'g��y����e)�#�EW9{яl6E�V�gp����k1�C���\�6Q�O�wZ2(_��<�=G?7��I�]�����&N��Ξj��10����L+��a���]�|�_�e��3��}��z�Em6�L�<KÌS/�AQ�m�N��0ZP�=���q| @��k6��uz��*�e~l.�#���=FWJ�J#kS�����vF{��o���M?��:�1b(c�"T�(9���M	k�d� 
MZy�����=5	������g�}�}t�r-R�A��/��Wʫ~��MT���ؽ.�0�$*4�1�9$ٜ��Ί���g\Y�e�?�7�`���1o�%����~zA�V����@L��2/���{s�2�$.�9�g˺=#E��7���ևFT��'M�N�:*��/���/��L�b���B'��Ja@�7)7O��wI�>�b��s�!Kܣ�~���,N��3"f7cZH�
G&��$<V��8h��)ՐC.�2�J~��.��~�w�<���#OdD�<.�9z�58��"ӽbJ>��M�>����qev\�^����/p�?�#��nK�ݝ����WۍkC#&ĕq\��`<_k���ʹI�40�|���a�j��s��{�מ��°��ꈌ��,����H6�q)����A���9�e�H��$E��1�.F��;>���;�W�T~��L3[#;��>��몂��Fw�ckt?�LG�q��/`� ��U'�[��ˀ��V�;pQcC�tA-<�=�o����r���3�m5%��46<��AZ�˧s� f+��~���T��U��0b��]��#}���W1�w����� ��ߠ	�nL.)b)?�TƈCh=� ���8���x�	072���H\������ٷ�2�E�҂ ����ex�ֿ��2K�򲗁����b�s�Pe}�l�<ݩ����}�@�	�kI��}�c~\!���YX\"�����j����=w� ~yG�3���4����8�}�1"��+�P��o;�e3���.If��r��R���5w��zo��,6�=H8Z���AW_��OE�Vۃ�j�ȼ^ܯ���}A�f��;�}8 Kf�D/T4���;Fh�/�ͦ��ʳ����I!���Ù!�r#���:��y��ׁ0L�����N�ų0�J`�E�n"�������qE+�5���I���ـw���$3O@����� �i��E[�2��ps�U2g��rQ����ܕ���n\�1Kg'kz~�1�s�
���
�-�zV��;�|�$H�Wa��\�|�u2'�F�G&R�8ӻ~H#����5m)X�D�mU��b�ߴ9���f��� i�q��/lUeznzC؃�y:0�P>5Kc�����0N��*�ӏ4XJۢ��ۢ���&�u��1[zbU�	�`'In�XR��y�!p�:�E\���/X�x�3Y�0��Q��d���ߜɞ��a���b6��m��@^׆�8ļ ��P�4T�Nh����mdZN�˜�~�i<�C���K��'䰰~��g{l������g�$/�m���u�fi�jϬbm�iuj
f��NJ�1n1gt$.�	C(��G��!k�������$�"�	�	 ��;7�;<��K�ҹ��[Uf�o�ޞ��̹�:$�4p}��j�7�_��9I_���>�n��ԍW�F�$�3ѥݐ-�Z�J~T�qu������c�VDNjF� P}�eM�Y|m�Sa�EJ=F���5��7?���ˁG��|��������~l^�/N���R*�U֘�8���\����z;�)cbH�) ��
-
�C��sT%mTf���G��$���Wx ��/3����h��9�?��
�U36e�8��
0�yǾ�mk�q����c卅A��&���"�3]%mV^�cJT��ٴ
���R�L�nI2Ir$de��:�18��0DUkng�oZ�Սޜ�3�Zw�-ʞ��L�!�fW�*�f��0�c��>�T�sp�~�- m��Ӹ�
wi�q�>�)$��Yj(�Ȇ�ۋ���_��5�m��sz��r�:��L�M{*�c0ҁ梈
괩@C���������1G�^�n���z�J�ߑ�vg���/>R�mR���Ocd5¨��r�)]xª�r�E"Ɛ�G�au��P��R߭��-�$����h�sw�jܝx��rqs/�${�@�A�
��K���7?���
z^^N7�cO� ����E�z.F��P��:�w"������e�s���˖��>�HV��d�귒 �it�����E�������ዉ��g�U���&�Ea�0��[x ���K9���.�@r)Vء]���k�^�J�����>�켵��.(~�m���Bu�`�̀*�q%���'���qV�υ4��"��� &���z<�~݅���jn���{T�"`�kV��b�;z� ��ٕ�N��3J}�9dA�l�?w�Ԣ*E�wZAX#gP�#_�����*��Q�~H�֝���F33�Rրl�#�ss��N�������*�R�ѵP����i-��,����-�V�%��_>�W���6p�?[Ty�����#.:�y&����'�:�
p{K�.Z�ntQgp�iX��5�%�0����&a����[m��켎q�k(�Z�A��JI��!�Mk��+�TV�YtH`�B��f*]��C�-���p�̰��������D�PԷ����1�]���Lz�֡���6�b��J�
\*fI݅����  M+�����O`U�:.�̮u�i�#��h�(Q�4*�n��ϙ��gr���$�C�#ZQ�������܁0�����7vF'͝K�(��Ɛ6��Ķ3�|�����=�M��.=�f���j�ӌ7 6��y{���>�?��eJ9�I&s}|��b��B+�ӳ�=sw��a���Y�7EU�)�ਿ�#��=�}U��D��P�pi��V]�{���[[P�6�$p+��bE{
�U���o�h��{�"���{�+GH�1b����9>![�_]����&��d������څs�Q���&%w`�RC��)�+:>-Rg��@6�V��+#�}���Ƿ\8b���)`:x�4�#��� �5�Wj��?��r2����m&�.��B�~Y�o�`V���K�S�7�1PI�pb4��&U��,/�bjC��C(Ґ�|�][)�H�2f���/U�}�����և�s����i��#e��hp����(y��yG��T�d�41�I���3';^
�C�8̮�r���:�`��1�$8O�8�tm'�\߻����'�������y
,z��
􊓼�M0�Wh��7+�@[��&���Q+ �<�m���a�����^ 7�aK�o�жd��ѿ-3*AB��Z�aP�����0eɄ�/��V'�Z��yo�o�/������͵w�{���~��
�p�g�
-~qJtv�� ��: �@��?�`�	=3-;����=�f3��g9��J�
d,�v�DT�6�4�5,JO���B��\Y#���2�T#R_����ȑ��C;i$�j���2��U���;jf��6���Z�v6��r
D&(k�S�۾.������J�ǳ�'����y����������o��"�:�E-Ku��|s�����I�~Fjf� ?,?���s�x�^�= ���j[	�?���$(�׶�z�r�t���K�%�;�j'	j�5�e��\.���_���o����?��R
�]��F�jT)����g�sD-��!�<�o	�|���Ɋ�H;G��[���P���,����o�B��8�30�=��|�!-��s��Ih��d-K�M�����Yub��w��'�Sb��N4Y���/�����s9#u�Z��q�"#Π��
��`#;�!�m��.�g��AdGa�j�9��g*FD��4��ųf�E��g�l��;���l`e�o�eg�fu�.����S]=����xE<�M�	��ڿnZV,�O��_���t{�ib����"�{5��Uc�M���+�U��.xy�h�Ɔ'�d|������Y�}Nݫ���l��-�(RI�Q�"���gqs"��f�) W9�3Ć-�ğ;H�,�T�8ɾp�Klw>�{^٦\m����A�,�|b�s�〻v�d@�;雭5�(��w��V��i4�T���$��ET��ިr�[�[�����ZBɹ����$��ǳ?���Q!Q>����{�3yq�PMb]lo��L�i�� ����o�!㦠��ƿ�)&�]?�E�,����A�y�'ϣp\ �&k�1�Y./6� )����c�PZi:��a�%����n���5�=��$w5R{��g�3L�S����U��7̠���F�h�V┛	�K�|��	��5��ye�,gN����h�� �^�X�ޛل��0|GE�����}�h�65��;tݡ������]��5@�4�����Yv5�?n7�u�i��s����pD�M���$�bz��K:�̖x��6��.�<��B�Z*l��[!�=CX�ٮ�sIp
u}\�3�{�ۭS��J���J\��E���v�f��H�]?AF��&����*78� [���AHQm��\���O�+�!�'��`9�=I�2�M��WP�~��9�AG^�,�k�beǤ̝J�y�I�Au���h�F�6�C�)��ԣTd���iԁ*_֧��v�T�<��<z5�O8��Vlk9��Z�Mܱ���Oְ���Y�@$�	�����ΫIE��ip6id��%�G�,�������. \PmS�$�N���V��{^ޑ3����+NA�k��ā�T�4 \���n����kЌ��z1:�=!�bI�2��L�V$�ƿ��z:�NW�|ڲ����'�������y�$?N�������C�>qW3&���^\��d�\H���!���ٞ^�D#?��>[���\R	���J��@�?S(������Yp�y瑣e0 HZK�@�[joN(p}�z�=��~/9�3u�p0�����A�Q=��^֣�GJ��av�H��$���'v�?u	�N���q���6�
�� ����S��c�KZ����QP�����%Y.�%�
~>�^p����V�� �vI�W�2'qwH"�r����R������' ѵm��;��~']e�tw�MY{i�2
��BC��C�f����v �m��yA_~᪈M|��{��6{���Vr�9)TU���3��u����eǸ��ǩ�fa�)�g*���t�=4:Ѥ�,4ͩ�Sæȇ�E�QC��|";� ���	E��ω�?���!A��V�<�P��{�e����Ⱥi-�2������W��̕�<�����{�1��,~���/�&'��p��X��ꂕ�綴2n��D.L�$�H��$�s �=��c�[�����>!�3�xP��L��'�����('Cj��}���H�)?/�Ay��>+Ę*1�5�ğ�〴�\�5��O*�5�^���o�?e�6֖����dq�6���֝�h�"w��ǃ���צ@�%�u.�� �l�����I0,�t��e���꒾�=�M!�o9��� Gm�첡$�g��&F��s��-�Ή�L{�)!qh�ڄ\�G�c��;�3rt��.4Ч�55$��-��c :���ގ��"��XF%���zd��1����R�B����s�f��\8p[��g g����U�`�<���� �1��E�i'_�b�*�/)�3����j|!n��Q`�WYU���p���9-�r��E69G{��v�ex�k���N�,�E
}�D��Zĕ���6o��m4��o���1Qľ4�ڽ��yb �|@�׹=��n��� �A�b	���eB�n=�l��>'��|$�*��
���
�t��5��v 1X�o����c��a��u"�(�N�:��Å�
m(�Q���P��ra�;�% N�{�>s�Cc�1r���,s����803tP��3=��S�5�Y����^�N�&�1$Lw^�����D�FY�2F�����!{�5�P�ѳ�f��o�3Yaܴñ�HI��PB��M@��G+3�K���-�VU���D���H��U��tD����m`��}�gS�)mS$:} Zt�P#F*�@vA�o�rymo� ���1V�!�v�o��c2�]�Hp)J)
/�"�#}D[�ӥXo�	�4�h%<وGb����>����h��th�Ⱦ2�S�m���*�6����_���s5қ��݊]:�y�'�sߐc�ꒀ`�o�d�$�o����d�b��Ѐ���w�=WsboT�A.���I39 ��0'6@��,�OO[(���.W=����U8�.���A27r�\�؉���6���p���#5>�dS���f�ޮ�ңhK��M����p� Ce�a��N&ߧC���0�a"X�w{��,FUX��{�Y��V�WR<�͔4"^pb�nj̗<�(�U�׫�a��[TRCE�^���!��Y����[y4����b�]E�����P��B�B&��2������QW���
�ȕ9/sNu�I���	��J�T;��֡5NU�����2!��F&B~���y������2��
+�mj�w�`�w��e�-�g2���!vO�D�yT�~��.6Ԏ ٹ~[���Ͷ�WEPC~�;e�#���Mr"��N�^���(�����ǰ���b�^��8L���?t��W��!a1׈)$pA�jCE��0�M�2��_Ϙϭ�B��t�K��,������Q+%^��hǄx�-n.&�n>�;�c�����W}�)}��j��x^Rg]o`����l
H��ґN� ř}r��ֱ|��S�-8�v]��?��R����rVw�*� @�z���帶[新s0�4�<���4"�h�[��L|7���GNK0,W�4b�蔤y��З�$o�Z18.�+���!���K����*eYʹ<e=Ύ��0���߿��\���؉��m���Ӎ�d�h_�]
�@��L��̳S��`�A��&mɦ�x����#q�b4g�Z��^�3�b��(��a�����X�#��u��J��R,�@�Ќ�/2�,c���6OC~��35V7�E+oE�f>�-T%����:���&�Nj�|�Z4���: �j�Z�����ő�ޟ�EM9���YY8��@�S�d�O�p����0��d]H/O��g?5�����1�F;-��);��+�.>v���� c����{�&��]�����[���t��L�}g�'hZ��E<��J�h��ȾB��V �>|�����̈ڈ9���ܳD�-i)��q�H)����	����\J��m����<����A�'�����2#��#������$��Ǒ4��'ў�,���H����dG������3��x��­�Lfn�T��u�&����n��ݠ��2�m4-*��� L��|=��3g�%A�θ�S�תx���W��6�[�_Qg�_��.��z|FBc���m���2�j��}����8��+](C��p�DPF�Aq�8h@�X[�s2q+�:�\�7�qC�ܚq�����a<��z�:���k�&óp~�� �\:k<���Q|�����3�[#I�=Q�x�S����"���|�E�t����ɽ�I�5���b�T�v�/M�9 ʳת�jZ�N�+
���;6�[L�2��N���%��D���]�X.�E!��A	r91zd�]�fH^�z�'vX���k�L^�J�T�+2_��}z�o}4�LN����|TSJ�x�*k3���J�'y��X��)�U`�`�X�;�^�s�e(d�}��?3mh��(��:��^���,�.����ԧd�ׇU�p�������t�'�N���rR"W�T���E�I�#cM�r7�Ct�,�FB�2�@��y��q�ձ����\��iQ.��}_oF�d{W8��k��o���ưxԴ�\q ¿���"��Y�:�xj��S�Йf����x�r1Cw%]~\M˨K���t]�
���)1!�On o�b	y&Ʌ-?l��{�:�R��1V:v�d5���P�|���g�o�)*�n �u�S�#�#~a��&/��e�!�ۺ	:��\���v�o��E(�N7��Nd ��V���	��oN��zO��	���)�"X?���>ΏX�]��� �Ol�z��y�E$�z���j�0�)���?Fc`#H{�@7�vbP���J��Ҍ���ÐT�C��3b?�Iu5��N:Vxń�K���kq��(y��i�"���wHw�I�,\��˻}��l�33�	���z(�cU��j��dLn���\ˮ߃�Br�Ѻq�~y�W�U:�]^=Ȅ���-h�*�z5����O��Tt��-���z͏���yc&�
T?��%��5
�"�"v��яެ�)��C�\��{S�.y!��~75%���&�}&��9J�����iO	��r��<|Y���
�"j��y�]�ߏ𒉑j�Z�=�Z-V��>��vm�ï=Q�ؠy�.5�׋SW8������]�>�����Ws�8CjzS*Cy�6�I��^��S�"S��v��������  �'7h�/bmL��$����s ���i��c:�����MI`����<?l�ܤC�Ǭt���'�i@Ϝw�<��#�_���k��
�4?uN�bJ�T݅p=Ig��9��Ⓢ2��O��ä��G�̣��\i ���j#�]5s��+; �#�Y��R�g�ϋV�轣���(�Ok�����u�ٚ	�� ��o���~2#1� V|b%\�Dh�pT��#=�߫J����OOfj��O���MI�J�}�!ˆY��|�6	m�oC���Ң���V@��e�椂$b���|�k>n��=?U�ن�k/���6N�^`K�R���r�C�0���8��y���p�>+l\r�P��#Fm�h
�en��*JR�+�?"�ICl@��
ߤ� �%�E����[��t���ŕ�/�K��X-��ѕR��s���Δ9ḓ�kEN����w��~�\���V�t���Yl�LQ=��ෲ�اk4��, �?6?������p����W�P�:/n������1���\���)8�>|�V�8�D����T\�O����慦<�n9�:M����z�L���6�ÄSv�2D@㩉b0.5�@ ����ԙ�h����t�}�����a��)��L�E$�I~`<Z"�CG@8���Ts.��F���b�r.���S��(�c�N�3Z�"ޔ�OK[!��sz��ԫt��n��[�D ��3�s��IီutwD�j�eᅡ���h'L2���Ěv�G�ߟ_�Q�e���o"8�������()�%��RD�H��2��k�������/��}�W��߲�^׾?�,�0V
��_V$&���j�G��.c%�Z�Ҟ�Q�(���W��5cro#�|���K������=-�c/���~`�0�C��'�l��Wԭ�0�־_qݛ�D ���xk��k`̌^���rm=u���y�q>j�Û� [��iwq�y��C�*z���$�h�k��yI���ZJ~�om?����CAf��6m�5���%0<�P�&�L���T�ҍ����O�N��%��!�X�u����x��!�/цD��p�̱�A��X�<N6bM����WF�Q����d� Gq�T3Ͼ������1̃�����vȾ݁��J8������}�l���6���A)?�l�o��7Ge\�}n"����n[�&.�C n C���R9Q�wu�z�
9��ed�*���DUay��rZ[My�O��Ǧ�h��P�#���ʂ�(�>k�،ڏ�k�l&$>j�����ck��t�������d�2��^�?��G��\ �mz���!+o�iӞE�Ϡ �6�� H���Z��2���� ^�Y����F�Tc:�kE���%e��2i;l7V��놀���je��֐�q`�P�j$��vbwI5��#�A��"'3���p���.�����o�I��.D�Y�{���J�7��:=���D��n������f�+U2_�gr#�ø綋I��]2%���;�����yP��b�9`�5 ਞ�b��xʷk	��|�3x15�It/�,�����W3���VO�H7_,4qo�m9����3JD��>�JNT"��-k��d濫#El���dD�5v�xup����L<��I�:G]�=�(nrK�GEGjI�2�̓]���4K߶�]��/�z;,�(X�9���e��n��0���I/:���4G�&�5�|�� ���[�
�(���㖟�i��2�!�M��-#y�D?!]��m�iL�u%�Ӣ$#�y�g�Wo�@l�id��C��rt���4X��0�,c3c��N������U�	f��s;<׀����w 6�Y�9�e��H�1�f:p-!zt]�[�vF�V�7�(��ry	�4��{���q�)43�*�U#�����;�3Ե�b�y��O{�ϼ��y�)�*����x�=����3��huGC�j"]DGÂ�K�P����1�C�St��� B�!����]x�0%��&,�p�8B�����n��z�4{�dHC6<+(��x��ΘQ����h]0�-�$��0���ܑF��J���P��?���-��Ek��}�ԫ����u��}�Xy2���qB��b�� q��%�v3����=��-�9=��)/:�3�5៦�X�z�Ӿ�l3�gJ��>C	���!��8����?�&@xT����S��*�pR�Ǽ#���ҍ��}�|�DȂ|J�Pm��*�F���~
D�)��AA�0��s��������p9�I�7�W���=m�j�[���8��F�����zI����V��j�j�v��eh�Ĩ�q�GK�OF��j����M�������`!7Sl�W��� xk �͡�hL^Js*�� �(� B�(�*�����oaz�C�J������wr���{�$�XC�>�@i�7���3�F(��B�k�1�I��I8�_��M�^m���d�=��ݫ�P�U$]1F�	����3ꢸ��~g��kg������i/3�E[���&/C�Y�U���e��(�Ԕ:�iW��_�c�&�a tH=b��,Vi��[4��:8�*I�׾Bէ�~VQ?�~\C:8l��a�"�l <~�ůc�e�z��L������ɪ
�P{׺sL�|�����Z<��� ����if���9�s�5(G��觓��_c���Nש�hX�*�.׷^ɹG=l��; n�H��]�wf��D%}��%D���D2G��8Euh����b#��&���8�Dt�]i]��#�������>&��I]Ǹg����,Vc-�F1���Q��* �/���y̓X�z哇;/��V�usS�>����.�Y�qͯ�"5�R�D6�����.��NK��U5dȓ�~7"�]l�.͗_v����4���
m�%��@�N{��d�80�]��,��+A�há�V]%U3M��'R�F��/v~P��(�˅�2����~fO�K#��-�f��P�l���UF~��No��z9]�G(y��L���?����Z��ؕ|M�o��^F�Ϡ]��d��P�s�;��]�^�S��[g:<4�i/�B��:�R�s�H���^�VU�E�M^~�X�}�Z��}r�� F����'���_�MX�8�T�x9�����ܝ�R;񪚳��,�d��z�����J<��	���+o��S�!��A����.Gm/�|���S�MO�R(M8�����:�]���cL]�S�(d��X�ǰ'�F>#��8���d��  �উ߀�X���%����mR�%yc8v����+ʾ��w4w����h��FI"��*�޾�w��<U���_�o���ȿ�GwS����l^$�>�`4��xH���<��=T�-���%��n]|Ѩ�̙��Pc�j�:�a�:tZJ+�pǿ�yX$��6��:�T�fM������~�`Vб[�U����knL�q��Jo���yU�j�w(K:�������������x�l]!�p���(������/�.ؠ��(Y9�t?'�-�ɫD�Ы���]#xקU�{T��.|b�.�J��5��q|�&0Qr$��=��.CӻǲCι IM���L��������uh�����`1�KO�"��MQ��N�������{�#x��/Q�����3��| �x�!���\�e~�
@{����7�X+	��Lo3a�B|�C���w�,xyx�:��X�2	�.w�Q4���a��K|�0Dk��܀ð"�F��2�8��6�f�]y�3���0��	F�=^���Zٸ��y����bq���Pʍ%ep���wT���m?�@�C,&M��w�/�����Y�]��)*���ee�c����.WF�$�3�uN����l�����&SV��ۈI�6>�2Bઋǐ2h�"5߀�͈)6�q_M7�#覼K�}���S�~�͎P����n�����L}�)�R+e9�_f�J��F/y�oJQp�k�x�)2�z��Д �w�I��>�b%S箻3��"ES��^��3V���Y�>޼�j夵ޏ�x�U>A2;8h���Km���+�d�)2y�S�+����Ґ_�y�L���Z�8�4���X��5���k��(;�@����SM�O9�>�x^k��0(�7>�+,?�-	"��#C�\�EM֥����q�x3{�S���p�)ev��Ҝ.��P�=y)����ɨ�*�?QP[hs�Wm�����h*���J�y�^�N�?�J�PR�����@UK�_3�b�(K˧��r�B������Q�^�_��m~��_�[�## +;�A�|!Y�PȠ��w��������c�i��ǀ�z{�Mt"�B�&�U��>̭���:Y�mg�p��#ګ46<]�1$�:d&S�������L�<F;p�"�Q�cl����9���gFY����v��:[� ^�Z4B<Rc�l��=jnVfP��?��h\�5��F����A-����9Y�yGK����ԼW~$�J�˚S2r��U5&�����ǌ�q ���@*��Ld� ����,T�&Mv���՘�}�7H�x98nYm�0�UZ/w���EQ�����g�~vBV�nǇ�&�	����|{�*�g+��'U6ʶ���&3����+�7'��_��2H�Bo<��)���O�.�ʵ��o��J��W��:�i�h��8��'�b_n�N�YZ��o�I���˔�[��d���O��1r�Xq�ai[�{6�c�Q�>���{�h�H��?2�`B)c?R1�8_����׾�"(b,���w�ڸ��y�U��4���������!ᩋ���!/�)@� �d����b[/�(�ثU��������i� ��ƢU|1p1�а�SX&����T�R���-��ŀee*Re�6 �Te}O�PKC���ƅ�lD[��%�P��<u���(�$�b���K\_�@Ie)י�а�d��������Ҭ7������X���2���h}��ُ8D��J��a?��:T-�ǽ�B���yl��Оī7n��^�A��/�ߐ����?�q��&3��k�_�|֜ɁZ(5�DAZ���YP*�Ɏ� �ݥ��"ՕPl��#�_�Zt�5�=:cNy6.�s��	�8�:�N�O���IB���>��wv����*�W��"T���NH�442�R�N|z��&'Fw&�?2M�I���{r�E��,V�{�>����3G�F?:����b5_?0�٘������ĝ7Ѥĳ�Q�H�:�F�o���u����4�B��(�k�c��������m{���h���;�ƨ��/U$f8��X�n_���¬ĵ��/���hWw5`�<��_s N/ �i)dG� �_�p��l�/��}\; Bbr?�/�9�գ�=�pj��.	�n��io�A#�Dڞ�ln��Oo��L�P�Tu��#��<WO���s�H�H����_��!=��zM���I��q�u~�
x	���y��P4��]x,V X��5�[�����~���ߍ���;B�>�ߔ��5�"2M)�4:�3S�k# ��������P��#�PW͙��Z�
^�ij��P�yT��A�K7��>cwh�� ��/}�l/4`|9"�4:���o�U�c��fde2��G+|�X���Of��o ��ۤ:�]?m�R�Z�Q�B�oѭ���ڷ��M��|zp��~y�� W���O˒��=�.��W��v�Ϛ�y	ڛ����J:�
��T=��k���_G�~�цײYw�����F������:H�/��Sc~L9���>��C!�6ӭ� ��k�[�4������m��đ��?_�`dڪ�%���Q���������/$S�����ĉSe��d˾h4NIvv�J���m^��x~;X �� ���hC0N�{9t3A\l��U��_s4(�P�MLytAg�Jq,ص����d�"��#c`�������(�t$�_��6We�I�|�Ͻּ����3���2�����f~�� 3�Ì�R�o��B/I;�����������*A�w�d��d�{*��q��kjj6��ud�YR,p�ΔQ�'��,%�ꕂo��q�@��>��wG�0�I�S��	J@�.+*���>���i���(Ͱ�>wM7[�{��'��&ZzN|�0Z7����ɰ�m4ˬR:cH�5.l�Y3��Ey������тD��Ƭ�F"���Y�������)_N������jO�cI����=l�{��*�<�ϛ��֧�M8d�)�g������rW[�s��������#j�}M�%y-ݷ{��Y<�͖�ڰ�{;pU�+R�$9WQ^��Y.�A+c�N���g�A�V#�^Q�to�E�����v�������.Z?7�xZz/��wh]m�o8/?ud��A�����
3?��A�ضx���0�5�}�mj��dumI�0����%�J�
�tO5�󺫋m	K�/����������O��l�(����0 XH%H���}��oņ���Zi�ǆ��tH�q��}�1���l���EGһ,�A]|�e��U�l=���ac�B7I�/��6�˵��YOǠ�9�I�g�'T�q����ڠ�!���?{�˶��Is��)����
J'����,E6���Em�
bJ[a^]Ys�nT�L^(#�	�M\pPq�Pf�Y��?�^�� {���xl��M!��_w����aԶ/�{-H�iR���r��i�n�ίb� N8ȵ��J�U9*�q[�a�����K����L�ߢf)1w0�����{�%M�@
*�vCEO��E�P�z]�9/��k�2s�ŭk��!��)?¿�Amx߆Lg�8TQ�@S��V��!

J
gS>G�>]�b�[��7���^��ڢ�`�]�3�A�7ѿ뿜JH��_mZbf�����:�ۘ��u~Wc����엺��X~�ز���j�̵���{>f�{Y'p\�������_�Rݣ�����	���y�H'�iأ�I� ��H�N
�;:��X� ������cåB5J��s�@�:�v�F�0f{�{�܉�Z#��,���"(�2|����K��8��(*�,����_��>4{�J˳/߀Ƹ��H뼃3y����q����-�;�Jz/��c��x1�~-CGi$�3	׵V�a���2��D΃�[/�>%- ����ǲd0�c���1E{�H������c�mDָX[��v?��:�`��C>�G��"��/�]�厎sň\gH�5�+��`�����L7����JR�3;3�����͟��^��OI���(
�w1�Z�eٷ�`���yH���R-U#��w���yV~Q�e�p����5�\��3��rߡ��x)�y$�B���{'ȝ�Qb��J���l���C !R��=U��K��PO�u0]�+Oh�����ͺ:Hf?b%�4HD7�Oy�a5�ت�(M*ܷ�z�c&�u�wU��]^�7Y|��hm��EB��G0/o;�,b0Q*��|����a�-@>��M�k��wa��'�u{��[��@7dI��|�_��o��аݶ�ʢ�a�M��qֲh/�o�d�6ς�|?���~vǜo ������L�N�R��Y���*�ײ���E�����֭��!�M��xp���o��}��,uEH�̦�Z!-��*�,�Ϋf�w�CE\��^A5>�Ƴ�_O2v#m4����j?l���{e|�*���g.f�u��	B�+hUJ��0wS(ڋ�� \T�z�M=o�W�"ً���l��4�BSː�\-T��R�֢�h�?�^���0L��k�9�?�L��2��+͂�<\��I���#;P]��]j-1����H�M�HH
-���`�N�wyȮ��ޛ8Te�y�.�
��^Xę��2�i��z�m�M�~��G�$����S�{^�%̓�R`�}
q�0��s	<�����\i��όx��'����O0]L+;sHU��Ϛ�mu�{fTf1�F���B�Mz��B��i�@.Ja�of?V bXgH��[\S�²����w�A.l��RHl�ݔ�<�a5 ��̥.����S�x��8<�>�	����DPˎ��}��N |��wd��5f�wy<���H6	��:��Рe���0��7{a�1�,�lN�n"��Z��x�%�CCRwN����{(�p	���f1�yH�WA��K?��\��\aŏP��n�U�v�O���˥j$ͣ��6�(�*?)˥��q�a��������N�F(�E��*1�P$/�Lﲐ��]�ޱ��%�mgT���v��3�t�ْ�Y0��l=]��" d����N��+jW0��.V�o�V���rߖ��v7��Z"�ρl�^v.�@����W���vH��^qH^SU��"y��{�����s��As,5��R]�|X~ͻ����d�4�\:�$�����$�|�<���Q���r�v�p���z��x�r���M������� �6UD���������1��z��81�K����Q%���_���"�����K��E���"�ӈ��L��&�uL6�Ж@�r����Y}~∈e�����*BX.�Ih� vGٴ���1{~��C����pF˵��,��`//�2�:zVk�Ĳ�'+}��訴�
Π=]�2\�n�a/�\�s5A��1�Q~�#!�S�*ϵpg�8 �t���������U��[��k5��#Y��+���D�n���
�t��*��vG_׋P��f3��j����k��{��BL��ڞ��d!H����A6�[8ew�������zŚ�J�#p��7W	
<>�!��r�QVc�6�كkS7�ťfδ��{Rh���t6R�#�!�-7��4�⻚�M�����Z�,�&�����x��!~�G�
�Vp��� ����R(���M��-y��{�m������6*��8�G��Q8\�O����t��0�3	D���s��c9�oc�ġ���Z����$#}�a˪b��a��a4�?8��eGc(,�� DJ�WE���Y6֎}�3��	��U��g�K������I�	NB�6j�H)�iYb3�j?��J��˫�9x��d�N�&�9@Ϟ�LsĀ�,���ւ�E�/�odB�ۢ��םB`��1��y�TbS?�?�F͗:Q]_L��O�H�گ�	H��0������ ��=-Q )���-5qU�/���hK:X$�>�1f�������.�?��A�e Tί�wA��#��������D?����"��Pp�։�MdJ�ϕ'��_ޛYV�������oo=ʺ�8�8�U��mu�6ҽ���烾�9'�G/��}_o��C�/�qX���Ue�H��_8h|e�f��]��HF�@�]�f\h��aԑ�n��<����`'{��0�+]��u���ݡ)��g =������Ʀ&ýF�er�UPUy���JKݹ���$x���m*�X����ӂ�y�_�G�OҼ�{��R���l~�ZI�\��#�1� GJ���\�>���=�n���� �n.=N���i�^�L9��h+��'�B��#w�0Cy3��s=aG*��|m%6|�"!(�O�& �K�bXTa
?��;�z/kC�@�'�p}/�i�_<�C�	�oL����.��*�d�U�OJE������6�e�g\�d��)����B�
_n�%���4H�2�����aٱ}i�si#n":c�^��0?���g���}{�g��K[�7�o�+8fiii\F!���\�c��:�A�0������$!�����#�$�O��3;z��U&<��e��g�?8��Cv�}� ��m	]3r��Llå�_��KN$U��h�[�R�@0<�u{�A�e��ڴ�f������y����I��U�<�_>��q�w�YwM�f�&�q�·�/d�!I�tK�b�hJ;�
���a/�; "�d���^�� �0��I�E==x��!V����p��S_�;��H�ǥEF������|:Vu��;�3P��|��x�q^9=�����#��o>�g��!�t~��=:�*���a��-B��.vFäF��*���Q7 �O����mQx!:B��,�l���>�@�³�"���'�!�?�.MP�`�lۋLJwF�p��}��G��ǑW�8d\~��ְ��"�ni����C�\��4<��K��}����qt�N�!x��5P��G\ǘ�;�5ȍ �3�;�ȑK���芘g���z�,�(ʳo3TZ�J��oE�t5�atr��:0�;C4���ƽ��:��)IL~�1�`nbo�[|��0?��M�b3(��y*?�;V�}���.��4�Q�Y�}�`U&�z��,��Zs���(�3B�OEO�w~�F��/$�������/�9�m�N�ơ�j4�˥y��͟���`�X�4v'�HFv���O�Rl)Ѿ�^����ԁ�~�7�2��î0�L�˾�K(��]D5+��P��Ρzr�4�Ũ���m�V"d������K&�9� ��n����� ~*G�f2��i�u@'�@�6,�	r����g��[�wi+_+�rx�Y���G^E"#��%��}��|�J 痧e�0<�ͻ�aU��;��χ�K�h^0�{Q��"[>���C���>�C��
��F�l�[/��re�*��蜧��6kl�~�BR%-���~�pI��%3���z�]��
 ���'i@�9S~5�񾽭+��iN�垶��[L: 5��U�;�0��fR���twGd���rM�Xժ�H�C�=Z4u�0!�@�"Ԙ�'��M�ZrI{�W7��go�����l���/��G��~缌XM]����<C ǂ�s�� ����&����%�c0'�G�b�~��k}���됿wڰ�m��y,��{Ƈ�f�O��/=�Ԕ�s�I�!k�k��|J��eK���f4�@ȅ��[~�"W�(���u�vdx�6���Y�>��rlkr`��{�`�PFl����vm�h�=Dbu��n�|�g<�lUF�?�.h��㓢��X���(YY8k��x������JZ8&&�o	���N�9g�*�9�&A��w���-��uم��a��f����=Q�k`��	��xW�T~�3O&��nOi���t
-br�t��2����뵫��0Wb�w���abq񶫣"PMU�SOv@�:z�;1���ϼ��Z��J�Fxa26kdK�rWe)��c��׍k�2� �k6�ܬw�/Q��|�k|/���k����~����^��I��F՜k�����.���gH繂��Q6�;�R����.#�X�9��&1��l�/Ԣ���>H4r�O�p޳|�[�ą�O��³���4�G43ƪ��/��T�:阂��H�%S6%X�Ծg������HĄ��ucm�ם�|^��l;9���N{�nT�}5edmͱ�o��๤�;�ᆳ��C�:���Vb�S���ʊ��d�K�f/�#2��XuP�c쪜��7ą�<O���޾G�$���(���Ο��d ;�|��v`hҊUh:�>t���-�*n�	�1x!�̆�xv?h�����N��	/x�P[��l��e��r�ק���;���,Rl-y�>���c����%猍�"���}U\#�
��`k�l�9��g�o �5���[���Kr5�� �h�R�yc�L=���6��mǡ(L���Yt��);dU_;ۨ�X�8c&FK�It *�R���ޮ��h�%Z�(
�z��� ���O�ҵ����E��5��%����<"��������V5���+�y
`0�ⲵA�80�JR8�~��C�~`�.�w7?`��.�Rf.i����dY��#/j�EN�S�l���^�#���|�����-��u��*Y��d��V�F���h�p=�K-��6-w��A�c����(Ͱn�� ����oF��n̓"5�"MXb��a�=��#Y*,�DU)����̿�� :��{�� �Fc���:B|Z
T�~u�	�f�SG{ZZ�_2u�*^��Gΰ#�PQZ^����x�^�����f+��w�hv4]"`��u��tᖧ���.F���`��%��d���Z�$����"	ps`����tSXQ늖;�V}�7�Ę	{�m��N4�TM��A*�+��EnEGV��^,n-D���X�8�;��)�ܰ��n���iȳ� `�����(�֩�yw�Zr�[�|.\��~���˪����oM�H=	�EC��z���o�2��8Էx���A�(��b�m?� �fb�wG�j���������{K�+O������z�2<2BhjnQϞ����ip}3���g���@�n��C��-��D��%c�;]v�y�K��e�,�8A2e�y�#X��j�B]w��o�ϴj#P w`�d,�j��V�(�2���5�Sz�SK�<�3��3]�a�u�;�[{��[� T�8 N���f�>�޲�3�/�"�V��I7��E�i�.�pj�u 9�6���m7��P�X�䷀T�>ǝ=i���ƈ'1��2�z��u<"�*���&f�S�޷�|�wo�0^%�y
g�Ff֧��͖�����`V"��v�m�����B�f�$����;����jW	%r|��O�+�APЗr�U���9&_�n���'�7�5+3��`	a�N��9 �̵c��U*e�b�v���P5�Eb���i*�w6��ny�D��R�JH�z��傽���Ox��f�y���?��	�xn`���B�4D�(dgA%1��
�Z��s��N�����Y����g��d>�3D2��3[��5�چ|g����ZjK��o�|_��ǥ+���1�� ��C,}�����伥����Gմބ��Ők��H�ƖVLe��bi��Q IX��&)�&���;>�G��1���wSԚl�7���:�C^9�����F��J�}p�,�,��4�hHy�!y�mg��k��6P��SH,!����o�;� ���&�[���4	mF�bȁ}�o��(�1s�W��>�w�]1��3���\�Z�b��=���m�ʖ�E�QpX�����NP��IǕ�R����S�YF��KJ�ų`�kc<��)��ڊ�&21�A��t篣�9���,�u�u4a��ZEAr�D��%���fr���"[���t��	��?j���zdB^�nKK��Wu'd�9@o���|J�,%��bZ.��
R�'��:�蒶Z���*�?�l1�n���cr�OY� ��2�y�E��͇�b��pi�;i<o���K&�*��[����a rImf�$�f����2R��2E9�L������|i�t����o���ޟ��n�=B�3%Ɨ��0v	*�7��X�t��!������K0��I�X���@:݄�����@���ܳ�6�<w~�~9����B)�� �����9&N�m���6�S��m_��A�<R`@!�+dt����;GҬ��p�X|��%��M�az}�����\�46^'�7������HD�\����i��f��/��^{Vu��7���s4���\�d����$T����&l�9-{���z�z�gĩ���vO��8�v�Dl���7 �[i�]Lv��d��\�j�
��_Z��8d���Ė�1��m+��p�w���q6'?_Ο��^�&�ˎؕ�al)�D�^B�!N*}�=�%i���2B}Ǿa��ȮB��7g !�򮦫�h�8�P�#_�.���Q��te^���&�;�����o����QxVJL0��mm���:İo����駳�yn�r��p)����>��^'9E{������{�]PR7"�cc���xcy4��f�)~��B~�K��ݏ�>7�	~ȉ2�͸ӓn�q����S��4m4w
��h�Y�Ft��� =��H�G�4�wj؝_X�#Z�i�b�E�T&�0��Z��ST�C1�d�s���$&���ёYQe��bؼIx~`��h�;:�-h�x����}q�DT������2�EP}�햎E ��[i�'H�Mp�	Y(Q9�Jc��4�)��u�����X�tF�au�KHl�R{��[�P�|��0.!�waՎÎ�Cyp���K!F��ސ]0�i�����,I�
%�4O��V6A��t0�γ����l�۾�6���Ю�vQh�Z�?��7%=R��9��P8
���(:�<�s�8�N��پH�M���f}"?�-B�@zŽ���,�.[�WxbGхE�S��Qi��]6��m(B���I��v��S�|'}I2�3�.��N���������#��)�<>�J��t!ɷ3�C���{�40"s�JF�Oњd�X�޿g��*�ѽC��VVnOY��C�4q�f^'yeQ����*g���B5�ww�C�wy���+�N�є,�g% G5>�#��1%���%��mY4�T�ؤA���b����8{�z��P��A���L�J�
�q2�[�lP��7���J� �:8���@�A��H����!ˎ�a���G��ٛaK� 룞��R;���A�]�0կ��}0��a����x	�5����X�j��GG�ނk�[ۯ@�_S�)��:��.���D݄;���E"WK���B�YA	|B\@�R ܉=�ͳ	9��L:j��s��;���Ж���-:�C_*߰�&Q������ȲDF4�[����B9�䰑��ܦꞎv��+q����'ב�°~��\;Z���3��ٹ����Bo��,9� �����F���4x�}�m��WV*~�u��e|Tt�G���2�,(��&ҷ�&>�
�DW������N9q��i���҈K
RF�;�y$ȯ@_M]�-�e���^�q�h���X����R��R�TEe(Wl�z�Z�OϤ�oS!�����%jAg5�U4ښ�_I��5A���a���K�ci'����;�y��$�Ye	��T�q����K~�]�\=q�\�|@�����qV�,^`T��@2Iqeg��1����f�i^��~�D� ď3�bq�bU-\�^�k2�FtHE�7�\��	�tZ�x�i�yƸ�vZO�2Z�U.����N��a�I�������� ����*7 )���\��:>d`�-l!U]]��q?f�DjC��c�GT�ܫx���7g��4�TpC� ��m=E�����r�$�[O���n�3Qvz�zB�)��ԟ4�
�԰x��?[i=�H��{AI�ةvĔ���g-6r>�S{�jq�V�E�("4���sm5�>6C��~c>��7e�b�)���D�*�ʿH��27���EԉUD�?�:4�Ŕ����l�pM��3sՇV���t�U�t�8��]	�/�~�%��r-'%	�r�߹�u����1?��$n������2������ɗ�k��Fd
��Z�Tx+يh]�1�Φ��%��l�����zd�������ynFM
�$���*^�#��M �t=�,���ј�=�un<����1��W�-�G�e<rM����c��@����V��!�z�E�:�*K�xi�����bC�Hm��yS����9D�޾��Y��V�y��\	�| '
���A���T}��� CI$ f� RDkx�u�|^!u���`�����j����<$sc7�\�7����ˤi���`^4�r�!����V�t�v8��v��AyS��m��,>��vx9p�5�ݬ��b�ǫ��%9�s��ޭl�;��<�Ô�v��!g1tw��+��b��Q��.����x�e��3�#<���C��������E�~�FM�(�a������5֚[�A�'pn!���5x�>�3~3�6�D�ܘ�C���+3�\E�/+�����,x��λ�Z���[U���P-ѕ�s3Nǟ�!	�j��#I)iV�(�Ay��-:`\ˮ��%�����m�mL`n��?�g솈��͝Ͽ�˘b3���Ǽ�7����0���N���4Y�:�Zv�5�A1g{+�+����m�蘸n�tG���/�q�'<�#�|md�L!�y�F?����q!�� �*��3g3[��j�|���6ml(G�w��0�6��L����DT�ϋz<˨K|>��_?��ܙ�W~[0�j#y�b��6&�f+Z�����)h1�?Q�	���������#�\*I�8Vm��x)���$�գ�8��bo�-> �U�C��oǐ;�e�`݇��iG�[ymmw�?'~i�@��;�}����wP��hL��W�������O���~�?������I���'���WN�d�i�*T�-JnL=�����v�>|3�=j+=�����z��/B�.��%Dȥ5�;�@��W�b�A�������Lޞq�R�W�x����HJ�� �y���r�/����/�89����k�������/��Ъ��s>�.0����ܐ��
\+��t���C�;�q������m���1O@�f� ���h\F�ѥY�`���iX��8¢A��V|U��eѡd}�vv�.9�������*c3Lya��Y���	��ݎ���$ ��H߂Ç���}&�0E��vF�}�(�	�v�(��	�|[JxK?��EQK�Z_��e������m8�z�	�B� ���5t�������HX�� Ʋ�`�+��:;��S�-�ݝ+F;�R8)w��*=$�~�
\O��&�gl�d�t�s�^ʚON�B=���W�.B��d:+qs;��=C��=c9�� �r�[o�NW�(~�����w?Dp��z-�+����4��g/�.���Ae��N��3BX�[�89]�C��SM��ǎK�/ �5/7�L:�b���͖z��f�����Lg��Rf>�zÍ�� %E�I1⣅����	�G5�g���)�P{vu�­�KEd��#��E���˧�ٳ��X�ͤ��W���^��0%qfֈ���uC �N�!�3S�h�n�sO�+�����灅:���8KCtG�o՞Q�����ϘN�'��{(���U"Z�#ʜ �v{��h�m�Ac��`�Lo&�{� 6�8!M4�q����i<��џ"&����A�7��ѺA�J9r�������xz���Y����v���z�
�?��;ÇL�	`�_ �;7�[c����+��8R�C4.W�� +6vLZ�2�M�s�j��C9<;�~R%yo����~.Z���,�Tf���y�w�'H^u���ur���5�m{��Ղ� u��(<%��u�k�[�������L�����;�F+��4n�R'��l7x��uзg;+F���s�bs�+��ug\m�a�hmK�̢�Gq��U5S2.t�nJ�R������4��1x�H2V��e�o������<��D��e����f"r��:�����9�l�>��ꆧ9��?É�żE�b�������/(6a4=Zh$��a|B#�w�bH+V��xM��*ur���DbJ+QB��x��9\E�}bC���.��9�&b8M��r�I���.���j����z�����v6��M4/������-���^�������_�f�3*��� �����%�>���#�.�2��ra�f�&67�����|�p�TQ�*�����݀ӴH`�y�|����^��**�\��*�y�CW�������R6A�鯩��3֘�c���y���U����c�ֺ���w�"��yՎ5��[h�ݹO9�P���41�1�cÖ��&8rY�7 �����
�h���_P0m�*k��,����[�֫�B��'��l���8	}��gY�ь8G��K���3A��X���@��� y�n���m1�� Ս���E��>̭�����Ȫ=��:�B�Ū�I���A�$,~�q��SR������p�
O�/7g��TP��?U��˝�	+�6�����Ex�d
�WD��'V�;�[��¹Q�z�zb���K�Z�����5�E7���p*���j��W� �Ӯ*��+~i�1��ƣZ����0A2F�^AP��32��I����cm2�!P��Y:��@͛�v�U�f`��z5J�{8XJtb(�G���߮���/���/6S6�?;7Ya�u��3�]���&����N�#j�S��u��l��U�0D�p��O���7�A�q�6S��ĺ=	vG9�@�CRC;���Kxjwg���8s�9,<��7{��{9�E���;82���g�$_GΥ5�l'P%5��R�G^�0_���)?c��ƽ�!��v�%���<=�� l7��q��4�@}���u�:p�c�6����c5]��&yթ�D⌟;Vp�Y��4������5a����%vgHN�`tH�G��-�6Ure�e��{FQH>H�BP�D�M��3�"�Ѵ�zW��C�<"}Ӗ��rV���n+�^E��� l#c�nr��@����n�r����9%bjO��}`䙺��W��+w�V� ��	 9	?����'_	��8��[x�tJ�]a(p_�<�l��`ց��vsx��<F����n���c�����E����Fx�S[:������"vpY��k��vjw��7��z�(?e)ɥ�������ڴ��� �w�@��pV�
^P��k]��n��2�6�
�)�\�i4����F���u��qZ}EZ�Cnƽ�Mg��$��f:��xVN�W3��晔�n!C��O��1 ��l�����^7s}�������.dZ��z�ҍ��E2����=�� b�=���� ��@a1Ӑ��q��{rF7�	����j3�HF����J%s��{劯=�ci`~ԏ��q�nW1�m�L�* �G*Ba; ��Z�ꏝ�xN(��a�Rva�+.qV�i�7�X����s%���i	��tY�BL�O@\Hi�F)���L�iqk�O��ݰ{���P��QǧoTL*{��ֹ��s �!��1n1��[��HJ %��u����3v��'>��.���"&vO&��u/��>],__d���������\:_F���ջ�k{�"��7ȟ&e?u�J7�I7؋W�b��xM�Y1�j��!�n�Yl@��o׸wRw+>�����o��\\WI��ҍ!Ph�4&g��d��(��n�A��| <w�_ϋG�5a�t��HP��-���Xi�Kb�ʼa�mȢe��.EY)��N�ᰰ6�2�c�������v�s�,\3?���'����>���t�S�0��?}��>�٢������B��V�T;����V�r�}aQ>��+;7�w�B����s��k��/�2S��s�ԗrB�:�k�q+3�>�r����ay_��ο�aq�o�S����=�D���RY ͋���랶�-��
��]�=�ϤK�u���CS_�����`�S�s�Ċ��P�a�sK����P�k����3؋dX͜;�]3��Qj�[(=��9S;�e،v	�Iu Oӵu�����лk.l8���d��8Q����wFy�1)�I�8p̆� z���[�H�G��/�	����hd��]!U�X�(����;*�mW7:��R4�WL���3�qZ�h�iL��Idע���ou�m�����d�)_�%$v�P$G�K��
趔%�*1�n�
[E-C��4��J�����I�.��x��V��:�N�\b(�y̏�Б���=���*���4Y��ߥHÙ4���ƦUI�6��4v�%���k_���Y�?5|�9��z�0��5]��̵�����\w�ST�Q�IZ�W���i�����/d����{���A�K���ä����y��C�k ����}��ނ�R���C�#�`L�#��w%��Z�Ҽ~qw��E]�DТ�`"W�
�7�\�:rE���l��:P`´Dڪ�	�U��`uj�
4��"���89��[,��_A������/� �wr��{�ǂ����x��a��Z���p�n{����|&�v.��~SY�#�D�}`҇|���Da�^z�ё( s]R~�W{�I^�f�����N"�<͉��[��74�u����K��9i�����b��zw��������}l2a
�q��^�f|j�o+�aљ/�d~�=D���Τڀ}�mo�}�f�>����m���o�Zݻ��W	���$َ6�D�P
���Hq:��o�I�����&���)1Iye�!m��w��2���Z��5��mi6p�5�jj+G��|>  �7��N�w~����~C�WPSBU�q�S|P�1�Xrŷ�����7�~嚐�H��6�
xV��5�F�3��R�/�7Tc�b���9дU�_���
)��lHv%"�0�=��'W͕�Z@�J��p��w�e5VK��,6r�(�׏��6{���1��Iwr�C��N�Ǜ��xg�O;�{[`�ގ�;30b������c�wQ�p���AL�����F�x��n��'j ��:8����`6{%��wt��b?cp��G�w��Y�0�M���Vd_���I�J�z-�Řs�H�mX�8��u��"b�Y+d���Y̺�%E�̟D�]�4R�Q���?X�XP��4q[��j��ad��(&m�Vj�R>�S}�?���l��l�����I-���ٍ��ї�U���H�����R9&��3:ph�w�Ǻ9��5�W?��rT��`�iТ��m
"eeж.Z�2F�h�N�jp0�	`Zѥ�~O��^����#h3�	w�c�pmDR"���w�h��b��g��!�U�Ȳ�=���G�^DίF~�����co�,;�_q����t۝��?�!c�X�򚭍}����I��
$wi	��$��荔�yj���
�s�����U�����`���o0!�6�pˆA���+
�߂�'*��;��{����c����o.��|������(�*����'���Ii2Ԧxm�X���5���7�'OP�7�Pk�1�����dD$=�g�S�h՟��ᝊ���v�7m�Mb��n��SZ��E��v=D�B )ό&y"�W�~7TsjF[0D:� �K������t7A1Cs�0�Ix3S��ɾ�E��u?�Y}��no[��qz1Ȝ�-�
+�5Ft�����^��7�5��(�j7�O١Z��#�B��M��;�qT�LvcK�.k0�x\�7`o��Qm��,����R�_��5)�(ϵ�@�Ƞ��ڛ�z���n�%3���%���X��B���CD��%��G�'�2�/䥭��r�wi��!7��h��{����[g?�����ߌ�)4�~k�ɱx͡���#� �B��m�VĦ�u���������Úĺz7w@Ԝ(���K��Z3��#"7:�i斤߉�qu21�.�5�qL��se��5~Ж0	f�EE���{b��P�ό�E�*%A?��l�M H�դ���u���cBYغƂ6fge�ēS����ٸ�D��L,��/$��`[R�a=\��r�s�d����(�q��#3aS�	>z�'����;9�u��+�v��M	�\��;����T믬��vj�؃�c`:��~)m,���ߪD��VW�^=uਡ�@�ӂ�}���Ӱ`	9F��u:o�T����p5��2�.XN�%hոׇ���2u+�[��66W��ȁ��ۛQ��'���v`�F�O���m��Rk}��w%�9�֘�d���nt5�W����/�FDp~d����yh_��V��K�	a����|T���G��F����0��Q{HC_����m���4�_�du�4��(���۵�p�|[�ފN�)_�@�ۃ��g��������L�!�g���Ȧw�7�E�/��z��?ηJ���6k��O�"��g���z�Ou��V�� B��'G�(�
5�<�<$V{Ϸ�~i�����Ek�Q~^($�@�M��9A�s������WXi{m��F�P���#��c�X���Xs�|+^���N-~<y�Δ���H����<7p������3̴��_,Ȑ�D)#�{�����_)��zt��\��܅+��yg="��Z��6����6�FO(��
y҆y��@��w��
xͅ�뀾U�qV�Ͳg���FS�5P�`������.���x�W����*� )�$��	D3��d:t�8lktrN+X�L����K��^� |�x)8JoT6K}w_Q3x`�� u�u����J���QKп��=������g��-þ؎���Q�t�z���[�c�z$/,;qΑe~�9
��������L.`�9�j��c׹@W�xr�q]��{�&��D>F�ST�5T���
�����@�As*�/)p)m�@���tU%8�r͑R�������Dx�T�<ߧ��`cq��ߥ��m9;��c���87@¨��0י� vn��>�}�͛k~�u�Ha��<��[9 +t��d%�f�o
�>���j_��0���X�-��}'�#e@Ez�sl#rC��^I~�ђ�T7l[A��lGƯ^����c���r�$>��'�n�љ��&JI�OGn�˝���r�7�,_�����IL�u�O�;��]cac�EQ�I3Jab��b�>�\1|E�2=u�j_���W�����9��n!'�#ޅ��������Ã���9�9 uY.ռe�|��C������5+C�q��0��m~�-�N�]�Z�+w�K���|�Ԑ�S�ݼp�˫o$ГLg�0�$�H��r�
����=�:r�����od����
���U���&�D�f�M)�%&:v�ʫ[
�]R��m@l��jl�J�� ���%{*�4�}wݐ1��*�`�F��x�艙��=��e,1z&�"����:m�t콳�]� nz�ׯ�M�:����Y�!�$��L��&��wHo�Q�}a�j:n�Y!x�p\q��1�
�i�I���ij�`�T���;�i���N�YË�����?��m�����0�a2�:�����tY�����/jU��)#�^����ȠҌ{��ţ��i
؀�KQ<G�����Q�;��\��w� �=4�o\�y���_��a�n�]<ξW��M���WVƎ�͇�,K+�k�zk�^��|0O�Q<�I�]Z[hdD__zt���EZH��-�i�?S�yz/����� pJDt�ڨSC�r���ahl��5|h����aP�|����T�JF�ޥ�I_Xue���D�rMW�x��F�1��#j,��QHdp��3m:�ܔװ"P�2��}�mp``�	�<��|�ܧq�X����V�W%��	���k�`c��r��/c�>r�����Ұ�}t��
���%���呼��6S��EYWR����s�p5!Z�Q�Ђ.zIh<{�ѳ<��rq��AF8�i@m������)�&��]ƅ�]��Ǆ|j,��͸[P�C�̣=��Ɓso~1�=l(�^�]x�~g�y;)�R���7�8_��-BG0��[[ck	�z�"Y�B��Ty5�d��o6��_�Y���f���!�`*�{��9Qr��ɳ������s)�B���*X�"�ԸV�P��C�|Nc�9��4ʗ��H�F�~�O���F:HX��@�^ϙdX4	0P��b����.�.hk�*��k5cE��^wg:�$&��U��"�Kz�e�@���C���Rź?x�v���4��w;������^=X�?X�9�@��1ǋ�^��k���h��%9�~s?��--f�W��P8[�&n�;�t��$XC��t3ж~N�$����/�P�Z���M>�w��5+ٙ��(}�tC�瘿Zˌ���ea~�n
��pǃ��
>����R�B�*I���7����6��ع7��aV�屝�@�:�f7mҺ���� �617�	�a�A��(u����A�=�럸REpGu��T���W�CL����!�ᄅq�-[���.��V2)�N�~ѩ���d�E�G�D�-����)�^<���њ�y�9d�%��+n�%7�>!�w.��E�:�NV��$�ۃ���<��a3\p��y�>7TE����Wb����]Dp)�rF��Be?����=	�ݐ]]HS��;A@�I�if�+��rU��W�?�i�oM�~���`������)�pTWv�M-���}��6;�An$���>al�����J��tT����GJ���֞��0�Ʌ�o�%�o���B0�1�$���9� ���=��e���<2/!:�bXؾI �{fj)����JQ,B�q"����4�1��A
ȮLr�RV�����827��%QG>M�V���2͎9z-+�a%6r��*��9��nmʬq�"�]p&�o�w} �5( ���G
��=��O���'��=l�%�x���$m�{�԰�=��&����"K�y�	��>_�7f��{�<G�:�`L�ȉ���O����se0�S��vy�B��TL#�bcPc�	�xAFc}d
y��C�M��W�����,�h!�b�L8M�����F>Pp*����=�Y�7�×�3!&��[@�U `��l�P?��0����cD�ItS"�h>n^]ܑ��ԍ� �¶M71����%��j�r=$�HP���"O��|Y^�*�[V��!��dBeU��L���R[R�ӴRT�uF����Њl�]g��O�r[�!���ˆ���c��`�=���f�i)�c��$@хCvK{N�dOk��D�]	q�>)���2�i�QoE�%Q��q�_P����|�ل��~^��&�Z�5�#��ICjU����������e���ƛ�\�����M=����: cޱ����	��%Ϫ�Z�ě�Mr0���\��[G��'0�}��o��z�&�v�������?Fa�0@b�#�� eg�#���L��)�;��bnD@��'q��`>j1��T�y�:�����6~��&v�q@AQ�U܂���1J22p�<��,t��-|mQld+Z�-��J�qccL�AFO㠗{���[A��V��Ur\��J���~n�yQ�)�>�C|��3p���P�S�H�+��kP�<�9��pS�'����AF�t(TGa��]�IE�(窠��:\j��ޔ6j[uwЫF8�<@���pn�>����mh�y�wc ;K�-왒Ё��P�*�N�anc��,$=߬�q0:y
�1(���틄�Ժ��n����%�}k3x�u�b��Gܧ��ԅ�i���!�"!�����c��^5�����V���XK�1X�X-VN �L���$W���)'�p��_U���i�\Hf,DI��G�\`x����_�H���C��;0C���t���b��*�bK ������s�����ah�=��'5���ղ�3ɻ��#:�:Y�Mr`���wT������bW._C1 �@�[v+�Yp�a����)�3L���̼��/���M:�' �+���&,����Pnu�5d-����
m�\�j��_�A\e�[7��s��8S@��ݙp$E~�w���tʗ��Ҭ>7��Q�f�ǐ��D�X�e�?�r?�D�
�������5����F]x#���Nt���pgH�
Py�=͔�G�Ϲ,h��`K[���GJ����������R�bsVW;��p�z�8��q����{�b4��T�J�d�L>�,��G�����[���c�����C�=�ռ��jz������������w3��F%1CB"Q룙�J1(�5��h�;P��@�j�fm��?�Wsx!!��[�Cd���Kw��њ4��Ֆ%8��eQ�A*?�����~d
W5��9�7m_�!�Wk��=zǩt"�h��}�ܤ��Y>����D���_���sRm*&�g�`�X��]��)1N�l�E�4v���?�1�3��G�lu�c�^�W-��ЌC�Giч�(7A��\#}�������y�[�h�X�ҝ�>��gP<��+&+�'c�+�s���r���Z��b�Q�'� v����W֬e��������b�Q� H��y<�����q%�uG�z�R�����`�d����-bt]�	X���^T"q��=I�h\E�m��Y�$
���s�5xYL՘ah�`�y<0��Z+8-�G�?Tڹ��CC�'��K�W�+}>.V�0*-ܖ�k��@��O�A<l
��%y6��l�cy��X��l���+�kTㅉ��,mF�A��j��Lc(��qZ�������zW�~Z(�_�
u�����E��9;G��v5�ۧ��r�$�^f-���ғ �<�F���� 鋃�Ma⊕��Ie�[�F��nY��� �5�I�U(�,4��$�8<3�m bJ
�wN:�]��Z���*����:Ky�3{�q���g[�-a�*�	�f�"��}b
����L��Nї� 0k�8���iQG���,}�����.6�1�D��5Y7��~�A;�`P�~R�Ǌ�cΩbcQӹ٠����=t��mGW����&k�i�ׁ'�,昏��ڱۜyG	/�C�痣 �x�����v�+�$�l1�x�S��-���<����B+s��ڱ��ܸR "�Rl�Kl�@���>�K��{��C��i��Pzc5d�)6�/�h�%}�����6���q�.CG�T�Lb��V��*���Ƕ�o�@�����h'wd!ijR�nVUPN�s	1"~�3u�룱���#��$�\۝"k�-�z�����1�xa�����qGt'�� H���b,�>;3�1M�O[�¬L}"��f���^
B��AM�m�Q�Zď)����D�F]ją�)��vM���	�G��c]�C1����^����p2jtJ4���}�)fG����9�.�_yɳ-E�����"��>	VvF1�?؍���A�h7�'���0���	�_i�"O��48�7��D����7��GU�{�/
��`�J���^=�?��T��g����R���	w�����:�k�CXv;g�pUA	៍��$�����ps�˜�����]��"��0�6u�г���j�ևA�!��f��M��-��j� 	���W�uZg�Q5��Gt"BlK��b�hQ��=:��uf;�p�N!v�(����E�u����?�*]����P�k�����5!5<!n6f1#F�q��,X��
��uA�u���Y��ޘ��,�l����tu�|��{�S�\2��iV?#��=�s�%�<��C��Az�HK��8'@ˆу;ԣ��j�����t��<\M���E�(��MM�ƭ��!�R�L�i-����`��x����!�r2�)U'�5 �R�$�4���K���/�8�����.��&4،��{��w�J"�y�m��N��+�u0 5�E^����UV����<;̥惊�W���F�e�^*�W��af[��*��_y��2莍G�+����i�z*�����^�����-�9�����|���Q�fS�r1 �E��(֤�D𹔉:D&��1�T��^cbg;]�����/S���x������ax�,9����}L(C,R�m�k���P�L���a<m�_P�/������=IjN?�P�k���S�X鄞��S�����?J���-��V&>�.��
�M���q��#����Ӣ��a]kR,��A5p1���'��R҅�l���h�� ���jBŻ�O�W/M3z�J9��1��f������j�!��3N�#���Y9�����#X�ݗ���t��K��_��Ģ�y�1�q��*a�Bo�5�7Wa"j�z���¶,��7�����
f��DU%͔���kKj��`���l�!Ξ�986B��s�5J\��Z�Bٽ��s�	8C���S��Ŷ�8;��չ�iC��%<��3�%��H�>������œ��,���ۯ)�@�їS/����7!�g�����8H�M��t
�κ�L�v��u�E��_�Mf����(�2o�i�e®���,�M��G�؋�'�$�[�
0���R�r̴��.�x]�3�^��tv癹�dYl����Ť�溒ٟ����6�Gs;kH�o�!���?.�ﵴX���i���,�S0gb70Ή�f���!)u0���䰛Դ��>�OS�;<�H1;���N�u��Q�j%�dTS�X.��M�CgF�11��Mk��kGw�).�-I?/����n)&~)&���$�Ͻ���b��۲�<BTA)����95�	0V�.�k�1!�@��Dh��'t!Vp����P�A�S��o��Z�"���+�q~�W�O�����Ϻ��nya�T(�vV_��>�N�J0�����M3+��h9Ot�"��6����<KW5^�`ͦ㲮P�kFQ��qtP{E��!X��-c��|vʪ�3mf6��.�q���M��4��W��>���9*�7p}��ߔ^�h��O|�z�F#7L��!*ɛ���M�N~8���ǭ�-��nm0���ӻ�`��g���������U0/�����
���n?�heT"#������\�(l<��K�z��(�H�A����f[��Sq�5�v���{{����"=��3��P;(�^�e���]�W@�R��L�{@Y�?���#��ꪡ�ᴙ�?˺}ɐ�ۺ_�*��T��_��U���/"_�,QT�_U|����*�S�-#hE�k1e�5�]�$�P�k�֩��ߴ����}��qee;��[R;y2�ed�������8g7|���x-uG�~�����*�\�P��Ǖ��g&\ݐ�J�&��no�X��¿����>�Wn���39�����kE���>�wt��.�4ô�� #�L�\yY�Ǥg�0�ݒ�L�IS^q�����D���o�'au���W�����q��6�aރ\��1X�DZʫ��c�/Qw��Ŭ���[N�1����k�Ƕޭ2�s��zׯ	�,�iS�i~�	$����A����>޳~Oţ�k8IcMO��.�YZ�S���5v���6��Qg�䪴\��$-�0�c�z}���%f��-��4-��,2�3��	l�rL��S�Q~:I�e�=)�n�+7� 1\�7:�q��2���kA�Q�Oҵ�#q�	�W3ߜ�%�=$��g�ȴ������ �mVA��n�.����|�����{t���t���ߙ�Fެ����|Q�/�#�Tǽ�����﭂%3���@t�@�����W��p+�0{�3ɿ�}g��l$C��[��庐y��@\^���@@�;�i@�ϿQB2_ת��q4ꞺN�7jMU����"p�!V��+IA=pLLNt��ڈF6:]�]� w��ЮO�.��;��j8�c��k���O��:�g���w���vGF��Ǣ��� �؊%:,�0�G)��R]~������u�F��D���	$�3R��}�_@TO��|�Ex�fP$��t�(�='���T�y&�j�g����^��#*��{Pp�g+;�V%���|F���A΀o,��v���Y]���'�L��S��Y�k���l)N�Ů��#�(%�9�6�bU�F4�?F69��=��݇j��K�(mR��)bϮ8	E��k1���|(Q�C�w�nR殨1�j��A��w�E�{۝y���t�{��B�=��/�+�2����N�����g��b�0P��#�|W	��0X^?<��2a8h���cn^)��]�t�}�Ɵ#��󣗢D��M��/<O�Vzy�f�x-��4���Rj��"KE��L%��@�kJE���p�Y�:���_�JT(z�#ݯ�7��&9�ܤf�y��N�"T���1�z�o������&B�:w�R_�ڱ�b�=�ZBŠ��[ҭr�4�M;5�j)�(j�s:;V�!�_5��R�~���l����!�}�ic��S��à����ɉ�ƀ	�$@b�F��y�-1��e�v9b`�i>w}�!U��x�Vz��ݨ���*��3l؅�b�ӡ�)q�k	ä�F=%`Cl��Y��nxLs^�2(@Ԥ�>"VVO�t����}1h(�[�ȨP�W]�*)7,I��o���˛j~��VP���ϋ��,w^�����%���oo��l��$2Z�.5#!��5b��5�LK>T��8�l�SnyɴoJb����|"]�|�s��kFiz��.�8�V���҈�UL{������/=��$`βNS�ľد#�M����}���|'�Fw�eU~�c<^j��Y�muPD^u�����D!���`췿Шmi_�|G-����G#7x��Ό �b�B<�х%m״&&u"�g��ɵ�5R���@#$���r�s��M�7���5��V�4�ͱiT��G���V��Eo�VF���O��B�<���Zn���S�%ȦS�,J���A���-����
�x�h�D�܂�'
� <��/~����=cs��s���[Q{+�����
�2�^���
#��ްw��tL��"�����4�kB�2�&2�p�r��O�-^Ǧ���&ë��Qå�y_j�+(�ڄ2P�UIh-Uhb&s�4˲����lzڟ�9|�r�_X��ܥ�ȣ~���P�E����c�u��f�s�^�谿�Jŏ��\#X��ꔢ�l���^&��l7`;vN����[=��#7Z��$h�������ڨ�n�\D3�΀I8��TD�Hq/�t�g�&)��W�t6�j�������ғ��>��
-�p,Wp�C5�ߋ�\�k�N�� �;OUN�0;		�I��ؘ^%����9f��x��c'�2P��+4�&G3)�d��������/�%l1u,�L�0a�8W���<����^ES�ϰ�q&͸f�#�_L�i�1n-'���Ax8�� ��x�D�
���a*�5Mo/2Fi`��[d��D���(�C��� �P�r�qqvh�4���c�T�&�a������1��wf@( -@޳���D?�(����7<Z�Rh�Ş�;X+1~��Ĺ�p��ͬ�M9}�W<�;���)�uZk	�H�%�0h���n"-i��%k�(#C��&d�ȸ���>p��Q_��΃�;1�f�JD�X�&���Mf#�8t%�U��b|�a���vc��N��^�y�&d3��A^�T�p�2�̿ы?g��5���FVk��fb
�1٘�,%�	���GhRno�0*~�c�' �e?�Ҭ�zU>0ۻXy�ϩ�U&�~L��m���!�R���+�I�.Cd0��]�U#�MW9@�v���Q��/�$J:�٘O}g��י�*��,V�!�{�EFZ3�W.�3�f@��y�nh��Roy�����,�^�vz����Lc���t�-�!S
^�5@	�6�������8�Iͥv���H��8����o/�2�I�A���Ϙ�9P�^��z����^+���oN�%��]!@��w�B�+M>� ���jq(�t�$�Уbׇ{���$b�ڨ�F�|����ND���M�˼���vN��mY]3�������\m\0�!������À��ٲP�/Ʌ�ʲ���������a�Y��fRP��qM�C�4��,� ��()�I���`;o8Q�����m��p��ПN��p�a�q'�v��f|���\0�Ԛ�upz�Ш�(�sX�wP��lyR�p��BXf�)�'s��tp�����J��t+"��Ak;`�yw��f-��&[C�p*����|TR��r|�6@+qZ�t��_d�
�?u�>��#sh�ǖ;%�B*Q�r�,�ھTC~8���~�Q|�Xʛk���D5��˒ z2��n�3{{)vm4�#���[ރ�ޔ?*03�@�5��KVĿ"k��[�g�:u��l{jԇ��4[Ր���-@vM�q랊r��*c�<�o�8TIT!��p���<p����Ev�wA��gL����=?�2_�jt=b5���nB��A˟5PЭ k^
��:w���M�`5�~ѽ��`�\~� i�m7���r1J��fQ���UT1��r.�H��Իɺ84@,�'���^3s
;E�����/��A(�B���R/]�H��g�\�;�L8D��l�W+��o�+s����P�F���y���E����)�_^p��:6��c�0��2w1���<�$��/�&�Y���Z�؜I�H�T�W���W6�	yT\zZ�!���8�<���<��0<�;a�_U�f�Դ��	n��a/.�QZ*&�5B�!b������o
�PZ��-6���X\&#V���f$I}���1ׁ��J 4�w-�ъbo�oz�r�y���1�#�Ƈ�ʊ�_(P��s�l�N�J=g�;��2riei��L��$�Rq.��������Jˏf�h��w���$��D��ӽ���}�7�1�<�1��򥦎���l�
qM��-�]�oS�;��U�J�oqJ���=b�.k�"��$Sv�$�W�{����kHN�\���]�aA����a#�p]��K�P1�[W���QL����+��M�	�1�#
��R���r��}C�T��M��<�{|`��uؼ�tr��t��̴��H�:�:`�B��4Y��o&���|����?���ό��;Rq�/\�C��',��7(�济G�1����y�$S
��|��`�v����#T�t�*���]��"��]����_�8g1H��� m���լ*�t��,kR�t@y���ଢ��H�b�ͫ{���;�8�i�������+���6���7޽�[LK	f�m����Y�Y^)OZ�N���P..�G`|'Ǚ�4_�	8Ʋ����Lrmp�#���p��g�@��)H�G����0��=g;-i>�m�v�JSѩ���cw,Eq�䩡%[|�4o�0�N:\�;��eL<>��5_0߃ho�ヮ?����v45v��r/���?�s
�7��%$�aD�"@3w�~
k:(����b���W�4R�#�P��hA���]r��CV'��UEr;�AU]��*{M~�_T}:�D*��q�YzF|}:)��f͆ ��rm��H�{̙ĩ{Y�e��$Tm�|Qiq�}* �[9}��=W4�#\ �~���:#,�L�!�꫾�+Mͷ�.�Q�����I!�⌙�� �t���r���#:��p�z�	3	h��DA2�{�d9�!4w�=��vn)�W���nM/�{�7�r|j�sO�8�W��XX�!�ߞ.��l`OƑ��]��c������m��EOsr�@a��	!\���c��!Dȭڷl�'=!��%�м{u��y��X�_�K��.��:�-/���8a�愋� _[]��=+%o<.p\!C7�J�Gi��;O(�޾�R������9p�G�7A�G/1\w�%|},�0#�l��O�ʭ�H��+�+�FU��vV��V/�8�ZP
;��S����`����_��.pV�.df��R~�+�>��Dmk�E�nۿ�W���:\�ї���z.ω���8 �/Mh��'=�@PcR�qb�Љ3�K����S��]^cz2�6���%���,S�/;G���
\*�j��:b��T���oR���H ]�gZ��:S8�C2��I�̋<�)dއr��{�)��P��%�Y���W�?;,�I���������\G�</�Nԣ�k��>WQ�>�`�����Ώ����|�J��-� ��Ygt�j���da�?H�S|_��E�<��	}������^'0i�q��O`��4H:�&�A�b۲��+�dQn����=�Yb�8k��F��j ��6j�&m����FD4H&�; �N�H>@iD���]%���H~���x��}��<:b�r����r1�0�x�`_�o~�x��1���u�1+�}�^/үi����9���.~8�t$Z�����<!��78^Z��Wz?V��mT-o����%�^�1'^󸊤C�[m��B^A�m,/��(d�bpp��̬<p��VE���EݖE3�H]$�����c�,�M���N��q�H�%����܄+"Lw��xj��h]�����#�8ա�酫
�P���ⴄQ2����D�}Pj{]�e�X�r�6~�j���D�Vc���,$4��2��6�
������ya|>А�rLu�!)6^�)�mݳ�� ב���?W;�=O>	0 �����/�	�%Ad>�~����t간  ��SF�H�k�����f0�k� c����CX<VG�ݦ�@ɹ���L�j� �4oo��
��V�*��Eۂi=d����^��VJLhwT3���n%�cbT�W�=��V���@���K��4������;��H�*�8��5�
�V���0����ny�wha���Iy<�������Q��̾���Yn��=0��E�����1a�0��b-*��]��>i^UR½`')q�5��ۯ3�M3�����e;YΗ1��y�?�ϱ����U�����-�;C ��웈�Sc�<�7��m{�R��ܙ�ǂ���C��p'�L�E������Q�RN~k���k��O�,B���mV��)#�~ �F	!�R�ZÇZ�0Y� T2��2�:��	�;���9�k���!6򷺸Ũy�eW��+��Bted��2�hXso��|_����R[�����m��B�&[�F�d�L�Z0
"��Z0�����b�N��?�)?��������)o���	Zz�rG�v�?U��q�氆 �w��6h��zX���<�%�R�(�^�; ��y�g6�
qgkȁ�l&61�'�;���13��\��$L�y���iWKa�Tt��y Cm/����-~�z�x*�ݙ�hd]�:�w
�Fi���D�\hӬ�`����%��n�X(�Jו�Q0��M���E�\��$pE�ү���Agmf���EΟ���|��x	��()�d&NK��_�53�1F7�WkXe��XmBMU�:e�+hI������"d��߁�T��8�N����j�m�� �\t[�\]�%���,����1i�����b�_�7KQ)y�IUW
�w����*��<K	\9e��̅�ܵhҨ��~���|;����PΉ��R�� Hu���K7��ت�f!o�������$����u�C�}y�>L�����N��ǅTʖv�|MEj�x��&�NZUZOj��8!2���h#�l(�]��Rc���ŋ�,�v5�n�T���whA`W��� [Ub��ri�D���V]��ֶbD���"V��Jkwi�=���&cUms��]p�%j�D��\K�˻Q!)Y��"��OEy�2��	�񫮑&6n�>/�w1��k�Qg���պI�a>��>�����-촑��d�_C@-�5�,k9|D4)���#�iα靃i3��N흈�$=l�;N�@t%��f�A���2Ww�xiW�c~��-�9�`��	��֨�4��0�ք���]�[�E�sx����8⦴�>h��=j�� ���-�K��(N�\iE"��W_c�+�|���@���P�4�ά*pv��O�����y�����+��>~���+�)�@�hY�V4z�ű���6�6+�1�~���r�?�̛��q�� �Z��>�<���F���ъ쒵�/�P#��������Zw�;���K|s�f�C�9��%-Y#e�6��D����1����Q_P+�5e\�6jrA��F�E
�W�s�xt�"<Q�;�M-.D��#��Et|��E]�h �2�#Yw׽������JZk��P!{Op��<�`!�ޏ�Ro4mx7����`��=����G���am<���b��-����O��t�<VEO_�+j}$Ő��D0#��Ӷ#h��2��_}�?+�\*�Mߌ�6�ޘ�!��\���}TZel���ٮ�i�����M�=�X�DU�_nVX~h�M���x��r1�sʅ]����'"�A��[k΍-e+��]���WuE-v�wd��{�L�u��|?2t��T���z�Q�r��>OΝlCe����fb6�x��'��������3���������{��/���&˸�� �?������?T~����>�V��	
��]ֽvsʗ&R0$��l0/VrDi��[�E1BN�H�aS]�x̔/��eE�!�a"��hAL�l$�Yx1oU,Mal���]&����������F�}�<8f��4�/��X.|x��>�<2�D�7�Ų$+e��|k�+���1G�H�_u��MNv�͌���'i�5m-a�Utxg�K��t��YU�1*!|<���VW�Y�K`�˶9����ly8������0h����Tى}��?xE�����3�M��6vs�����|a��_h�����@��m���4l����Xǳ���j��@���R�Ʉ��;}�B�kx߀����U�/>R���3??�s@��dW�R6� 陽�v7=G��/$�����{z�NTf���XMf� >rS��[���Y�PUn���p�E�E�'A���1����Nˠ��2�,�Z:0AM���\'�4�g('�GZ,����K��f�������Aė�
F|��2���q-�s���[%�ԙ��{x�=_���C�Q���}�T����֙�� �wa뇵��z�Pt���V& ��U#��Ψ�Ce:���4_�G�Ѻ�p��
݊:�����P�sdڲ��u����Jl2M���_K&ԡ1�)U��r�b��5�R�I܌�ҩzA�"�<�ݮq��U���?��掖kg0S�B�*�[:k�|�yD���I�G��Q'�i��mZ<M+��|��N-0���~��}e����q�W��$����bYPOй\_`��IA�*�-<v꽞wJ�>Q������Y����@p�������@�Ct=I������lf7h3�a�0�ٮ��l~�jC�X1�|!��D�-��@��Dg1���	�q���$d)��[��[��.�	���^���ѝ9S�-:3Ƴ�9�+�������!>��,�J��+X]?ʡ�wA`��c���d��cW*�d����@T���{�>�V��U�E�x�0s&�d-R�R�u��k���SF���$��G�
�&��3ֈ��a�DMiz�L����^�q�>w�bRW�#��?I~H�Rp¾u����`�^���J\DG{���v+�yn����sF�܉�[��M��W�h`�����rdrw����h���v��Oa���X#��][@���m��$X}��
���ƥi�K=��4��>#0���g~[>>ovD�y�_*��>gh|N_���8�'r�H�T���!�	r�0J��O��U��_g�[��1�I��7' -U/SKE�{��b?���/I��G�[9~�-��Cf�Nm�mO�a߷�+sJ3���	-�V���l�n���sX�̕Q:B�/�%��p<X��ₘۅ�n Rö#'pA�7M��O��R9Ջo���|Yb[�՚��e3wsU�f��j4zA���|�^�������G�P"2�������=������J�<��5-$��*ə���)@�_����6�������X�:�o�_+b��Mzm,�)xZ�?;�\�%�g����E௅�O�<�XH�i��M9���J%�� ������A��EV'i��*�����D�mmU1�h6�u��yd��aL[�B�c��|6���>��~$�K��+�����V2n�#h�h0P��7�!~8vٴ+�%��,e�2cC����:�����RI֒��}�4QMVR�ۡ����7��{�xP*�1���e03뚟�3���!>���>��2���1��N��g����74F���;�̄A��޸Q����l� ,\���O!�(2�d�F5@7!>G�~�\�!:v��85������d�,Aڪ�4gW� �}�B�.���W��͢��Zi�I�|b"zpC�(�g���5~�mL�h�E-Q��@9(�4�4����!6�����d�}�F�J����#G7�\	�B��׾�#ǅ"�:�!A��kayJ�SÁ��/��~����j42�xt"��%�-Ί�g���n0˽��К�]w�Z�W�6��̜"�z�)�9ɭ� (+Y�sؠ��j�;ݧ�r��3��">C��8�*S��n���H��S�I�,\{B�[������҄�k.� ��,dz���A�K��������BC�R�;%m�vՆV�����W�{\�#�@��3*�t��������;43��5}zzH� <������l�U3B��%U���`�\)����%����l-���>��A�I_O?��!���N�b�N�it-����c_*�.�~�����|1k�$����z�i���E��:�Q�ڭMt����Z�_5M�'���b��|�n�ʧ�N����c�PQ��`n����
D��i)9X�y�\}�l�o�+���הh�{�����������,u����,��	�|U,,������qzQ�yN������y2�+YR�����n㱹�A�1��v�-�+֎��KkJ��j;����Z��Q��	��"n�F�yڸu��0&v�r���k�;�'�����g/�y�=���	���r�C��-e���y��F�������$�ۘ��zT5��/�a+���0
���/��	dԤ䐄����U���v����/}��n��fw�����FpÆr���Jb�m�l��N$�=��X�[�A�(�b��4)V�^���[��BK(K!NQ�t�K�Xy�5ц.1䓛,ū����d�}!�9L?���gi������{�<{��"{�E�LI�]���j�_�}�����)xbf8����
~�v�^�d��
��@#�9��p���
~C
��e�i�Ӫ#="�(�|�Q���>��cgu3��ù8�ǁGn/�n���m{����?�9�!ɂ�OsU�� ���e�� �,ټn1�W9<� �SYL�(	�t#�R"�A���];��E:��#L��=T���wް~	�0��΍�>=@�o�8э.Q5&;��$sΣ� �?����C�mH������E54KC��ܧB�	m�:�|�{��x�+Kj�A(#��W�A�*c1M����+uղ1;����0ȇx�76F$��j"�@A܌>��dOS��ߐ�i���׾b4ozx��A�Ȋ�B�D�������9� oϓN�t��%�ze��K�O���x�*u�|pj�=�/!�$�5�nJUg�=bo��U�Rz�la��� Fh�����?$H0�ǝzE���X�U�a�u���+���os�f%���]�����T;�!�|~�R��K�-�F�� ��Ӟ\��Œ5��Y��B�П���#��Y�KP��00{��f�
��c�]U���L����ZH�遯�1�Х<��V��Kp��*��~A%��ֵ	�H 7 ء�U�Ӭ��Ȕat���A\i[��!��g(�e���'A��7�{D�o�2��H �C�* kkl�I8�Z�����OPc�:߫wFYzu��1�,�֜�����%���N��i���E��_Сr���F�H��Uxlg�w��{G��� � �1���fdK�9��E�a�GSXϰ�ƱSjC�~ƙcyYt�PX�	��o��Y��v#TU5gMJ��ֲ<�t�V��}Ԧ���=ӝ��-�0���j�:v ��a�.��%=�AM�<�Բ��v�7�qMn�&&Gw��s�b�f�B�`��j��T��S|I���t��;���ƥ������'�� b��s���`���?�zd*����v�C�Z�$I]V���d��҄���Po��R�9Aͤ�<����`��+|���F��`�G�YΑ�ي�=�q���.�C�[�R����l͕q|M?�m�;T�`ط�qj#k�$6�t��j���ǪH�J#$G�6N�����?h�OJ��"�1�@������E���a­�s�`�|�jA�X�n��9���ju�����t���Ȉ�
��?�j�0�k	��R�"�ʥ��P���Jɹ��XfE��&�i�U}.J&b?����
�r��YG���X��?
�ڱ�ڒD��.�՛����'���Xn �M�LyS]`{\fc�d��ʱ_ZM�!Ԣ�1��o�T7� fW��;���$�)V;���Л��פA.OH*��a*�m��L�p��9xL���!�� �d9ey:`�ُ$#��h�Z�w�v�t�C �)��Q����`A���ݸi*l&���w�=P�aV�m¶�B!BC���N�M8k��:Ȱ@��s;x�Ñs�S鳡�C2,�ł��L�j<b>��ieX6Q��Qb�S���݅�hc9Ԑ �=RKoq{K6n�cYƐ�8f�^��=�n�(���T����;2d�o�ɏJ+�C�Q�;n�mm�A��|)�8�/U3m_��@lR-���*��t�~���u�΢�Ĥ����7$�F�����IB�Q;�aC����S��q&�DEfk�]a����Ƴr#7�׀�f���+R�+��D}�-�|��r�	vS���Z�f����ޘ��&9��L�6P��C���`ͽ=K�%t�U��ՠ�1���sӚ�H"ෲ`4�� !�c8�2'�b���;�c�&�N_���<�v\5��&1.6]i�S�ZT|�D/�Q&4H|�$��D��\�Z)�V�n��@�|^Z�.�Z��L-8Y˲c-�;a*|��$7X@��w�@���^�#s[_��GM�"F��Ė���j΋_�]r�"di+P��lП�*��+��4=��5z���4:�{N(�p��,<e��1�w<���d�b�_]u�Г�A'���`�h܁#~�Csa��&Q]-Ƨ�6u*����G(T���S��B��'wy���o �2y�$d��vh$4�a��[߾F��+�Fwr���V7��3I�,�'�7�Ţ-�Wѩ�h�v�|#����L����\%�`ִ�E�
�)j+08�C���И��6�:+.P�m'��Bk���`�����U{SZɜ�^��v��t�{�&�;��)"�0.�{���}�����u�j�S����@�T.�&-*���S�S�k�ze��R����5M��BH�c-iRI�9�=<yf譀"�ѷ*6���*�z@��T������j=V�i��lpP);'�}2� �N;f'13�Vn�e6��,��B��<@6��D�?�Z�m8�	��4Ho
:kt|ed<�1%������z�O��z��-�c�㞩Fྟ�i"�WFY�v6�v�(�G�xQ�T��̊�`�e��9�8����`���r�Rdc�IT��#���M�x�(��:�K]	�*g?;O�l:!
���5�c\��4Y�J�{���1�f����s����*��Ks���,Z��hDC�f$���7I���u/Qe%����씥��]Dkw5A�O2A[O�c��<i��ɏ�B��=�Bo�#�q�<f_Ο�빒��C���|a�@�+'a/ý8�������B���f;2�6�ҸB����d�H����� ��g&(^ۑ<9Z���ۤ�L:��X\�#zC��itva+9n��Uu�~�K%�7@���MHР�[K��T��ڵtL��S��_'2iP~L��b/�5�] |�N`�Gn���A�n����y^�8��g<��F/h*d����S��{ى���	����.�s�btc���?ȴ����/�M	Ł�p�Ӄ{{��i�4���i��B�̣-�(.�#�C%�n�i$.�Fa���|vԮ��+yOg8�;����$��;���x"� ��zft|(A������e3հ�"]���KDA�`��y�fkb�VgR��F !�H���Cx�o1�^l���ĸ��(%�G�o�4�ܧ�,�1���[if�,O0F��jı�C�((OM�T��Y�XI��NI<Z�j	7��w��C�J�2��r�ih��wj@��M�k��%�+�70b���� ���J�%��]ǯ�є���W��Gg�ՠ9�q�w>I��>�,��9:���������'�:���~�F�0_M>��ٯq��1&qП���4z�2ccw\���$(��Ny	߆HSo8�KGIHt��7�j�F]��{-���<	�n]��LO��e���@�l8����X7�=�NB�N�F��L	��t*Ϛ��GJ��|˕gG,k8z��-��l�%o�>D����*���(����D�/��a������oe����E��cl`�{���w�g�P�$:'E�EMT:�z�V���I��y��W��ʑ���r�`:'��h�� �����]��+hr��jє*ǿ!����D7�E��N�$��Y�C{�6B�BWh�a�Q�&�0X��"�8�"�'�1/-?uJR�6ReAm��7��+��~󜣤���;|�/�tܪsnFh��u!6Y���o��Z���O9�`ޯ5s>�+j��!�~���p6}怾��#s��a����pѧ΢�+O�ߧீ�#�VA�̍��z����l�Y�a]�	�mP���34	��'������
1��r�PC��Ɣp��[��ꋊ�\���ٟP��SJs���U[���D�z:v^X�Ҹ)���p�)���v�S�e��B����_�4�|O��(m5Z)b�ڏ���V�f�G9���#8f>wԗP����� �@��&6)�,D���_��?�*�t��,&k1y������G�+���Az2VJ��ODE�n!��%k��'��oҝ�>�<0rL��=��[�!mvm�-�N�a��xt�=��[��وr��03��a�';�Q�T_�T���]
|�U�-��U�߸�[|8�l����a.�N������#��l;^o
��~�:%��r::vg��J����4�h)%�O��pFo�l�s��X��ôl���%A~����=}�ߜ~�;����C����jT<A�'��^�D���Lg�6�y���zx�n(bz��o�^�G��4�O�H>���-�)40���F؎	Z��f����W:T:�<��7��2�N� �[��<4d�l�_홋��|�P��J��B�r̕�_f�@=7���<q�2�T6c[���d�"�gw���EZO4�=����Oa�d�W�`�)Q�L+� �G�d�R���3�Ƿ(4��IC�������E�)����A[c{�L:¾�����,>߈���$���E�`�R��tG���
L���7Z�D˹�P+ϴ���F*O���)�P��hf����v�Um(�ڻ4��x�^h2��hU@R�%�l�رo��ث7�1����<�:�d��2p�
�$9��C�nnZ��1ZH6ܦ�Qmj�z}��|@/�)��we�c�f|�Z�L88�hx!,5�ѐ�W@�BH��&r���,��tHbb%�5����:)i$������o�0�lU�Ӛ�Խ�1�␈���@���Y�#�f��g �&�f�N
�!t��-3CF��������L��5K=��م��Tx�8m����vQ�5��Ix�����[�GaOe�{"��ve�6�Հ�YL8����F+���r��ѵ^;И�@��zX��/���$�b2��oť�̥�g1��hG)�����H�6�[ �IU�+�yy��0Ⴣ&X�Y?�a����E,�"�6F����q�?	�^�J>(v��3!ް��+�i�h:ˢ�����e)����ǆ�[w��Z%|�UQ��V���#�82߁�/`����Z�����<:��Ֆ\ϡS�8W�.
j�y�ƨ1ȓ��>�Ɣ�P(�����n)�y�H ����3V�,���@�
#M����Ly�(۞��U�
��
1����3������t�ȿ�SK3SWz�|!�71���=��Ѫ{р�8���ĺ�˟@�+K�b���2�(���1/Uݜ�Y�Zn2���P�����\7�Q��\
 �"��~}7z�,g��%�������������HQ����d�G��Lk�̚���΋����s������5"�cE*zKD��X�i�#20Y�ӛ'��O����@���؍Y),v�j�����{�ﵗ�#N8M7�9N��>��&B��>K��B�����z���N�eC$=bi�8����x7g�����W��q�7�xZ���v���X� x��|ĕD�C��P�i�g�_ٴ� /
�V�p�79����bȯ�S<K�[�p�xn���(��ܨҊ/��.��S0�'�(����y���X.@p"!I;3$��a��=��!wt2�&�K�{奜l���q�ܲ�&��ޘt�Օ���-�&�3GD�c�;z_����<�q��@�scCZD�rcj�$@#�;������|H�qIɋo���:���<�Ρ׊��h��)�����	5�B�o��N��	h;ޛG��*?�d��}^$a�oyV�lzj�"�
'U��i�)O��º@�|ym럟 a� ,��_?~������,� w��W���r��Y&�#��*�� �����g@A���4Z�t���K�6���f�P'&S������5��y��x-�䵂cUBd�B�g�#%ɍsEY�ټj��,^�ڭ-�.6ʎ��?o� �bO�� YQ+R#��y|���!^�	#N3��?�Ԅ~�
D�����.j�:��蔊����j�v� ����S>�!862�77�R�mM?�*��م�B.�c���Ր�4�4�P�:��x)^���1f5E���.w�Z����	X��x{����e�c��N��u�mf܍G]�����S{�V�(��WBV}�;p	`��z���2�p����]H.�ֱ�"_" �Q���-�ɳ*��;��1��Q�8�_1q񎢖x���[R� ���F�q�%g.�Q�Q;����j!k��{{��	�a�L��'+K�s�\��(�����쾀;[�ਓC�z>��z��l���kg��hX���
�؅��\p6��R��l�-��a(m�A�\���*�@���5CEh��β՟��R0�e�~Av�p��-���DiZb�_CR��G����T桔s�����VCs��j��|��<w=���A�HB~1�?��#	:A�?$���-)O��y�9"I���tEK��4�뺿PK��x~^�.�zr�ep��9�Ҟ߿����k�|�a(�׻͏t�GN��xgt�	�;p :-xb�͓�� �(0!��?>��u*�%�(~�{\͛�n�:�0_�)|_Ƚ�NwK�C�[͠fU�����gs^=��6:�u:� <��MT�oM~ON�U=�C;{��������P[��՛��G�c̓�����w����cL���V0<��v#l�W����9T����N�
��sx�ǫZ��!Kb�gB�͵�?�����c^����d|����<�UtN� ��X7�ƕ���b�({2�p���i} �h:k��ɞm��@�����D�ң�j���V�X�H���S�X���ـJ�<�DU����U���-�F�G]��d�Av+�4r��$|�,_ƪV�Y�0H�B��Q��
@XM�o��V�g/���P��E���C�ߝ�2�
��g�B�/��#��Ѣ��j>vMè��܉'u��V��L͌<�>%U����i��4�kE\��.�:�vK�{0��_�T�O�}�N�ilP���V��ZRCq�>!�5zS�F�guBdt��L���B�C�����%H�/''?4GT�PHz�@m
 {����v�>���s�Kg�3{{�A?4v�PA�;�I�pd�F�"0G����LB+k��W������I
 �8�w������ܿ6������o��0�F�y��8��6h�s�mǿM�Ԥ�t�K���9aI<`�i��2���ȄNZ��өpr��hs��}HI��|Q�(�SQ"π́������fE}���]t$g�J#�4�E
anLNk�7�z��3#���|���'M�C9�}0iR�>�H=U7e�y��n�DqYT�F#?Y%,��Yֳ}}�)�4�%��Mv�@��I&~��a�H4g�3�G�!�����G���H����~����K�	V26k�V��Ob��@G�����އ�Mԁe>����4�P^C�ģɋ���$⌢܄#�!�r]g��{wਲ਼6��F������ӳpQ�)O���7ozf���j��������9��	
E� �h�^EJ]����,��/AJ��45w��}��(�"��)/1A� ��/:`���P�'$��>��vP��ߐ����� ����̐�
� ����Kz��'5.�/:���$��LH������ťH�ʿ*/�t�')�M�)�H��ʞ���'Bm�#�Hw|�ga��s7�a�p��D4H������[P�:k]�ŞM,&_��-�hB�[!ۿ>�iRo��Ċ�s��="^p�?댹]9o_�e_�Y�,|o��;z�f�~��"ŝ�߼�ypJ9����~A'�2M��<�4MR7����M~^�T�����I<��	rV�]����9a���{���UK��s�;�����B�ZJ��OQ������
 ;)0��ye̲"-����éx�t1/��/���Ir�d�i���s���DwW���})�ך8� ̊� �6�q�_v�s9m(v	�$\-t���.w߀p\�����R*b���c$��hJi8c�#|��,8:��R�MH����f�����lM5�Y��-��]�?M���/�Y�4�g����s,��S��iIH��{�E27�)%�;��f,CفРX�\�Y��3n:wnW߳��Dļf_e���1n��"�mD�/��S����X�[�lð �J_:�|�T�"�ܐ��^�~�f��1υ8�cYŇ�#��榺���6��+��餩J������2��f�	T7����L����պ�|:ls�O�D��蓺0�0:�5R��f���Y۟kaz��ۙ��0�yb�_v�Z�xe��/���}r6�-q!;�/��_�Յ��/^ ���F
�?��`�vXl_�=s�����R}��ޥ���!������T���K�6Mk�Ĵ*��?皏��S����l�8� NI�����/F(]��uc�V���Ďi�x0���W����J|�|����ǟR�9������خ#�:��w!b�'Gw![�\�ġ�����a;��w�n���vLRɛ�B⁞�_i�U�����8���p��� �9 ����p�_1����ie�J�A��Z�j���V�1Y�h��L4�7�׳Z��.ă{ �Ӈ��m�"jJU��1���J�E$���ၛ(sNk��W���c	���[�Wq}'-?���FF��%ֱ���jE[&�*��dVEx�
����A�Y�;Mа��&�>�� ����&��]��6,�b�x���	�/<�~�&�������O�X�$'�'��ޔ�-.7�A�[��%�R�����i���Ӗ�:g%J��Ф�a�gt3����j5�e�-P{Lo?�?�./h���rڴ�s��q�����j�����������G�ZMoVmi��-��c
�<���wY �xEZ]���W�r�C�n}ʣ�����t뱎.BÊb�Y�����y�=qN�m|v'��xd���ŗ�X*���RQ��Z�&�}d�Iw[�w3��K R�R2?p<�k�@���U1n-�hWQ�g�.�\�H:�W'#V��ڤΎg~���[���8x{˂R>4�L"0��8HUϼ��0�rk��7�����?�l��'���^�C *:QU�?����os��)�A�b5�uNF���{�}ӂ�s�5�A,����d�P��M�^N�}Y��b��,�����{���G�l�_�� ipw���+�1��#�-�MS�C�OA��op����BB$lt)��Al/[�MheV�h@�.���H�cDE����{�*�K�D0y��'r�bK@j�bV���3{���\߆��{ ����W�N�
=ǝ}�G�+���a��s�Y��[5���U4R*4��`[ц��hXf��U��Y�2�K�u� �CѲ(�P��# ̅P�OkK��U�u�@)y�*��A���F����V����B/e�ㅓ�ʈZ�@�&m�*���.!�#���M'��N5�<��=D8u�Lq�>X�{!�s◜�4ك��bf���@�7�&��m����\2� u.�=s���'��*��܃۱�8���U��vTHK����0"Y:��qg8���fa�vH��L�<$��X$�����0�u
/6� ��.I�1QY#���a�].K��H�l�ď��o��� _;d�AV}�s1%��, U�c��-�%�2�w��Qq�`��9}�-,��L�Z*�+���Y[e��4��UO@4P��	�s ��`��y�q�?c��v�Ϛ���}��@��x�����Ѡz�*\�9ɉx(��v.b�&�,��i�b�--�p ��DP�>q�/���
݇���\��c�%�\s��jM?l����q$�3���w�o����V:	RA��n֬����d���;�}�7	�v(���6��HA��}0��R`i+f����p�u�Z诛�(��4����������N�eZ���A2�F���fJj�@d^�W`�����ӧ��mI�I��(c�p	# �9|��s���1��N%
�!�$�!�,�y9o���Q�+"3��jN�}	+۟�������bMN����;Zd<�b�0^OC�3�'4��ٯ�#� F�j*�a����eĨ�Z�xbs�攘G��E�hIZ�ƿ��t�����f�]mX����������c�fjY�^b��R[R\Ҳ3�[P鋓H��tt� v2�ME�U�p�fߧ����F��teX	*���̩7�bh�Is��o���C�H�"B���� �Xu�������� ό��ڵ�����okW9W��m����n���biG7�vt��j]E.��t��gqHEd��N2�E�}�k-�6y��/]Y����Q�|��)=P��Օ��@w��"UOdWa� �z%��V������He�q(�8��O/���K�fd@��A���
�����a�!e��P)�ߖ�1�����{¬�nK+���5����f��ߺ�"A�6�6��Mw���V"4X���?jl�E(sF�t9G:�����$K#�[�^ű�Ï��r%s�Xh�8��Ǵ.�$�{��4XV�����T\�g��?�4�Pԩ��M>�ƙ|<
�J�G{,%2�� ���%1�L�LM���P��E��Z]���q��?��j�=/��@z����*i}\�z+�|���S1d��Y�_y�h<�+��2<���Ϋ�)b	 �>���P�CeT�#�����,�&`�/JK�%��`$�K(��|M�ix*��g�Xx#u��+�E5!*�x�w�n����D��7��h��1>���ήcs��7Y)��Xr.�l�5bvF0}�_qg�u�rͲϡ6/� �Żc�����Q���!hR�r=�|'�{�~-E���=�]�k}+�D_`��dg����%�Kb	�.�AKeͨ3n��S�/���um����`�[���M-����8�Y�� ~�zp�4D@Dܺ�A����z�%������R��q��$��7���s	��}wq����G8�����\N3����܊5�������!�h�:xxؼIB	a�=�����\��ul1�=v�������a9+'��L�'�W*hٷR�/���.�;O�?�N|\!F�z�y+'�������ߥ]�i���̺�I	�t8EN�+
�J�������J�A���w(�����m�ޱќ,�q�}3K��V�X�"q����ZJ!pl^I�q�H�7m��J���
��fZ�Pؗ��=�8��Of��)��e1Ki�PZ�?�X���YPvQx�д7�B���*���A��%����v���o��h�&m(��q��RtS`cf�֤�P]L������ll}���G��0fw��Xc�������It��%� ��a�ƮA�{ٰa�*Ls@,Q[�jn�
};�G�t��"�$���e" JJ1�:�*�Av�w ȗT���,�q_��F08����"5M���jj>�)�i���=L=/1�y�]����l�;�nʲ�q5ߪ�Ž;��-���a����7�2(��"��fE&��.��`"���MQ��O	Ҽ~�	�0G�3�G����B;fb�#��y�2��f�����#d�,�Ĉ�~�Z�Gꆖ�Q��z�d{�\U����`�F7��"���)�>�h��w��X�.9�i/��]�X��\�9���b�
�8�k���5a�NQ:���de��.�����)���\���T7��)�::l���>p��{�3� �p��c��������U;f>1q���ԥ����䖞�_��1�ЈO�hE=#m�$�7d��I�<0�k˟;�0�]u��>�]�\��+`��DE
�j��F;�k�_���)�_!�������g7c��k巒IS�{@v��8����mi�	_��|����YI��J� `8)�7�G�0)j�.��b����&�3��ڏ�*����S4������Z�{�ՙa�e�:<c�Io�EU�awh���@�"�j"�<0Κ����X����9�U�
�?w�ĭ�C��c�u�%�︄ds�/Q0O��������(��m�8��o�l�ݺ�D$�A���\le�M�uv�~I1�	!���UW�q�%�g5�ė��\�[��w�̅��v8�>�)�`|��]Y��v%i�Q�U�����Gͧt�%b�G�P��Ԑ>���$/�ִ�D^rƸ
.����P;&v�]s�"5��4#���۪��5ND#��|����r�o��H�ۍ��1A}y�!�2;��H��,��v=��}UT^�foK�o!b\�E�[�E`�%v����;	���:�ԅ�-�9��ʜ����жp�R�fv�Q&}\a�>o���~*}����\AK�D.��+���Th�1�����̚�;�E�n)`�A<Y�~�����Q��[�D��!�@�Ap�W����$�٪F�B���=,R������j\��~��*i�<i~�:�)đ����*!|_�.�"��Q�&���WIYȭ	��M�9�^�IO�0:p �y&��3#w�v���7W1����EU��_̶��,��@�76��/ͧ���%?Y�^u^����ь�S�PՒ_�d?����0�%��� ;Ȼ�J�}��0���F�j�ڭ��@�J=��Ї��27h �)���\�u���)���T�(*���K�gg�$�"����sd�L�\�ehT;�e#��Q�Χ{V3bI� <���fpmkXiq�����L>��Я�|�pE���n�M��w��X}�P�0�X��v��E����T��>��i}h����s��9�>]����14�9yh�Q�8s>&#a�hNh��d���@����@nV���<��FH�󒿞�7X$��zl�	;̗Y=�o\�`%����}X���*�.�5���@����ĵI�=�?��Cޭ}7V����5z|��V��T�~�
1������7�e.�������	tU�"*�N~hr�#��g*��Q���PJq�|���?�m���8iA�-�y8�!ߞBB�>�F�M�F8��tH��J	����>T�?��G
��O8����nN4�R�t���F��5wRߐ��=���WH���B1�a��Æ#���z�-�!�㎵�[0vܑ`��ŤaYQ������"���"��U|%j@~�0�WTQ^����z�6-�"/N�	�`���=���$�(�U�,^��w�܎��
�84�x%b�k�sES'|]����?���2uJ��n����v҄OfoȰ�?VdD���Wr�xͩ��wK%����!$���&xbm�P�:��y�W+Љ��*�=�]y�����!�`z����~ֲ2����W��f�m�?���*�o`��d�x P�����pb�2z������(� =h	�ﯘ����.K�WŪP���Ƌ�]�"�pR��ws2��dB�5�}�����`�*X�x��iXF�<�b�MC�}��I��v�[�SK��`ҚŁG0��f��V��΁�����'=���mV�"Dd��S�T�����s�}���2���c���i�O�]K����`�/�����1˺!�X
��"�v�O�Z����n�Z�ru��/�^��k�b�N^u^�d����-q!���X��^���Q�~��Ԡ4�2!Q�Ι���V��|gw��<r����)�/I�
ۢ�s ����)r��i�K�����}o0�Q�S�����<������js����ɠ��<���ۗ	��O>/u���|1�?L^�V*�����r�
�|��2"g�5���b��H�q�h�D�d�Y��D��������˘Y닱N��������[�#�KHWp�>���77���5K
�d��;<���q�/a�ތ�b�'��__�'������'G���0�~��o�Y�i3-&|���{YLْ ��(�܃�>!��ճ��@J�w���E���X�Rw{߽6fW3En`��t�1��x�<̫���3I�ĴA�
	��=6`���m��c��Ј��9y��\��yQ~�%�F&�3v����<������C�.�)8 H��n1ƛ&ZZ�:�A�e2�ۨN{
bE'f���׏lͶP�O{/��86����R�A{7$yP���U��.8�K�D3�m���_Ak�J3\��,����;4fO ��p��Q��Ju�	|o�C�#'�� A����VB���`�]�kF�JҙF_<�ҡ'w�jl+�M�ꤑ�|�%7��G捦��Zݱ��|��fr��� �ڷ!��	��5LL��Ѹ���N�a	�[����33|F�S����ѽW�ծ�`���Q����b0`�����|�Ӌ	�1�^߬ r��S9�����50@x(�J��YX3������ʾ��5���!�e����Xc6�/sC"Ό2�����B�-5��J����L��i�����
�G�S���v10iI��3��ʞ�
e��aH�#���6�^?��O�ښ����s+��_���I1��c
tXh�����ތ�����d��<�[��s[ÇcsS�a���v��F[ه0�I����+�ap�Z��;fp���'.�c�Uz�@q�U9N����D�R��!����j�i<�GRә�I�0[X����@��47��A�No�� !B���|�������2薊��sV�,�A�v $]�zs�M,)"��e_:W�.#O���";9T�16t��a�?�8�dCQ<��a{��r�o��o��j�ڙ�>6	��!h#p߬ugj��ݔ�zcRNI��(F
�Dl�E�N@���
�ԛ,�]����`� �����-u���6H�P�QXC6x'�6	�8�G���@�l<�1�;bSYƩ����7@�9�U@����R;��[:�����Բ��*1??w��:qE��� #Ci0*δ�n�u�����z��Ü
]��f:�B@��̯D���NL* �>��9����B����+O�;d��#�V�a䶹�͟���ě��o	�oJ�3�N�ϔ'A��,_+�w(�>*�@��9���l.y�b��w�����_����vŜp#膮�x��2|H�w���� 3~��^P�E����0!��ķ�'F. �[�  $��u�B�����L6�P�Y= ����1��s�I$����ӟ��ˇ;�Z��I�A�2Z�Hw��NW����g��M�$����1U�EёH*��9M�$b+�e#�	�ɂ�y��{f ��kʦ���G�!,N��>gmû�HH4���j�ό��ȍ(}�@Vn`�RO� �J��2�eQ�J��7CEf�=�U%�"S��E!��|�t�T���$��ÔT�K?�Q����V��{ZY��I�v���G��Q)�Q�+�l;&��^�m7���GQ�GMJ�\�+�jqYpK�*w)Y�g��D�q�
�ۻ�*�E%Q(�[�T���
�(a�e'���uX�������'Gn{n��ky"�f m�?�C��5��H��(ᆊ�����D֥S��ϴ����FzFDB�ZE�n�E�i�'�Z��I�� Ƽ�����>�`�����v
+շ�L��,��_�8�����s�`�O��|ף'��$|Dg�^��x4��R�~����&�)4�fS���R?N�Ћ��w�'��
>�o��2E�$\�c��0^���nU,=Ϯ�lQ����%��X�X��w6�̓:�k�D;���ak�Ñ���edF5�&Hƪ��4�ͷ��2~��\M�C�c:�`^�M�D�$&�[X.�d��C��(99�2��Z�oT���%�ͭ5��,��.{&��U��ry,M�fE��[�D?��o��ȍ	C��r�NC�S�tU%�j7���'�9\�6�&e��WpS��>a=a��$�=�@CL�0�D5+!�W��$��Zw�k/#�ｪi!*1m�?�[��Ĝ�F1y!�� �é�4ʼ���,L}��{��~���a5D+��'^M���:ų��E�H�%�}��S2I���K�4�It
�K�߉7���S<���(��ó�y�!�qn_1���);��$��I�S�~:��Z�ޟ������$玠��~5J5�Z}�
),�/��]��Θ�!p��>�
9q�M�z5,t�:DL~`�s���d�J�D,3dd�^q>�	RD�Sy�,����u�r��Q�ʌ;����령(���s��i$@��=Kh��/�_zf��uV9J"<�~T@ە.�r�w��mF���Z��]pe.ϰ���@�aw�����W0$h;þ�����^���Ä���e�m@Z��˦Nݱ]���sRO�س9�C@ou�;�%��M�H�n�������,Ѡ[�[�n������f���dT���
�D��l����G�X��������h����w���:Ek{���+Ŭ����t&'ꜦT��F�tpF��o�d
�X�n<����L%��^�6�%�9 ,�0��?c�+�7cB�ow����]4F�R�`���q��Ut�����
ǭ��<�`c����Vy@ꖈ��!�,V���T��8hOt��-��]������&�rǏ��Cd�g�8�.���A�̟�T8NN*Hw�J��#�9���n�[�O�3Z�*��&V~H[Z��H�S���]�Z
�+:QEb��9!_F?-�X1۩���i&�,R�6��~厒w�� � �i��:E����o�Je�@��f|֛$#p��
r���Z�Xf`�;�4�ZڑU{��H���o� ���E&5IVO��Cc�x�O�m����lQ�,�3/�,b���ϋY/?J���M��۽����9^��r; ���;4�ܚ������R�rg��?DZ>I�B���䑺1���M>ݨ��ˈ��:4�\���QԨ�~�@_Xfz��V�cö��~�B�E F4h�Q�Y����j�qG�>���}�$���s����n�)�
VW�+ݡm�m���
ΰ Fr�t?�唺�_Ė��� zUB��-8*z�cez��Z�Cb���Zʷ��fߏ�O�^<��3�&����ʼ=JC�_���{{p)L3��}$�9����V�u����pӸ�$���6��I�)���Z�v �ɭj����u#6&mH ����s��$ N�w�'���<v����_X'�w������Qv����X�ֺ��wЧ�[��Mh���r81:�D��������ȍp,2$�^G�H�3xT���ˍکc�3�ː�fuw�=���ރ���B��F���@��D7lђ�f.ϊuZ0�?^����d���9�5:
niC�
YY��&?��wV���3a� I{�&��ˤ}����<�8��as�Oe��s�װ�~��k����V�%Af �sٺov�?�������L�����|��c0���+��;e�e~-�kFk�3p�Dz�؂d��,֞�g�.�����j�i
d��%������ˏ:qJo�h.�����
�/V���_�ҵ""�x��Ϗj�B�f"�(��O���~�)lS�����{oF��<c�'wGl�����^��n��;��=�u_�>��T��@�@�/���Z䌲�d�3��c���4n�1����~�0��U��dm�0�V�)G��6�+Z%-4�<��J0�#&z�N���i���)?;�о����������S�f��{@�d"�AG�O�4��gd�hN��! ���6�$ ԉν���4O�+��^kF���|a��B}�T��CD&l�c��+���iH�lU*��i��Hb=k��1xYD�*I/�,8#8-�Ɖ�KA��I2ӥ3���������lĞG�Z	�b���@������ٺ�.�^B��G��?c��^�����^�*�
���L�g�� ����R����%�t��(Z��?3A�|T>������+�kI��o����i��y��t������-߳��.q��"����6�+x�$͍�몖������=��(z���n%l�a ��n�_ MD�n��;t��'�����-�2�=���=[�$1�5k@��]L�q=,��o��l����l�����@x�]��s�8�P��ϥQ�e|[s=W�x�ON�0o��R��z�`FooB�|�J�_�����ȑ�c^�>�lm��O�C���O����O�d��c�Q��*����zF�������Z�w4S<A��G���={�� 1����^r�l�z彾���Ҍ�w�A�=7�z�i���[�6r M#���ETw���&�8�
���FbfD�.[�����M7��T���h��(!�%`�qpW:�m�������=�ȗ�1�ժ*39n⪞v�r���1ߖ:�o�$�8��\L㱅㷅7 ;�^t�\͟�u�����jF�=#�%��?�b����6C�����.d"_�3IVV�y^x�?Im�8�y�/�y��2<Crn�_L����μ����}~�_��9k`5Q��M���a��ܚ���g?�i���ǽ�h2�	��xX_�Ý}͓E��\�٢�}�¹פ�ቪ��9'�FD���w~6�FVl�������h���;6���a�����K�8�'�N�FH��\��Ì���5O���y���8Xn��#��O��HZG�5�zst$�d���@����)U.�7I��z�ޙ���ĳI�<�s�c�U�,�6p9x�e�B�$�Kldkx=� ;[�YK���c�?��Ğ�Ua���SX�i�R��lH����u
0h�V�� ���g*F�#|�z��������I%���;��o�*X���$[s� _���T�V?�z-�E�0
�Fk�%^�o2��s��dX	��샰�<�<7tϙ�_����~gG�k��^��?[V�:�7��zm)��K3iҦaW~ �����6֓#�y;�},Eyy4�YH�1@�[s[���Y�W�]���J��ϗ�����N��u��c0�GJ�)����`5�"��;	1�V]�ـ�J���0���:��5s�����Gk�)U� ���xٌ�E�6���$I嬄jv��.��k������$.H�>��
q��J�!�m���>(�g��m��8j ����X\�]$/5���}�o�R`�k^���ܨ��Bۊ� FXݺ�\w�C��<3������?'�۲oc��+E�{���4@sYcU��  �G��`-f��w�c2r�͉q!#��.��ϦZ~��Lߏٜ�5����`�OB;�~���s��Ǐ��-=�UR�svJ��$����G�Y�l<�����Ξ��}���_R2ra��UC���ٞ`�M���n��Kt�k�H���W@���A3
�a����]��p���>��Ђu�j�'랸:!|�W���fX�;���ա31����0�d��2���^��j]�<��ud/F!5�Q��*ʏ�ٯ�P��J��C�\l!�F�d�#�a��z_�qO��.�K����ώ}�Ɖ�
��?SOH��ΪGৃu؁v�V}�L�wԍ�w���i�ҽl�5a��	^&2�w������|ղt7F0"��ƶr��i��*�v.�m��T=m�Z�^��6�(�A �k�%n ��Ŧ�#Ux���.��:��o�[��q�H�SǗ@I1�)��`#@� F'�Hs"VR�!9it��o����O�	
��>U����Ӥ��������Kf���n�e�W��Z�F�˷	D�'���ODpR]�L��~���ӆCQ<\�?��(�`rrt!�D��q��Pk��ʥ�G���IS��hԟ�{0<ς�R-^��k�?�G݁%�j	O��D�����2��JQ���<܋,iJ3-�P^�7��-�[Qg�D`R��Em�:��w`�1�s�r�
�zz�\��dpU��?49��I�(U��E�Wq��� ���'����!n��xr��˩����o!�+?����v2�žO�U�
��H=ȁ4'3����!�����
�Ip�r�"U�߄�a��f� k6%�o3PNUT�&2�pw��q�o���
�4���v�-�q^0�'��yB]K�
߂Q^B�Q~�.�Ԩc�6�TOW)~ c�\t��Y�P�|kƒ(e�9����Ԉ|.|�pl����d6�_�z��&�V#p`8p{�n�0?��z�D�y�K#j����/Ȟy��@�!����l~d�n��*L "⁳���8_@ӁƦ#�e�G�,�G�?N�Q�"�r�M	.׊=�}3�Zou�j�R&�OJI~ّ�;���s5��wUt�7Տ$6�jU+�W�L��CJZ�(�ͱ�;���V���KaU��*�B��T�[�T�|'=s=�SHNYD�]��G����q6^ܼRp4{YB�&;tG���+u`����j,X�A��r-,ȟ|�'�η���K�0�ON�i�p�Y��6ZY������W ��%�2�O���m��T_���Hyk�����߉CM�[�AO$mo>��(��Y��üdn��lP�d�����e1U��0ԧ]G;��;�*��֥�])�l�.T'l���q̼�D�J�K=�~D�7+6�ZԊ�JT����ԝ�.�}1ZLփ:і5�J�XF��t�$Q�A-`gx��)3��a	�&���~�����VGM�Q�s�B�d���+B��P[�7��5�T��y�Lp�	*�k0�=��o�-���w�D�rƃq;K�b>�xy:lI��?/��ك����.�-òm�5���l�ma|Y���@�S��h �LP���u��*�R�۹�y�Z$4����%��H�-ۡ����R����mӣ��i�����g'0ٷh���M{�����C�i(�]`SPSe1���7w&d�a vx�=A���J�1�$j����YVG�8���Į� m�}�I~�,ʹA�W����U�g�Z��d�t�K����{�jMĨq=|�Ϲ���X\x�f?�a#R
���Q������T��[)�q�bE}Ԏ͐.��.���$���I��=�o�.��̗7����;�T/�w.�Y��p���������E�S*T���JG%���ej�V�!��ѵY�
p�t�x|C��Ǒ}�l��NqK%d%v1�v�Є�Q��V���9�F��U�W�G�c`�[@��`�1�.h�!�X��٣,y6�D֏覔āj��X�i���/�ϼ�A���	 ���a��#	�D��S,��y��-�A���Ϗ�8f����\�zJ/��|9���ߛ��f
�����:�:�H�Z��Vۖ''2>��rL�)�@_u�P5�m�$�����������4=�q3��ܝM���~�_|9��~�H}���jUVs{(��Z0�tA�Bf<(Ջ0���eJ��Q'� �V�SU��h���Y�ML��d��Ȼ7����x���Av'H�/e7Z	�w�kD_#���5�3|��s��H��+t�{���2_ҳ�=��8]�rF3Y.bW��<�,?����~������|[�n��y�:P��:Av�P�`����f��Q�.;��%�)�V�C`��i&Ub�5�`A ��2��-�JS'g
��K��qe�N�;��jy���~������&����ؘ���.-\���A�b�����k����	��3��\���Ai�A��H�!����T;6N�<T%-_�3�N�pyك�M��Ľ/��qj(l� �*K��`�K<;1�����utv���٪�Y�Y��vZ%'�Φu����~9�G �\�j})� ����f���<�`+��Ի���g�����@�f^�~�%e%=~�G��E����f�>n�EI���w|C�v���=�"�l��E��Y�8���Ǔ:�V�/	��&�L����T	�Yv��a�G9U�����5���t�����Z��d5�S�����q�2���t[�T��@_��htz�����o?
�-�Wrtm������`�$M,��BDL��C��\�"%6��#�#�롞�}>���	�i��=���9b@ɵڙ+f�L~�\Y?�	7�{ 2&�4�o�+�A�_],Ki�$�GlJ��ןzʔ2am�z&�H��U־ד���Z��=�&3B��@yY��m��N��|b��I*b�0�AB*H0�acC�N��T��))�)����ڇ�׹�G�Q��(����j/��wk��ut����`�y�L����b/��"����e E^
U0D1U%��"��S�%{���5�^��k�;�y�/��N����Bf����zf�;��{�c,}��t���:����Z���6>�q@����y��s1
��d��~85��t)�aQ%J1�(�~�^*EP��
3w���6b�m��*r����L:�^�I���򒋖O�RH�1c<�^m$���5�J��(�-�<LE�����F���#��,^9-��9҇������hx�")j�h�)65Û*�C&d9�Jm�f�7���#�^��s��r�}�Zf���`�r2�/<.��z����ؠ(C�ef߾W�~ƭ �{x��]����2��*y,D��GX?���?y���ٍ'�\��G&���+����β^���>��%ў�q
��W\7����(��r҂��6��Y,~�pl.�
�%�cq� ��ت��U�f��]yO�q)���[��hSe�χ��4,R�?>Չ
nZ�d�V���>�A��GO�G��}G��F{^��;�f���SO��C&��1��hi����q��0l&�sr[�?T����0�_Sd�Eg��BU+�W�ͳ�"o�ph�7���'����h�ti04-�m.�W�2b�X-F��T��d��_
�����D���M(!��8���d����*� �پIEy�
Eh7�xq�"K�1f���*�)�5��3�� �͐���*%��YN5����T�H��� ��ߑ���I��Q"��"~э�C9��<������2�QJ������N{�d�Z�'���dH�xq�Ns�WH��$M٨��&V�7Ȑ�Q�����}�tE�ܢXۂR ���cP���eEp�>ZC
��</�?�~=�J#N��_f��򽼓z�[�����b�m�y쀇�yH��õ�t�\O�<>���9���U����B���B�#}�ѐ��<�^���hJUg�T�>�oI��X�d;5LBbn�q��l:���ۤ��S���w�����|yF�7��9w��������]�U:�Q����X��X��Q�D��b�A�����3�̆�������'M�ٽx/��&�%q��P���g�whO���t"��v+ 1U\����=A�j��˗h#�D�,���;�Gs�[�j�E���z:�%�_��el���c�W��-���A#өF�ưF���v!�=O�
�j�{չ��M���K����ׁ5lw�����\��H�ٴ��n#��&��8L�?��{�-=b��Xhe4�כ5�/�u�o�����ܥ=���?��z�������R����z���� ���h��V���	:�>��9	�y��4�x|�}��&XH)�{E��$;Ҝ��DI�VB�=V|"J��ι�ӫ;=��X ���?�5@�rT��ͯ��"�R�m��[`�x�B�<$�4ڧ�4�0�Ra�f�=��\.����ϺB�i, �+It�_��	z*4��)	1��'�40�In��gklK1{�' �qq�'=#�_�`��F\H�0ch��L� �ߛ�h	놮��Y��8���5��w�N�����J�(�x�b�U�6I����k;���b�J�6�-��Fh���M�g��e3�[�ۥ�� �ݫq� �B+A�o1�dd���|��E�b{��h�l/4�5�C��g�E��R���4YSg�M!���T9L��_��~�6L�ɴW��0�]d�qP����;�O(b�mtƨ�KJ������
 ��	���>�;-.$RBbX0{�̬EUe=���S3aC��?ۏqL�g?|)�Vݦi�⫓Zrh;�|����1��/!�U4V
�BUp|D�G��{���4OH���ʬ�kw0�.��L�.��f��,���~-Z�\՛v�t��]�$'���	��3�"��d�\�x����ld�&/�DvXalE��NeKL���-��r��&�
8^��xJ,4o�4�3�wk�(諄W!R�H�BO�}����Ŭ�{�̼FĽ�J�v�Zs�1 �P��Y'��V΍@�(�Cu�Ş!Aa�h��*6G�3C�L�K��"��3����}#�Bĵ��W/�c�)�W^ �K��?s׳�A:@�yb���<ȩ}ctz�t�!kHF�8]{y��8|nԤ����XB�a��hk�t���.��� ɭt��">k}�T�d D���9��6\
O�w�
�-�[��5;�[��������T�-��j�g'?!t��p �	�C� Ta	]���t*�~�;p�kd#"�w�P�S�/��e�[��E�겫+���C�K͛T�^2�^b�x���6��V�mo�n��	\Ei�
����y�$��?�����ݮ��acW��l
i�ͅe^%��E�Sr�!{&�������G�W܍6��$����;T�������ǧ�b�e>q��0�k�g�r1�� �ߞ�W�Q�{w���20�ky 3%��Sç���Y{���1�*�1 F�ը��+���e���t����⿮H��D ��m�Ɣ_*-�3�K�)�э|5�D��[��d�՛�HwR��IK3x��w
;H�Jc�+�����1��BZ~�D�>�(@�O۶�1�A�>�Ǽ!2mQ� n�FGBa;}�OK���m�0 ����E����$C�U�v�����@��
2��DZ���?&F�ԭ��-���b�kOPm����?�jm�\l]���w��54���?g˛����P��)C�����4e��_�H�m3R|���S�%~��;~i����4���,6�DQ<����hAV���5�/���'�]Ih�3����U���S�N��y�tWg ��t��D��N�����Iz��P��}��	�oc?!&;�ND�i�Y�O@9Y~���z��#9��z�~Md��	J�g��^<�Q��iՈDFB���N�ƕǳ���>���h���CN&��Uᇚ�JuA�Ssh��j�nY�֬�c����Zw!�CR�ᒃ������JѼU�2���"8�u��?��z�-��[�_�7%����}�e�}h���j�'L�+�D�Nm�?�@u���A�k����,B����P��9B3������v`���
"T�t@BsЈ��<�P���ⴙ�w#i�\�������G�F��=���5���AvЎ����cG��&���	�"��)iXBE�
$��Јu�ߜ�Dqjz��w[�vZ~�ժ�.x�ah��v�,�c�8	�1��F��k�=���FU�m3�K���R+�=g[��{1��.�����?��1>�B�唌�Iǃ��Ư�ʊV�a����%�s�v0��#�&�����/��_� V�谜CT�Ա��� x�+X�T� nK��=��\
ɗ"��_������ �ƥ9�����t���x<& j^r�㢬4-��[/R�I��V��ǇV��o�
��ؑ5nt��C���:�6�%��ڊ����q�}�p�u	yc�k`�)�hQR��}R�j��??���P � �Ƞ���LNo��m�k��@﯒n!�ےb�-��z؀�:��TS�ɜNՔ��c�G���k	��F��g����	4���7�#�n�@����I���j�;��/�Rr�7�-��6��P���`�&Diƨ�7�bcy��j���<+�h�ҙUKy{��z:$ڵ�Ç���톸B�o��'��/m2����1�{�Fˎ,���	�|��^{�:���&|��A)u��9g�.�9A��< [-���R�zup�#���G!�7�wǉJ��) ױ	��~����A"�i���a�פƽhyI}ãȈ0S��k\�Pj�*m���t؅�yu=k�F�)���70٢Rnx'�eGs�5��D�wl�޴��G2����se��y"F��ڪ������)l�F�̆I5Q�������}�V�q_��d,6������7@�Wt��C#A��
����7�8�chTf�`��>W� �c'�Jg,�m!�z� +}�p�ih�^xJ�r<��ڮ�o�Au��G�@f&���`�	]��f�Jl[L���pK���ʡ��V� bD$B)���n�ٿ��״�X�=��X��d��%��l\�n��������:��t�%/MIQ���!�&ը�u���n�+2p��fl����O�jr�Z�7X�F]Y篖���	�m���jF��4���Uͳ�־r�kw��p��K.���X?-��U72�g7������M�Άӛ¸�h�I���ȩX��!;vݴ��OX��W[\�;��x�m�߀�[J�όm~,ĤB���&E�u.ުn>���%⦏�/�������腪��A!n�C;){��̯��X�f�ޭDw���o� �Nh��P���B̤Df����N�+��Kي='~���!�׿#V�ZJ�+N�5�9 ���!*BW'ƺ�h�x�R��EK�~��a ���a����F�eG=~Φ]�R� �g-���b]�&x5�	�|s�g����V���+��i���5�	����}�����}Xz��sN�}Ay���x�;�l���VG�Lp5�qHUF4��lo�&g��RoQ��8i�.����{�5��`|\��9�n�<�ëJU�����xM��5�x�� 0�e�;��_:�z'���?@�[,7ʘ��#��!�aL̈́�`nǰ�^���9L�����96��9O�PŰ;p�읬!$���$ʟ�*ɞ�.��v������T+�d�.I6�Y�N<�'f���n��F�ar��80�_���P�^#��ǽ~�s����<i�}h��x��B�l{�R[���c�2��p�F����A�e~�����pH��	�J�06����|�m���;һ�5�����]������:�~H������
-�@���B��A^a�h�6Ə�]�H�Z����F��� kK]:�.=$�I/�`�A+I�x@�}%�)Հu����.ߺ�u���a��^�8�	i+��̭��:����Yߔ?��߶Mt���H'�t^��8i�J�8��#�4����)�Tc ��\���w�ک��dJ�?'�L�)WK=�`�RCz�����Ŭ�[��,#��7g#�N��Q���q>���U��8M}q*�(����u���V�Gp(}� �j@�:�g�\��2�%�cs�N���Ԕ(��-7*gh��aYd��6�8}��R�� ����#=|@M�U��~�r瘥���8��ҷB^^|��T`�e�y&�Q�[��q��PP��Z�ź��.N$z{2��Qac1�f�(���QL<������9��٪����a���+1�9�$ֳ�΍]y5�-��:8����!�-e"	�Z���rԂ�!0Z��/���m����]h�m�>�l���Ԡ���3d���v��t���32���.��Kr~�QE�NV��LG��NSM�r���y�'��B���;Q���0~LP�I��x����Yy�/4i�<7)�;m���y���}=	tTK�FP�t��{���j'%�`vq�G��O ���C���<îpQ#�c��V"���W>G_s�A��]=���]1I��(�=q��E���y`�}�P�\���e1c��#(e������S0��;y�j���N^�D� QD�K�B�|?#C"_��!�X[d�&OL�*�B��鸀���ˋ�^m�A��k�}���o
���� qSE��W��_	Vk�H��1;DaxY'
?v�R�IAt;b2<�. D^>i7\��Ko�����Ɵ�Tne1�8k��ƫ�dky�:?������\�,{�����ub�^np����Y��ץ����%�	(jX�v�w�X���t�r������LDf��x��;܉�̚+���ʕ1>����YD��6��`�#
�[0[�ˋ�pړA.)X��t�tW��?�@3�(aOس�4Z�I��y*%T�=��q��_!d?��'����jA،�Q����L��`��*hL�d؞'^^��.o�9᩸՚e(��R<N�[6V5��p�F��Ӱ�{��J���*:�`��C�a1`����S�Z�K��?3����X#r^j��T��A���˯WW����f���NF����rR860���%X�cߡl8��%'~���i��!:��F��6�@ן���a_>��c������z:�qu
�Y�h���RA\��}��#C3�(��i��xb�>D�2����é�*K���]��O-��耊�N1��le)��Ct�b�(��tĭ�	:o��1�+s�ĭ�PJ�9��xʛ>�̐�W���aO�C��.}�@;�zR��<3��L.P�#�n8;s%�y
<�uU��j(E�jf&@������Aυ��d�N�s��J`	�Q�q�d%v��4���PYq��+�U�j��ci@�z���*@Cd�X#�,^���.~k�_>P,�$۱�q��Ã�7��i�#�i+C��(W��q]�VyaOw�gFLQX���9oM��O,�MVD���6���L-*F��IP�b�o]:PDD�+�k���W$�����ja���,���n/�Z�4���\���.l!�T�P?���,�	���;�*#fs�Ô���֠L�zV���t�������G ��{���oG���k�� �4<B�x�r(�kS�9M��h�k�T)L<�e7{�>
����v��H�5sb�=w{�y2��
_NÏ�;��&Ǐ�7x��rHx��o+�&����7��x�,�Η\*�ҥ���������$\8 }pBtwc=u7�
d�~�	����/�pΜ�G��D^�40�ɰKo~�Jfɦ;���R��>�&g%���b���Bt�Y�ִ���T���C�XH�%��Y�|钅�tp���o��TB8�oDᰄfن�x\�-UC��ґ16�w�� �=S��yc^K��{cv`������μ����`��D������U�o���!�L:D��D�m +D��w��ij�E1x�aG�ǯ�2f҃εP�����B6/=�+ӀD�p�|��}=���©��� X��y���#H�)���H��B�f��{Ya;l��:C�RGGr�}��������*�����c��c�kX�}����D��WT�K=a?@NA���N�&��ͣ��O��sAb�m��0?���E�GOel'Е��L�f�o����i�l��M��"����>%d����(�Kx
�zc���E�[���L��KL��?wP�!��������gy-���>�4fR�0%�������]���^G�\.៧m<�U�8�0�M�(6;F�|�E��5��ٳ"��/�wJ�H�x��s�Z�±᭩P�?��v�$ޗ�C�'ت%a�٠ؖ�t6��t!��=��'�Z�>�+�R�JS����ȡ�į�`���q�L�v�:��c�qJ>��t��W��(=��qʍ��R�%d��R3P��͌�$�Yc�ڤ�������ۄB�z����<Tx��0A�������	����|�dh7���.���QR�_����� Ϛ(�쓦8�o~��q?��f�,�:<�m�;��}ζ�M�vT��c9����A�������� )�H�@z�e��ԃ
!��k��0 7 ���rT=��v���)�r/DA�E��n��~TM��M��ArL�uV��\�%|g,��1T�4�c��(�҃�����.�bLkFuI�z΢^�9mN��g%$2Cu���Z���Wbc'\�Vm񌕾:3�>�d���>̌�i#m�Z��c���w=<��%���;}�)���@�ҫ���ܦ7��`�-u w���0��t>���4-z�K����f���s�;�ֿ�d�#�����A �T",Ł}r���$5'T�3�{�^�Ǵ��j
ֱݒt��s_X$�/哰���˚Dzi;O��áƆK�:j�a��	�M�ٖ��.y�i��<�1fܾ
�&-�+OH��E�pf7h�!�A#�|=Xɖ�H �Ī�:�"��hwZ�e�[^�p��,�1�w5�C��!#}�&��ÅY�#@�ꐚC�����F�9�Yȱ�E����g�21����t��;Ft�hX�&k�����ԣ_�2K9��m��|�e�Y���mD��P�e$���ߕ����x��`����,~�a�FS=��;����t[q�U��<�F�)k��|B����ão����+�<�j��Pᛮ��E�*<��t�ʿ���B�2;�|F��z�����\)�(�\� ��tG�S����|� +~�h��##۸��mu���k���M?)�|8���t��h��Q�@��#�w=ռ�/�5]�M�ҙ���|Xƽ���S�iRD����i��R��jXl<��L�@�������=�j-�\-��G��4�����"�!łV���޺�����ZoEc�6�<�O��:X�u�t���1� ��Z"����J�?�fU?i2�C��6:��zd�Z�;�6i�Q���/��w;��J,�ǉEs�������Dsڏ%Cc��y@7m��b.�8Ul�pB�#oV�W="2��{��E��7"�r1X^l��\���rm�<�h�yRj�6�����x��M��L�E�*wg��L�uV^҆*՘I{ù˸S%��P�p���Y��[pz�������T�/��ʺ�r��� ����`�LӸ��i���������{�I�},��}���K�ˍo������ ��Ht�"U�oG$A|��RmO2�����ɩ�,��%{;�c�l,ෳ��Z´34�f�6���$����+z"��Hq�P�?�y檤g=G��%�y�\{uO(�q�4*���{*��Rr�`cj����y��))=�Ԏ��Ƞ�2��s*���Ijrݲhp�ΝO�φ��(���� �iΖ�XS^�E!�������e`ȩ��.��[7xtej�����+��Ӆ
�ˊ:�W�%���K�l���[��@���W]�ϡ��X�[�;7p�*����c�'yzc�67�S#q'o� 7�,9�.��ð�ɦjIn��i?r�����$#$nK~N�~&M��U��7���jՒ��Uc?S�*�Y����j����v�u'�JU�@�D/�����E��E�H�����c0]�n^��ҽz���kc����������$�d���&5�}O�yU�P�;��y��OMn��=�|/㩿Ds��~ݍ�z9�!�'�ūxh��"�n��q�ư
Vc�z�)���Q��h�>�-G� D_�a��z�q����S(�l �,���9�׽�Q(�wo�Wuf����GM̱/�8 i7�������oE�o�h���;׵�lx�ӹ. ]]��Ʌ�¿�ӵ'�1&�T��3�w�kk=��Ѵ��*�;Xm@�]+h��6LA�l�N8xPN��i���IV�d����ނ���X�a�䧧yvq*�5����]-�Cۈ��@}6�*���0>�]��-+��=��=$]�hLC�i�Mk�������䬄}4��\�v����7�X�?�k�Fd�����׏�r��i��M[����6[��F�*��	 �]��BGH{���;��l�s)Q�1c���[I?]���@X�R�v���_H|=�ټ߷M�x;���3��,�dƃ�Ә����%p���&����E�c��A���'�|�)�C��Ԏ��NX�.��᎑�vnC."U����γ)�A&ң���\���8�����h~8�K�i�s氉�V�F%19���A�D�[����[�[���)�Q{Nl�*x!�	LoMi��;���H�bf���UY'�s}g �7s��l�Bv�� (��a����\|�gaD�z����g�|���@����l���E^��\^��h.�����A���ȍ؎���3��7֎z�r�3Pd`�����mM62X9]z�]�>�9TK��3L�E_O��i ��8�)���L��U���0ar��7�ө���v�����fc���`��M�J�x���N&�D�goY]&֚!�{L�nZ��!c	)�di�f�]ɹ��Y�=��J6Z��Z���ng�[����#�����o�J�X~Of����X�+pK�L��o��8�/�L'�$v,r�c~�='>��b*gSZ��������P/��7��*���鏴��1��1憓MM�����O�����μ�`Sp�-}q��$����sb��<�ߪ�wD�,c>y�M��Q|�R�m�/�[a��7���U�-�%���4�s4/6
����g亢��&�5g�;�0����� ���񏸗���0�w��A9E�Wf�4W+�k�g���>��0zv�!Go&�� ��Df2~�E�������n���������\R���\t����Ԟ�ԶhXO�1���p�Q��0� Yi��J�T�Wc�7�T�$#�5EՄ,���c�g*�[j/ �%�V~�8�~�\���f9�V��aj�&�"�XA���7�V�b���L�p�7v���C�z�/`#�ը.M����2F�M�oh�a��3^Uw!�>�y^��;��F.]#d 3�	��2�p�=���
��*���W6{\r�B���KE0����Y�>�ک �	M��@\��<�&i�x�W`��(��b��&�vi]sDko�I�rF�iw%��I����5�,.0���Z�W9�*�jo��� �w@�����WQ�MLݏ�!�I�9�s@�T���� 6�Ѥ�N��3��ϝ
D�����t�i_�$,&˯����t�f��s@��Gp^ �V���EO���=4��*!�r]�:z��E��y0aO��\N�[�=���U�Xf�F{"[4%o�["5�8~�_h���q7,k�A���tb:a9��s�k���˴�Cݰ�:+����u�ܰ�B^�Lc(��b��{,�ț��/�@��X��)OI����`���)N+����?F�fQf	L�����PfOX�4gy��􂒄�(�k#�M?��ZL'�P��B4�a���1����������F�>�/l�eZ�o.BU����  +-��l�Lg���Yc�+A���Å�����!N����!���X�q��f����qK5X,Wc�xՌ��k��7�u��o%Lf��yI�Br��~UF}.��.���~}c����V6�vn�~IρJ��������*��n����5e��{hb�9#46���@B�t)���e��b+��{[�k;��){����zcb�WĖ�K�J}>��h��g;���E��~�b�NJR�- �kn�.|�Y1��-T2�_+6�j��g�ç��;���|E3m�+�dM{)�>>&�FG�5�l�͔#��.��QԞͤ���+1UO�x�@G�Dv�@�l#pg:��v'"�%[�f�hC���@�ZOͪ�y��5����}ʬ�3PX5��: ��\_������2�,���6_� ץ��Dc��}n�jý��Eo��jy�H����`q��]������m���$�2m���py�1��Z��P��sy��zQ���jy�>�F��8�Il��ĕ��/��XE��(���i�0i���$���C��I��sD
X��w����f tw͐�)R<˟Y��zj�pm�v���YJ�V���(y� L#���>@,Ϳx��C6�VA�ȼm���3��M��{k��D���xx+"@2Ӓ���R�~E�*J�"�3Y�=�i}�"���F:�Ƙ$����L�[��י�����LF6]51>1��}9��iku�7u܌r�yv�G��Pn�55[�Ib�(�T�s:<̢�����"/����W8��0Өˢ8^ �:�g������E��翵�_qUbDN�E.S
^��:	���/-j(��h8A*7@�r�$j�v���K�����$��cP������]TT����I�U�\�A݉+�8�$�<uH��Q�o�
Cʎ��k$h�)�ٍ�Tz��ݡ+^���ڜ�~1�� .B�M<��\��Ѳqu�F��[�⹾�$�Q���DdU���7�衽���GF���(~��߶i������]����,�Gf:����*��� Ȓ!�JL%�Ѡ��M����xe���j��OR��nz�U���!�t�.�:&-H�����
C_�X��e"��aa�Dl.�2�1��"� jl�QOS]�ќqk�B�v�V�#?/��
�̊"o��te���*E+-��0a�3��7+��0��`�@��~����km<�Epտ���e�l ͵����x�����;��#�'�l�|�F&�W�pVWs;N���$z��FNc�Zٹ�&D�SD+��RNv�"~��'�����mt.A��pu���Q��� ��8�R/����(�蟏���W�t�ZP˦͙�>�D<�s�HY}q��m;�S$i_��X�v���s�I|Ǉ���:�k��J��ZŃ�/a&
L{�y��\�Ǜa�l����Tԩ���A����?��dUI��������onXa�f�uB�Z��y�U%������(���?"�h��4��U�[&!���.vk*{v���鬴^I��x!y\w;qhVBά5�F6���� *�����r�a���sI]G��9o8����J�xMh=,g2	�[�jl��ݞ�}��(�xό��� �Ua�e�#68YjO�>�n�]ɜ�w��^@<s�WA��@ÐCj.m��ѕ4��1cJ����4��2R�Z�}�w��I�T�L�==��s���駅��g] `DȘ��q�����#�=n�v��O�"\�i3��~	b��-�D�E���iu[�b�e��k�Ǥ�2�a?�߶���Л6�P�!�W��!Zᩑ$[ش�G��>��s�������"8�sE;��FM>����`�x3�D�!`�^�Gਲ�	�o��U�|�Ӌ�־�+��k*�)i#J������M��A?���ӊ�4w��QiѴ��;�Z��v�9����G|�\��H��
zޫ��sB�4�����k�PJ��Q�|���!�)���<iL88%���I��l�ZL�zx6H,	�h�r��͙��������j*�l�W��"�'�aL��bQ�@�s%L_�zI��P�����f��#jHR�a<�;&��hZˈGkC�ԅPT�me,�"�r8j�5kY�J��7/��q���r�1?(}��M��ê[]@C!���+g�G��y�ܭ�>����x�@���/p6���
�v����ܙ��l3�XHG'V�N��q�bl�V�S?&�?�5汲��Մ�(�|�am9N��A�7��f`�3Wړ�W�4�~W���g_S�� v��S�lk<����Ii4ތ�9y��*$��Є�]�;נJw�$tb�0�>�e�%N���\D�� ��O?XR؞d_сH^lo���<����s������tR�<��,�A�衟���/ ���|��۴�,��H���K&tMtK���vup=�l���e�$��퉲���ʻ��q��p�'��*�S3~@�[	�R�E1.�W�0���*t�B5H`��KZN�.F�]�1�XJ����?�� ��>�@#m6G��I����<j�$��%Jz��Z��_uZ`\��XO����6�z��l��4Ċ�{���3�ͼV��d+�A��W�i���Ě�	��+�����! ͭ�
jl6��=�4N���-�ث=��䍜�s�9��m��I3g>
�cX�\��IF���D
ĵ!�^�q�e-f(N0� ��ķO��D�1k�����/Yv��Ǖ�rS�r��ך:��h��pڥF#�h�h��h& $�٭N5��+��j9O�3%0�^(>��4�@��O��{��&���y ��e�H�������l�@��U?e�r��2<����\{��
��n	βt��\ݑZ���(>?4�N�dkW:�����-c� �d	dK����B�h��B���3���n�l��(3�8�ٌ:m�M�=��c����japE���oe�ɾl:b8sU���߼tǓ���Ʉ��E���o���}U9 >�XfM��5*����B��tz�&*�e�����<ex�A������$89�����{-�Y��I�_���!��U�^W=�|�.`���,�RK����G��x�5����>[���"JI��z@�%��G���d��iI��L�޺���-�.���j�&���e#j�"Hjti�􏑱�:��)��%Lîicmk~c���e������b�����th{Ͼ?q���`+&��܏��f�,{#R�}	��@��A�O�&�a�_��NP,)"�{.۝�B>]6����|��T�e����X;c�G�וAFnБq�ݳV�T�]��s���W4B�6��]N�`w���u����SŶ�Nq���<��|y�ܑ,�(�@���hZ�\NoR���E7=���D���8bA����cv@3S"?Q) 8?�-&��W,6��J��@����ބ#�n:%�u��^ﱴ��VE�$�m�C�lE���R����d�_*ӧ_��$5%5��@��G%�i3�"ATTWLT'b�B18�uM�u��b�n4�휓h�-����Hyr&��9a2 �T��I�֘Թ�ɱ��EJ'Uw�c:��3�A�7�}�.�ٖi �����⎴��8��N����I޷嫨k�R�>��%㉍��0N`E�]8������ 7��8�����DX���B%Բ�21�]�1��<A@�bl��v�E�Ti�����R�qȂ�U)�� ��<R¢T���`�x+�>䏬v�&}	�	�6��`�?�T*W����}�� ���G�ؽ��	��g�Hs̔�c�JE �)~�À��<N%Ψ_�;~�e�G�(bW<*m��Z�:G�� D��~'�-��\7h
�!&8�X۵���5��]�����T�.�u��x��� �|V[�%�	~t	�MU��^sRK�jj1� t悎r?m9k�����Z)ZC������	��z�&�g���L`K�G�>�_V���_��oFD��iKVu�)�}33��]�����擘�)����Q����Qc �u�"m��l�vH3��׽Ϲqj͢�[�G���r@���ت���!@27���R���&��՟u֡���	
C�Nl'J��Wq�(��@k����Cܑ�-/���H]��f�)_�W
���4=�rc/�!z
���ﬂ�j���]>w)�g�~�ӛ]C�Y��3����"p�i�!~�8�×+��֜�/""�&���s�
&ۀ�saPwic��;2?����KE(�5�Ka�h'�3c:��{���:�����!4���-}顤6jm0�\�̘�3�7q=�� ���.<�U��u6w�W�}ɼ�T���p���O�m�8ZX��0}/�$/�|�23{��rf|�C��˘**- p�.ad�\3w)�9��ӛ�ұ%�=WB3!_Ps�m�M*Q�g?
a_hG*3ZH��k�Z~VZ�Fn�H�ݽ��M f֍�X΢��M�2�o�Ӫ�ং�� ��_,?�!�:�"�G
6%I'IVʦ��,
I�p�iKu{��˫D6N��P��M����6���Ǫ yO/g������I�#���Y_5�V��4ՍM��	܋�~3["~?�B�j��Mh�}9%���R��FM��(��=�����J���2���o~fIE�$��8YP��塗<9�LCJ|/'\�-�����h@��'-�3���;���}�p�%V���^^A�(�y����ܤ_]�����H��C^@�fsB���į�|��fz3`g)�t6' 3ݗA�⼓E��0�S�����( ���3)����o�&����93�ϕ�݉�r��N�t�����;�;������Tp>�1-��:���Z�s�Uߙr��0��2����`ٍ!�;���&��I���-MF���DOR^D^�2C}���,*>u@&���ݳŠ��W�By��$e���cRK�i�(gy��-Ck�I9�B�^sh�������OKct���#�����9�*���R�s�(�!�U	u4�e�k����d.Ů��#��}���_aT��s�,P�(r���i��h� �h�}H0fgZk�#�ۋ��&���M��]N7}�0u�rx��.�y����!&�X��;G\����u�8T��$�@sXYgh�y4���-�<�2τ��"A"�Qr1R\�ul($���[={d2�{�F�/4��p�59�`H=�qK3镄���̒��y1�q��L�9+�M��hi���=���ӣtZa�Sv�(29c�|&����soРm�w�:�8;�Şj��y�=�����C%�[L,�N�(������.� A>��N���7x��<��[6��AC�l��"�~�ߐ�VS
Dd� ;�`��	i�$��-��xU� �/���,���@���>���^�P�p�EX��o�p�FZ��Ġ; �:H���m�8�m���C��;*ɩB�%��`v����i_��Ϲ�Cr��/]�X a��%|����و$�:���j��Wuko��@;��Sw�cM�,hңU�NV8�q��=�i&З��*�T+���Gf0kg�,F
�P�2�{��: ��y����> ��4T`�ń�E���T�e2�:���'��_�h���4Fׄ����(����9Z�h��|��.�����֩(��:AJ{�T��e1�?�C�,掱˯.#��Vi���_ >>�_��A�+EFݬ����`�c 1\��tJT�B�ӯi[7{�����v�H�q�D�*\�ul�q���b3��#\ i�W�E{�B(ە����G�jdϸ�/Q����P��y֛�#�z�+�WV?�|�ҙ��M#9�e�0ឺ�t�p�������_���
�Ժ�$�#����|c���_0�p��Ia�"��,��$�������ݒ,OPS�C�,�5��J�<P�r���#(x��5r�����} p#�Wue���� ������u� �l��-Y�r���Cv|��?�tXu�4\�F�q�� M� >�G��8��Rz�P�`Y8^ɥ�����R�6U�Hr��p�wj��5@b��m"��g�븰{
��Тe;r��͎��g��3l��M�#q�(��$&�nFX�� 4�`�U`�h���M|�	8U3|�X�Mk�Ni���%&V+�7t�n�HҊD$=�_���`ᅊ	 ����?Ěx)hyR��?����`6rr�E (i���j���D&�������7S�R�@�U�q�֍rOJ �{�s��VH͔��[�$��]���;L.Bۘe��Ͻ�L=��qC������4:��Y�_'���Kc���;�M
Gq��zmb��jS ��"ؗ���L���Ǜ��U�+����	�놾K)]bޝR���o�6�������՚����
�lf_�-�l�vI�xȀ�dKH8�t��/?���<�["�/�<D�ƔNh�u��tx(j'�����&n��3����94`�e��l��ھ-���Is��X��ؙA��=�"��f�S�ws5���}�� ����b)"y�\c<��l�������Of�zf�4í��{����7��^2l��������>M�����t�YY	��+Q��̻:����U[i;._OR��y��;lh��&�U�������ܑ	����#��q5\�9L����Mse��o�G��r/���������Ќ%�
8"�:�%�g�)���W��{ܽ�c���M���'v�������j��)��/��W�/���q^ߠ�-s��W�NG�gt��Ĺs6��@?�?�Bs��Kk����� .� 0�Ng���s�BD��Ww_�둧X�$��'{���d�R�זl<lڜM�h�f��x�!��ֿВj�0� w�$����H�1���R]׼]%��ϔ��4��������[M�c-�L�|Rk7�#�X��;�i��{P���8�DDP�鉋�c��vף�s�؛�����e��0V]Y�����N���S=5��r<�F�V�%��Π��)O�jz��[80��s� !�L����R�a/��R�x�i�ąU��{�J8����� bZ������Ǜ��?7��>_��r�'^������f*���%�5d6���[��V�+_��Ӷ᨞.���Dί2��t�0�Ży�I|�е�.i�\�4:��%$
n@�ԟw���u��]�f:��~�d�{��[�A���z��b�S`E�w� �aWw��?�Ou��A�P�� '�'��}�Q�R"�8t�+Г�x��K��,�b��q���s�3�9�;źa�O�/����I�~S�8"�y(��y3'�j^���=���+ /e�q�L��b�T���,�x^�6��A���a7��>�|Lp����6�~����`�kp�ךE*� ��u쫁�n��(���6�E��5	��w��NГ<���(�Ȧ%�M5̥\|4��ku,�k�ض�E���WOd�yf6������	���dZ&�kV��� s�~2�neI���O�Z�:pY�����W#�]�`
�y�O�+�����ȼeB�c;�i5���qU^��P����HM�L!3�3 ��*P:!��sX� �l.]J���ug�h�ٗu�ep�a����k���\/�Sq좀�eml�b�x�<���-�X����i��iՎU=D��9�a�PA��V�>F���	����E^&�8	9����5BfD���Z��t�`���t�C�*��Ͽ����F���C]�u��j{GY�e�Z=�@'�R�J��Y��.3��3���iE�a�MA���C��U�0�!u��� U0��;|�?ic���`���  �4-�zq���h�&o��MJ������۔rg1F��h��7�@ӹVJם?��[����gh�6����q�'RB������*O�wh��<�Q<G��Y��R*x`�|M릴�������51�;�3��on�H�d���>�nZ��Ĳ36ب\/��8��L�F[k� �Æ4��4��M�
��vLw�J�����#q�x�<��O��G���V���I��'�%�qL��n��|�oun:���a��g7�KM��I��لJ��2H��w��������2��%��q��	7S)��%!�nŏb�\ω|U�%iv��L�O^����E |�qf"�`4�m�1ͤ�@,_������s�8�=U�tP��Q�c?�����]���M�}��G�-��lW�_?W�W����,��^����B��t���c1{"\�ȕ������f^u�y��:`�$8k��c/�fԲ��k���̄o�A=#��xh��L������>7"��?�J�p��R$�Q-p����������@�%v��L&:�{;"Kܛ{�VG&��=��U�Ph�L��R��,��B/�-����uCGi�� 1+��^�T�c�F���R��:��"��Y��ӮӁ\O7��mzybn���=9��L�t�qq�h�uۨ8Z��+{X
�S�(`��2�Z�j�:EC�K��{�Sݩ�t��FM��pg��&@9Tخ0�W�T+/�͹���0g���w
FI�.�λjKY�Sk�e��+��4ʣ���WZ<��9q���'BI�^�9�467�I�{��2Ef�O��/]upgO�%ss��(��6b�X�,6i�����$�f�c�u�yl����r�&n3��y�)�k�&�{u�|�V����b�c���
1!~S�ˈ�! ;���Ҧ�R_�N�4'�\W}h1p3� �so��/v�Y?�!j���>cpK�4���g��-N��~�/uS�?��l�"�e#�5Ɠ��T�Ax�i��G"�x#������{��?��I��s������r���ހNk$�K�̘S�d���
4MX:�n������7�:<,zc���Vn_ mگ�}����\k��@�2�P	�~ x�B�q�	�S�ӑ��Æ� ��~��ʠ�:HY"CϏ~!ke��KY���N���G�}�����ʞ����e���a���W�� ,�A]���hк���@�t��/�.ߘ \<���r�` �G�c=���o�]�4�	�����xf|����d�Ǚ�𘲶�&~�fݭ���A�]}��=I�����|?�"'iT���	�'Mtץ� �0���K#C���bE~�g3y7rU>����T�v�ɍ>����p�V��=`����8*�� -���]w[{�q�����T�괇8��5���24�Кh��� I�%�<�uC�|wS��mH���{��9pH��~����E�� [��v���^VH:s�.�h�CV�п�XF�vh,��D���<�U�� W<^�ߤC�G��Y����������� �`�����[�����gf%^���ډ-��hc`��'@��;�R�Ӫx)x��=䊰�%_�m8���[iէ��%��+@�o�.]6�v�-�+�F�f�ye�I��M+$���~�J���'���{�%�X��K	��d6U�m]IC��Mi/F\|�,Z� !���ek�B�)�R,9�ʻ>Z[�6f�o�-��N �2{�=3+��.��}A� �Y"�̥��_h���,�>��.-���T�mK���|x�Bn�e�*>%�.�Wn$V�s�C�[e�����)^cL����QNI� *�Ք2rάdl��"�'d���Tߞ�o�f�J0�gye!٩'O���6~����_ܷe.�ϰ���6ɋ|f?���;B�ɯ6n+ |ƞ^i~�5��T�����ʵϊ�>?<�9U����*�rĊ�U��M`�Z[��{�����*H=TTC�%�QS,dAe?"^L9��r���_@��s��pN��v���k��}��	�r�t��jN��5�*�tK� ��w��S�����V����r/%r�ki��v ��5��A��LD'��K�ˤ޺��gA�Fo��gj�@�ry��
�1Ê9��tw�;�S� �)/�̭N�<yB�f>�O�X�I�mT;��#6����h�p��y���8�(;n�1Π��$Y�
�X��믉7��J�0ʷSB�̉mcO��ѻ_�br�A�_s0���L�B�VU،�l�O��,T�W���~���3������Sq�|�F&p\����\��a����4�;���e���/���*��8�o�$g��%2ݧ`[▃�a�y��+�}�7�u��\γ�[�d��t';� �1��QEz�i�(g�hI�U/�~>a�mO���������X��5Miek�>�Cm��M�;+R՞�J,	o!�s*Eh�!�y)� I�����T^�ʟڕ`+�FΦI�1"�iy�3����ݟ}܇�O� o��F��$��/�����i{A��H�&�e�:`��^J��T�]C����7����ze��%"U둬*�K����
Tm�E�#���h�V�t�e��]�VC^ioc/
�!+���+�5���/�-�Y
�a�J	z w���?0���� ����{!��[�bB�F.�e6Z�$*
�y5�O�J�s�d�.���G�����2�(��,�Ю�)r��={�����3��d���jI�����&�p��~B�${��6c0N:���Ĳ���w�#�����5L���Pǎ�9�ꌣH[a�°=�Db��L&��1�lU��{!��7�ֱ¸<�d�h���^�2&��Ivd;|��� "c�6+����?��gn�I̫��Y)��ަj��:8�+�N;Μqp�m#����/����R�Xg�*�TB�[�äj>`& t 1Q�x�39=~0ٵM��A�����Drc�����{y�z_��OݖC���4P��ާ�-<m	���qYх���r����<��%�BZ٦Vq0� _R@�T"םj�Z�_<[�.˰'��?Ď�K���>h�$d�*��\ۈ�y�E�=~�\^%o����5��$b���%H��H�75�0_>��H��ȱ�	gQ��!"��r�M!1�)Ke��M�G9b^��֭K��.���^�3�U�$�������7=ٟ� �?��5!���Tm��K�������0#�cXd׬�6��ǥI�=A��-�ܘx���<~���q�\�EwF�Q�f�5��^�q����@�]���.��#X��f�;�/(��j�gi}��,���[so�s:(QC��1���4?�����*>���X���R�����J�~=������^�Wˠ��\�=G���������nϯ���\���}�%�,��kY�u(E�<�&���s *��8��MN`�b�/=�!P��pM�,|_��uL�aݍe994�s{S5Z��f�#�O��Ղ���9"i���r�h@t�S�҈�@��ңn9�EO���(���t������w4C�	��(��F3e�vh��;�jE/ElWa`J�������c2*���M�U���KA�
������$��kc%2�Xs���18����b�e�o���8�A����.�o����祥K�N�D6p�`i���M���5;�Z��eR��ө�is~r���I�v���'��x�X%?��c�Y=�	}���#	8��V9�����k��(tSG�L��m^�v[+��gU���NC��
����Oq{����-����4��6ć��;Y�,d����1}�s��%�a�)%�k(�|c�7穟g�jjsDZ˥V�D���E�,�ݣ�Gu�bO^
-/6S�=Jc!ߪG������T�ܥ�4�Ċ�6Ŗ3>=�*^(�r�%?�ߥ}Q2�s'Ξ�n"b���=I����:�KYX�'�`�c�8�)�fG��e8o�/Wً�����	���&d�D1)�Pd�Н�}Q��>�������`�D�\-z���9Jp@�����}I8`�_�l�@���20��X0��u�Osl���,q	�
�C�A�#��U��M}�Iq�Z�u�q�ʶy����㡏�z@?j��xR'=Ϻ/A�Ó4w��T�����Y6@@4�z��p�W��;<<:E'w��r�ݨ\�h�:�cI�.P>����?�5��T�����u�$g�N괞��h���� l�W�=�@_�}Ԓ��>���$S�_W�F7���͍H�xS��%�����a�!z�Q!�������v^} ��H��?��6��8_����)�|��v\2@��5���ޢ�F�E�T��8dQ\���:�����Y�"1Ҿ�mv��s�F�2B-v~.NL.y_%��Ϟ�`.f�JF���eg��5���!��1�AP�Cy�ц _0����>�M*pԑ>=|| �U�5ed���'6B?��� ���;d��,�O>R���%sTi�|;SR{Ux���6?�g`��Xq��ؽR����������b�SL������Ƕ����b�hy�2��B���|���6P��y�{�2��׽2Q��6�� H�/��4�A��͟���I��9��ijH�g�&R=�q��I��� �b*��w�!q�d�lB[ �4N��|*�ki_�sI=�3i�8`(���૖��,���t s�$��v�~+Kux���c�l�~!6�5�����Q(�B��e7�	�/M�����a�?�Xb1Fm�M�.�p	P7��΄��ۆ
��5J]$�&��}Z�$z�v4���R���a��]W<O�<n�� cL� �,�,�L4�hJ΂�5{/�XmRuAζ����B���;�xfI�v�9G����،�:���̕^&H\Xu2M���L�.�G��ل.~��꧃3���:�U6�J]��l�t��ɪ��$cerMP� Q�̘2�'n=I����K�%���[l9�紙D��F�1z�VZ��Z���6�#=��'Ǝ���(-(?�cM�ՒN�Mi>�	�U�1`XC�o�I��J�Й1-�W��,g$P�kP�����1��9Z�vX4�[��M�p�`���ڃ��\��zG�]��5���p�4�Go�A�)�`B����*�pf���\H��0�dH�����q�k=֐V�B4T�9FؐΖ
����Wy��qL� �l�r�4�@���{1i�����K��~��	=ő�By���Q�r=r�<�����,j�5Ko5ߴ%Ae߶���v�ޙS���g#�o^�O��� C/�H)��2թ�����%�q�y��������V>���e_K_@ާ&���e��xjS���63�zS����+��֒��>�rˏ��}���w��V�������J� 5A��v2,A��Nڠ�=P��FpI���ܾc�n^If;�9�K)�kӒ����\@�׊�E��_K�}�a�z^�ԇ���f&P!)�]Rt�'P�m��':K*���-��V���A;\TI�Y���|�G.�����R`f��Q^�±�56���/
����a�H���o�(���B�W���j	s�[��cKt6.�q	!�
a��P�Wa#����NT�ŗA8Xz�����T>��Al�c?{�Ŀn�Z����i�c�=}�;N����~�.V�g �~Q@F�&WJ��Q��!2�����AW;��y *�_�u
�	�z�Q��}�[��E"K$$*'�c��"��˞�eoOG��(���_a��{��Xvca8�<}}bߣ��8�QM�m�q�Q�~��Y#���~��jS�0�nb�VG�M�Δ�F?�A�ף ��YLU�A�|x��?�m�D��	]D��	�����]a��g_Ii��zﺝA��Y���`��QpݸbޯZX{ ž̧,�}���P&�M�f�)����>(���W/��k�gʫ���.[�/��%m������� {Hی����N�(���i����պ�r���ؚ qD�ҙ�*`��D<.��]׈�2&�:t2$�s�H�є�f����?��>A�*>��;.�]o��5������x�a<؞�6 h������ ���[6�b��a�e���_��:��D��b��DHz�#�0�Wm(��y�ѱCD��-�,�Ց�h��P����K,��Q?��T�e�,,+�lGSd>��xI��EM
�i�_���<�t���q}52��W��~u��;���eE)��T�����Z���]��e&�
�5|ZqK"�����Y�f��-���up!��30h�%�=-?s�T���"x�Mz�G�L�QB�n�9d2N��N���_��8��;����J�.�}9�UF�>�^*>�h#8��Iہlΰŋ����/��g�B��	�93���cv:.]��I���%H��w����.���6�`�͡���/LU�;���i��QZ_D$w4ւ���[�aX�gԥ:B6�C��bk�.��VDA������v�W��#5���}���o_�I�ݘ(E��2e��O�g����9m�^�/ż��x�?�T�7l/
�L���s�y�A��\PəS2�m�4).?�C�A󙇭8�^�9mc�+����Gs�ش�!��C��8���� в�C.f�<&����}�T���l��{�y���30n^��Qa�Ҳ7ǚ%����'���a�9 ���7���6��t^֔'l������\�n,K1���ɜ�nAvHaٻ C��z>:��S�Ѧ>6v`J�hw��L+ṽ� �yz�e)	�Ѭ �EP�����U�����{��Lb���R��4h&�6�0}&-|~�j#����b�o%q_x	��Ń�bw;�l�]�3��?��[g.�I��������u�a��O
b>�/l@Va��+���-��E��þ����4���q�Z��KnE�ӽ�?SR�!(6���B��ٰ��²��~�=p9r �֑';�j��B�+?�63�"�hT:V99�W�Q�s&G��ӼJ�.�
>Y��EsP���.A�لs�Z�mֈ�g�
��9��Iec���CF��F���(5��V#�܃�f��^h6��r����_)X?�њ����4z�i9�Lf�֓�@��*TM�'Ԍ�w�������A� <��9
VQ����H�>���C�����<p��j�Д��O��0���h��a���=%�˨�5.�f���:1�Z7�?oi;d��1���3�Q�{d����^�-�	�k��PW(��y�Yk��>�o�☌�d�W�j�<(����Η!+ Q7�p�鑗]���%a�0�]���b�ݎqG�QZX��,���T!���&
\��l�xQ�ZM�4z����������Y�㍣���#!��5�îPb��L�rZ��KH�(�nCid}P)�I/�EjK��O����4��_��& L����)���p3ҪL�i!>Y�b꼙�QV�gd���,
_Y�i�D����&vꆜܐ4BB�)�0�ԙ\X��V��nuy��jFV�GHZ��W�U�&lN�����K}%P��8y�DR-&�wY��88�W��hgR��Ǻ��"��״�vAړYV�������˱�0�x4AG@+~z|��y����qP"[����h��p/������u	z�?;ﶽ�Y��Vo'�����̵6�����@�b{�M��ꔬ�U�՘�.��|�a��8�%.*+��2�"�!�x����/��{�"i�S���[��ʫ��	�L)XL�S�C-��WC�&��wL��?Zn��`T8c��{�$���=�ˣ�Ȓ�EB/�M�1������{E7_[� 
B���%�:[^�՝V��X��Dq��+�]�~�Oj���.�z�Mg����c�c+�x�U(_��&Fz�"`���4�r�#��HGN���N�W�CK���v�FM2��eR11�^x�&�����g�a�Έ�aëࠀŽ����E����-�ң�@��ݤ���Z)~m��.����$6)7I*$��</ܿ��ԅ9� `��"̚�1�9"O]?�j�O�L�K�r�4�L����.T���m���%ϟ�xL7�:�����������Qc������y�,�њ<����V�l �Q�ur�]�����þ�P�x.��sZ���&ʳ�ꚉ�)m�3nk4�Ra�e7�x�S4��`�Dm���:鶑*ka�7� ��SY�s���8)�C!f!"���6�ļf)W�~��,�G�_���\j�<3m���j:���Q��z�$j�t'J��������`�e�$R�D�|�!,E�3�覟I�
�
�2}��/z���u4;���ydC�Ɣ�7����^R��)%����<���h�7b�D�K-��ͩd�,� �Z��ڍZ��M$50�}�,����z��b%}˓�1�@��������IE���F�f^���`����ܻ7�F��e��gq-Cø��M�r�z��_��Q�J��ؙB&'9�������@%	q�c૙��)�t�����`h7� ������˩�%��J�d�!���\GP816X�ZGaq%��M�$�h���9�J%�2ς��T��h�o�@��w�a��fӼ�mxx�I�r|:�C�N���@�)��k9s��t��2��4����d�@�co�Y��!���r.��J�#8�:�n��&=��<��eF��'-�R����{H�|Su��)6|���nأ����]��702}K8�3�u�2���/�
�����`Ҟ�l5����w�� �\�k�^�
�<�r\`���I{��oΠ��Y�[�|Ѻ0~ ?��]h��bE฽l��ّ�j��I���
�֡�$��\�s\���>6��K1�2
�d>Ua��v�L�\����6�
F�?1]A���v��4Ș؍hx^�M� ��ri ��_]��}߭��r�d>��y��J��2��ڔ��Ave�˞���f����zڟ2c��Ye��1�vd��L�랅&!��(��%�ȯ�-��@4���EX~��g�w%��%6H��Y;)�%IOsI����{�p�	�Rg�A��R����1�$�pÆ	 .������@��l��9�!�S�5����fH�u.M~K��cjR�V�e@�t�ú���ӵ�ß��Z>�Y��On`�����h|�ۿ�I�����<1��i"�\<U��+w��@�䫔��M���z|���6έX�$;�sɫ���Dv0t�f���O�6�)V<N�dE��}��M�#�w�|TPgl�-�V����%�t�{:b���p )cW�=�b0�.L�)�k�bW��˵÷�*+�lqX��;���@$��W��K��H�v:K�bu� `J�=���Pat�G��g+5/o=#T��]y:�#���<Z�]�F�(���9��ȟ�,�+O�'ĎGh�����O��"3�*�=SL\�cKlh�Ե?`�����nŦ�B����Վ�����J�qv�JԮN=YGjd�g��.��Q����d�#7��L�kv��5��6z<�����ը����>*w���MI�q$�� �����B�_Uz=6Fg�<
L�4�ϋ@U�),�H�v�a�7�#��2\���aTHz"&ߦ������I�@���[��+�%+�9�/?7�{�e՘����=Z.ͨd�D�3���lJz"R�=m��{ޅz5��P�����5����;�˳�
�3����<�SB�G�����3�����<˂0¬*hM1RHk���3at����+��#zӧuD�N�]�/a�0C >(O�J�������d[���X*��PG�c��C�ǲX��nn�E�ح�3f*�.�s9��A3�OF];@]�? �e��93�c�Ij�}cL��w�s3�T�o�<��k�M�3B���� �,���O���nz4vh��s3`�'K9mpD��a�b7�����Gb� :���W+.ȭ�E.���ʆ�?�$}�L������Y"&�xG}�� 7R�ٿ�fg�N��:����<�2w'�mr���y�^�H��c2y���$�O��P�aC�w��˕E�T�Ǌ�	���5G��_��ɉ�8g�H��)g}z�mdzy�����pCn�V�|1�?C�7��As\��皾z�=��lw|e��
U�.DaDu���1�z�t�Zcg��R��;�����x?�^J�Z�"3��f�y��o3U[d.��\��{c��s��u�`�,�.x����Dy�˙���|�D�S�P��t���z��:Qxnx� FN)�6��u�2���>Σɔ����K�M~�};���L��ӷF�!D�4@v\�F�\�����Ո�a`�A���T��%��JQŋ��ӟ�L?+��]?ëm�{P�2�%lW��Vf�8@ZA�|
�W.��\O� ����*���lO�y�y�2�q��*����R<�HS������p������� -�To�9䚚5N��blH�!�B��?���TZ!���;|�\��g�}�u%��崎�!�<e�J~o��cU�2��*��� ٭�ZW���p�Ah�J���>���`�uS�C]^uz��AF*�D~yb:��ľ�9qah���T�z�C�uN�=�����2&�@�z]���w��_�~'<O�d"��|�z*~7"f��A_��@`0��D����!k�s}z�F�P4	U̽���j��gR�������b�%J��Cpn:g��y�aHo�0�	�[j�<�]�_�|V�v���nY���~j���g�Y);{qܵ�WL��1\[f��h�����IAg���	m婂I��P4��+\�62aC.,=�{�z}�zJ�w_A��WR{S7�-oڜ��K��W��\A���pe��v9�WX��f�������J�X"�5��X���B��V׾��?�f�����'�t�=��yP�AP�♢s����osh4~O�D��t1����0}�^����O˨�}nً�Δ�Kp��r���I���r�������.��_g�q�i=+el�d�7��	��$B�HЕ����.�"Դ��u���s1�K3���&�����n'���/�E|Xa''9_?chڧ��ڱ$͝c쥪M��~�m�:���f�P�&��J�����ƛٯ&z>�1Ү!��)6��T�}�̫�a	�	�\�B�n�T�Ӟo*�=����8�w�b����!�N�ڔD�{Au0W:���?wW<O�_�RK��薹F�+�`r�"|��H�B�cDd~���fS�6�B��ה\�3�K�ǵK�{�'<�v%�KJR4��?*���gp�]��J�2���M̈́և��7ZCg��q�I��wW��k&�x�6�	�<�ߠ}�u5[r�'s��4ؒBJ���R�����	%�1db<��
3���}�P�G��2�#�ql�Pеbg�ſ�:��'��R]�֧�1��R�1��et]����r�PY��@ï�+�Q� �5?�6~	�)Q.7Z`'�2��CM�����M�_��c I9�R���p�R�~�Dl���\�N���¯���E*ߎ�|]�0p��"s��)iKG���A]�XOr���Hf˘���iB-��,������,o1� ���U�Aq�����k�/[[ȃ�ܒf[�<;�C��Fպi{ؤd^;�&��
��%4X���F��>��n�[�g\�B�[��^w�+�!�ԏ+Ǘe͝P��B%FC�E�c¿
7]
n��à�N��C�4�d-��k���t�p�0��eV��2���	_�<�HD�{Npڼ/5������_e�$3��Ym��#���׭���i*˲e7$_fgG�$λ��%��W��h�-��yt��P��o�!���|�A�=��ݍ��wcH�^�m�g�X M>8O������"Qӡ"�~{��$�����Rl����a���>����ev�O̚�.	K���]�<�� �2��%�?��n|ɬ�v��:b�T�Y��$$=���p��ݡQ�!��zK<�~Z��R'<��j��𕃨��e#؄!##N��_�r<g�Y��"	ςT9ՙ�h7�Y��·�S��]'~sI4���쁊?��4���3'"�t�e�`]"Hbvg\��]����6���R'���$��`OG�m�����9O��B|�B�L)�$�q�'S�M��=Igf�c�^�U/��;> D!�7}8�>{@�	L���^%�)�.{�&�|�'��#��j��{1��,)ǴR�zc
=��}��u4��O�'�����i7�K�F)��`!#�\k�l���O�m}D
�`
�<;a�AOS p���Q�7�˜�~捽��d��=aH*8I������dsț�}�l�N�5�V��/K�,��_� X�ג��o:Xv�zY��-�f@��u]ꞖCI�]�ߚ'D�4���S�ob��H�SìI�)Bܱ+ѝΊ�Ժ��/@��B�7ڌ�~�*m���3"����b�뺅��(�*PK���(�M�sUQ���$�2�.�Ś�S��HU���Co�Ģ�^�	�"��쁻��-��t}���_cV�l���xұ;*dn'
��{�kC�r=|����bh����n3U��&�RRY�Y3�g:~�a?�X$^�R86.�m�����T�ɧ�� �����W{�%��/�����7t>[+�,�@�}���m�%���Dk�lZ˂�Z�m�}��r7-��AH��#�ڗh3N3���G�-2��(��[j��BV��9�i�=�)�1���jN��8�ɤ��2 	�$�݁�A�4v�1����@��՟+qap'�5t�b�j*����wd����&��J� ǔ�s#�Q
�D/������B���ޓ���{a��<2	|n��)�1[6H;��;��8�\���Y���w&��	����Z9�����O9�x�W�u�u1�]7w��x&,V(٣B��G�G���6�7N(�2s	z��F�3z9�A�I��� $��&w��Mž��xF`vp��(�L�4��e�!��W�Z��6;s!`��#���G�=QqC�w@�8�_���Fm�U��Tt^�*��T�j]":˅���k%	��a)a�r��Zٟ4�Pg�5�%�)�?VYt��C�j�O*��#:���m4�P����Bs�4�<'�6��Uy��U$�x���⿞V�B}ʡ�7�]e=� *l%+/�����K� Ą��?M��t�D3j�ք�s��,8_bY;��]rb����+�K}�8�W��3��	�x�Q����w�9����+��,�@P�QI���r0E��[F�OD��s8jf:]'_&��K���9+��o�B0-���gƶK�]�1�Sh+̸	�o�������0G�"�x��]��Zo�l�فs2�����z<���=���ӗ�c�RN�l8/V�!8C��ɰ�F7�b�r���p��/oNS��+� �Ӳ�y��X�d�\�At���uA�3ڝ�:X�v��-���-e�������P<����4�(��(K���w%٥B��;Z(�l�M�
 �b@�Ab�}��:Ŭ"�|Me$��K.v��2g������C�^X>Y&�5H�1��u4�GHxq^"��%�����k2R5Z��`��f���5��N��QKZǅBJ�Ġ����Eږ�����ǻ�~�(Vcn�E���7CB�����^.��!�I؈<5(z�Z��w��.aT�Ԃ3��~��l��,�$y�����y�xU�o�d\���q���V+�W���&�����n��m!���ܪ�иx7i�2L�Ù����=�A�����6Sb���1�bR�i��dv�=�NϤq�yc�ᯤ�`�:�	*�Z�E��s���юQ�p3��4��m�͓���\aٳ۹�A�#X�F�aج�M��]�)`�K�^�~�c8X��d��� ���0"�D-�ɶ���߶��%��ʘ�%��h�+`$�-U��'��㙘�r���-�Q��FM�8��]boA:��Z�,-j����(�w�l~�2��� >�Sʺ�Ѝ�	��epx�O���3�����BY�wQ-��S����� b!¹����%IO�3-��+"(�W6J6��6zn�����������[V{^t���(��B�D���/�}1w+@?3/�l3֫��b��\7L�r}�c�;�����e��>�[����N9ԕ3'9�N0�ݻ��t�э
�S6)�����4���M�cb�E҉���K����ۋk��� W�Ȁ�>ʵT��T�`˽?tV�C�l��{"�d��d7rE��t
�ȋA<?��h1�7�*$s��'��
�Fk 9Qr�_��0;nH��9����(�F3��Z�Γ{����C�%O:V�%3�Cw�$�_L�k�L%��fMԪ�'��{���	-��%�}Q�݈nt-�]��+��y�xov��b'02҆�)��^������|؝61�0Ƕ�ug�]*,\D�b3f�R?����}g�ݎ*f�I����$O$*�j�{���6����q�2��k��t��t@m{��Rb��~ȳ�!�##Ū=���K��d�:��	������=75���!�l��g��YQ%Q
_/nn9F�_�Sd��������Tަ'T��I���O�l�(���^$)曭V!���=aT'��jrV�L?x�uW� ��1��N,L�j�`��#{q�¢!G�j�?x�=�����I޺j�A�*�79�^�݌
���h�)�]����%���Pm!e�9ӗ^*設ǭTD&�uG����tynA�<�C9��p�N�L���	�2�d�FC|l�A?�=G���6�;H�⛹Æ7�C�z����8�3Oa���R;QGyi��z1byYq��Eo��t�id��$`A��B[uuRʬ���
���΋Y�����_G��n�Pp"��PA�3'�7\D���T�x���Z�ZUQ�P�h�B�_ `?k�<��Mk��_ ��0��ڨɨ=�z�A�Ȭ'X����sj6����o�h�}���3Z'���U��Ơ����MڍdMK���##��zg3��F?�2�D�8Y� �k1��߲=h9i�Mr��Vk�)k�d����'�T���&�%������]������[�.'�����H��&/�q����
g��rE���Dq���@J�ݤ�����dV�N`E/*�&xA����G����k�;s[p�L����F�������:�W'�Ũ7u��KU�h����h��� �������7�k��,�3�H��i�����[9'M���g��a�����y�ņ�}�U^�����A��h���ESl�M�c�Q�,��q �H�dElPko83��fP��O�q理Z�ջ?-tY{Bg?4-V뗠	
�d?���G�.F܉P��(��4p�2����龠2���*���hŵ ԔNSL�[�_Fw�{"�R��,6�������E�l~�pc:�ǜB�Y�~=� ����Ys?��g��w��!��Eg�١Eu��z�[�sn9�t�.���n�CxÂ�)/�gt�=Ǚ����8���6��k5:+��(�_��Z8�IIk��;e�'��T=��C<;6P�n��-���1�\�o��!�u��x3ԻB(�yR����k�| ���X�o<���4����mh���P^}'��i���Uw�����w}��3��-��&Ϸ��P�\�Zh��8���L��pg̗,D5��mIq/x���:�;�BAMQ�_܃1FH�&��,��y��cp�ܻ�N�k:Y��:��?�Գ��Ѻ jg3Ͼ+�O���^�$L�����4��O�x���Z�mg�|&� �/rJ�y�[WY�4VL;�V��XԳ�s/�� ��Ԟ6`���W�E�_���~�r�7�� ͛��|�D�{�l��M�X"NZ�P���������\
�}� �$�Q�A6ыiෑ
��s��e��<�ǒ"[gRJEw�h�|������C5�d�%���0�Igڅk�*_��UA���$~ �荈}QO]1F�GT�#��8dQ����Ah�vyi���W��'���CqGI�����%��<�~�E�������G�� .J��A|eTvP�
�X2�QN��i����=�B��/(%$9j��TTF6��K'0���^$�X!-��T�@�&.��k�!��l�7����0�K�q1���J+m�?:Og,�8V-fv�y,)k��k�.��@�ei���R@B������ϙ-	i�S���}���|
�x��T ��jb=A����lC��B{�J�O2����(��7���|�ul��\r*��HU��M�=��n�dP9.HW���v��� 2m@�� �$�6n�{w	�up�@x��ڀ��t�D�>�z�����+ ?�~`�2;1g�=�����}��HX�~���b����g�W�G����'����<��Q�Y����ޤ���"�/�BP��Ӝ�{�)�M,�(fox��	�Î�!���3כ�(vH����J)c	���эJs퀅%]P�?�١faM[y�s��*�l�����h>B�3h�
���ی��;-����)�;�qϖ�X�뒛[���D�5�!�Z�=O#7��k.Z�'k%�M[�1\�ħ�-4Z�Q��W����fzH�p���2B�S���ܽ<k��������Z�7���}|?�ǲY	��3r���r�z��SVݫӟ�JI�򐶐M4KA��6-c��IWp2vy �b!�}r���IT���tN�t�4���85���;�U�z�t`�S�y®��u�!G��^Yd0zBb9ˡ��v	"R�$`�o���o����|5��\�����;7"�#/��܌������T$�Q|(SX��J�)�2��w�"a�����̦
GסvB�:�i�١X���J���������$�G�b�،Q��ރxp�M�J'�V�Z��|�(������9Nc�e��b��BϕY�Ct|e�s�r�h��E{��b����,�� �Km� �׸Y���{U�7�1��~�.�����j�Xh���O=��[�';����(p�I��%���Ί�)lows*�~ډ��ә�+0�.���s�z`�T�DǇGo�W�m��d�h?q��s�R��]�	��n^�����K"k��\�o���J�(�b�.��ơ]�Ńk��<���0�n�[���6"��(�c	6��]E�eA7ś�Cr
ۿl��Q�XΣ`�O]���/�	��nFՈр;Z� ���s��#m�,E��TS��@GmK�eG{���!i���+S0eXd��v�a�|dd��-��
%�ye8�Ph�G0�H��A�K|�Q��Ԥ֏Y������%�u�t�g����G_δկ�'t�]��EB/>jwiP�a�6k�g��3��I3�ar<+LS�]�0niG��Tȣ�*;a�Q�i[o ����	�9�4�J��0�#��b?h�$j &���*�Z,"��ܳϏo��;h7��
ŶU0���?#���
�u��WWv
 
�eV�y=��a�������=��1kk���Ar�y����;�J���� 4���Π�E�#0��r��-A�9�8�E�>[��LwQ��%��c,
�֎�cI���	��(ˠ8�ĕj�	��"t���n��푈��3V<ܦ��r��1:T��|НPV�d;Cc��à`�ܭ��>D`����w.�薹eK6�19�*��v��ү����U,_(Fp���%�_�-���kv����i�����ƹQ�V�,�y2����Y�`�NϮ?"(����AXx�.J���gT܌B�ʡ�.�����u���^PV��t�7 �y�!G���U>�6j�}m�R�����v�̧du�jr�_�x��)ɀ��Ņ��@��a��}�N��'w�^�n��b�:yѾ:�=�bER�#
������Q������:d�֍�w�3=s�/�t��4��Ǫ�iɟ"�������]G�n3L�����[����c��e�J@�|=�����e)sk�̸L��>��6cLoY.�MC�㫑�/��+�����US����Q�E|Wy�5Zr����pF�,��\�`m�q�WƧ��V�)�9�H�Fd�(�+$� ��8]�_��nܳ-�,#mx]ط����{�v���B����im=~�ko�X�!$j�����.9���vq������p,���r{�t��ú���Va<*0�8�~)��u�],[��"�A�zF,:{���������a�q�A�_0�\�5[A)��kw9%�?5(7Y�+�U1n^^��_}Y4t$�/9�]H# Ǥ��aG��3��7��I,W(��t	�~ȹ�G����jPk�W��U8�@u��ZP���(�gBCY�V�1�0��­��, ��I�'R"X�;k] Y�)2�a߁D%挪���r���_$��PΜ��G��x�E�����0\������L�w�I<��wS�AM@]x��CE�����mHo�=�N��,���3�ٖl�7�Q�:h�$��q5�����6Mdv��y6�)R���D6�[gH$7�Zp�4_��~S��S��`����)��|+�vԛP�)X:���.�j ���R	�{��%0[��-+�N��Ȧ'�����a]*`bE�;��3P��(�XR�N��,N�by�3BJ�'�i�~�r�Ic������<YV����0��'a�qcx����*9�sRSe
���s*\9:s�>s������ ���'[�pFb��az�!!�e��K:�/�Y� ��ϨM1uĨ��0�?��e9�����u�w�1�ܜ�btd �mO�e巹y����.��O2v�f/�|,r{jp��0�1��k۝꼊QD�p��䙊����<I��Vܰ�!2-���߷�u䢉�Hx-��'�	e����a�<aX����W����#�T ��KP�;�G�!���xN{�ˍ���]+��Л�T��S�|l��;A�1�� s����p�O����f���������y6�{��(7�[�f���˚�#�O`�w����ٗ�v�+-�Z������?t��qV��FFvQfQm)i[P֫�:Ac:�S;�E�W��ԧ>�Yt�w$�c��%�d��zm�����IDۻ��n��!qRyݿfm#w��n�L���"�2Q��hcp�E|)��䷶��߆&E���Ըx���4��(B!�a������З�M'�e3��O��~\��#��$��+���R-wL��($7��.�;o�8����t�*��#'���0J����y:��P|��41FL]쑛Qc wQ��������3�� )���M�QWC�T�M�����f{�X�S�o��c��Ni�z�ȥO�).l�FΘ���2H�����s��`x&��b�V��$}��� ;d,8��Oh�5N��$M��,�i�<	�Ņ|��\����%�.��Y�i]�����A'샸u�%�O�3��ҵK��+��@]����N��J�/���HLz�n��3 ��㱻��0 ��i��ݡ�E�ҥ��Ez���.l�g�1Cw'œ�+ i�M�9��`��4��i�vנ��o��j��Q}���Ǡ=~���YP����YP�^ad�t:ڟ���CZr(#��+q9�_׋r:����r��[�*�b�4���_�DC����I��R!q���ˌc9�Pe/e�ft&I��$>F���J;d���FNNz��)��F�)v�!�����Ug	�Y���މt=��� �����-4�� �c�t,5�� f#��q��U��hu�z�u���dj��Z���5S�w��k��Eю�Ť+z�9[��N�=搙�;����D�m�i
 �z~��T=��a�!�!ط��6Ix�/l4�����>�0v�f��E�Ϳ2\��7� H0�Iz:�f� ��l%���ѩ��o�!%��\0[�1=����ů���O^�0��q���c�[���|�^*������Aʸ,6œ���QǤ?�|����-:�=y�H�N�_���#L8�������X؀�ؼbx·iY\���oO����j�95�r�r��-���!��f�$k�n�����D�����8pK�"�?�o���v��������9#�j[�l�$�V���Z�DE��O��I_h�A7����e�d�읡d��2&�T��������T[�ѼO/�m�m��m�C�Y�4J��W^�)3l��C/ɻ�鈑��H�E�T7_�����H5�jvSi��]u���a��GM��2ZU[����r	IX�0u�1����k��2�̓�	L6���C��yNh�#5�\��*�����@����f*�@��q�����%�0%y���s��\���8�@�X"�.�#H)0�f��L�Gb";W?T�I+s"T�T�(g���:�t����܀�EѪ��Oʯ�Fy������*���Zm4x{4���:	a>�V�*�������V����F��/xG��(pf~�)F�V0�Kv�˅���PiD]�F�`r�9��7~#% ���D�R�Z$���jי��$/�`�\�YV�l^v�/��6�ߜ$C���},W�@���D3�mA[�iH�zG�{1y�x|IN�!Y�^#	�;�9���W{^�TY ������W;}5����#!�azݘڕ*���Z�4����8K֭"dH��\&�����2ɨ�f�FO�wA�e���*Q�2��?U�����r�d&��K�~�?}w�M*4lxեh��=���P��=�OG��-�⸨��Z�R�/<��w��4��ר��>Z\�C�j��&�nY�Q��(��@*n�����&�|\�n���_#h���+���P����T�.����D��{��Q�J��c�Cf�5X�rЌ�5���?1���&E�4��x�Q������d{5G�|���q�Y��h"�ܛ��x�rK����q�P�a��7�oN��×\�xi���C�.��Xz���]�M�@^6T�~/$�uz����'��.����id��t9��V�����m��үƣ�0��T�{�A�iZاڼ٭[����o���T�{�]B	�SY���\����a�"xU�Ca��Ԓ��6DN.ݶ	.P@��v�pmMV�� ���;�}�������D���|Z���|���0O���g^Jk��_�v�:�m��U�҄�m-I�Ag����5[i�8Fp��Pp�I@v�RI��@��ƳVp�;��ď.h�kM
��'��c��w�9�i���"��@������~��ag�43��˶�P/|�5�b�OH��Ӌ]��}�;�G�A�O�_A�8���nE��K�6f���i�O�_���X!�:�ʆ
|#no�+Qd�3�7b�T����Ԥ��r��Oss���6�|6��'�=��6x��xB<�Aچ<+�*��{X�߯�xP�8B�M4P��&߆�f������v����d`�(<Y$��~�ã?E�4{�5 ]��;�!H��^��Pu��L��[����ӡ�P��V�$״��I�Me�&e�+��Рx�����cP1���]�G%����-��D"�HϷpj�A�J�Iv`��EƋDFdf(R/c�U�֔IZ_����Vh�!�ܘ�Y.���*��lE>`�L[����H�up7�;�7+�B9��W#�3M@]4�!A������$IK��齳��6^�}5d�U�l���Va^��?�2H9SY��2�c�nxU���a~2߇ws��8(]c�0r�5�a81��$�\�B�� <��`!f�E9|�D����Xm�N��7-⭥�8��x>4��%��Kn��c�@bzNd��:�g����c�	���ӗ��Jy����U�Be����?ӑ�mP���I�(���t��
�Χ!��c&=(���SoG���d�Y�Ng$��1V�3�D;]|��;��6���9���>����r s�z�qCzw��Ѣ�����6b��,#u�)޲T�����C��2W���lrу>��ɝ�K���1�2g�N�C{2	k�s�[��I��G�'�@������������r�������ظ�����ڝ���vA�[�4��������`3���k":2M���P�G�{�81�>�w��˝�x/RT����h� c�:�Ͼ���;R�#��"��*
��EI��͑9\�g�Awi�e���� �=2�"�Ꞻ�^DiJq'��`�r�>\jZ?�s׫��Y��a���ַI��jAa&(Av��ǜF�k({�Ԣ�;��}�'F9g�˰��E�NxC(��J����z���'1��M���+i�reE���_X��X��q*`T���X�����w�^�-�`���N%(k��<��q;5H���4�φ�(�e�Y!"n�1%�:`��v I:�wv˙l[����5����c��_��j�d���y.�i��u���a	�i�4���� ��<���$��%ٗ�(�,��H�+�GU`�oUXnً��x�O��rFs��+�߯��>@
Y��ϝ�:3j/�W>qe��x�Y+T-��[�����$`�T6��nj5���#�&^Q���D�a��9����O����c�����݂,>��eq�ň����Z]�)G����w��|h������j�lw��F}�R�3������y�J���I'Fb-�h}C�j��轍��Q����xupQش]��W�����1���_Ɓ�����`艴z����c�@��s��i��RW�1�AU��,5�� �}��#s�WS*p����%� ����2Q<�`η�xu�Ο=�`@Ku}���E���ٳ^b��8�����u���� @�J�k�N��lf�}�;Gٱnǩt��0�/�d�:`�W�iJ�Rw?�,+�BV�>�R����t�t�#O�.��+.��}0�9
h��y-�钗���4[�@e�F!+�����F6�Ut�7��@h�R��w5��{������L�o*_�)��OP|0��sᥨ�|\1`j�p�-]�=�+X:v�6�O03$
p�n���4%C�(�ɿ�^+*�b$��G&�Bc
��g�=S?�I/{y��6�~xi��8�p6�X�Q�<�GiX����o���Q������TT�-�w���]��<��m��TT�<�L�W�k��w8��W��i���o�
��f�{Z���)p홧i~�G����i�Ȁ��>`�O�9Ҙ�����x9�W��#�Ȋ<Eն�ӚӪ"�T�#�F}��;i��~�f��F���oj����멣��>,DάN�AE0�4����o̽�U`P,��b�<�>k[`6c!P�7��wa6� ko,��k�
�c�)��a05{����ybGj���R��rw���4z�"%w$U�J���D�,fVi����*	?���.<��Gi��t?e(�����:^����q �xm�?��t���&�y���kW�7	�r�m�Đ�W����Uԯ��f6��(_|�˅�A����B'R��y~��Q�'~�7	ſ��v�M�S�d�*����L���T�J^V���sg�';��c�39
��<�#���xEB� P�p����WLalS����?ǽ�����]�7�i�~��!?\
��s���	_�I�&����@�R�l��0�!���)���9>It�胞�hC���-��Y8����E�ف��a坢�~�@`�/R�d�4^�-?+��,e�K��G��������e����bR$V��|��K�:�h�=^T�b_���|�����=/�5'pYU��kX�� ��#PMx]�u��R�\��i��� �5��m����2��<�BGav��֚\|�,��s��c�l�q����s�6��S����j�d�>w}ҭW�����Iź�l���m�@c���b��^����H��R�~A�=RD��%�0Y�O�����z&��lz2����G@����i$f�'����FKE-�X�P�tC�!~�U{d����b�E�#�2�ήɠ/��KTҠ8�}fMT.r�j���}S�6I�O����%,S/����y"��R��+����G��&���v���)��$͔�3���~d
�����B�7��'��mn��L�e��1`G�$ڧ�����⊮	�i+��d,�\a�A������,�⒗x}ȹM���vE�Nve��J���0���+
�Hy(�%=��F0Mj�{߁�HQE���A�p��Bp]4�v����R�dI���F���*����83�ˮ]tG0.=��ۡ=⿫�2<�����@�5[G�=.�2����Z���aO�������)�Z��Be{@�?Q��\�̙��ūճ��0�7P�
NxU��P�� 4��$_�Nقo:e\sF�
���S��vU���;#
p��u���N�bD0;N��:X��[������;)�Y-��r[ě�;�(����3��e '��Y@�������V�[&�A�;�q��#�ә�Y_^��J��V�Q�M�#����M��P�:�\�	OH�����R���aN�]̍)�+��a3�MED�e#��&Mz��~��6�K7V�;L�֟���8���U��s�֑��e_f�#f�;]!�ʔ ��:5�)6�;n�K����+��~���o0fD8�ԃ[���F���S>K����y�@Īd�m�>����l�c"�+�q/E����H����ܓ)��/�����次�KkB�b�!�P5��iQ�E[x��`YkK�H�!0�r��x�������i�({�м�����Q��iۊ�ڹ
6[^�eb!���L%x��˞5�QK����ގѠT�=��dİR/���=�
q迠���m�&�jF����:qG{�y�K���v�[�m�F�%YE�T|�te��I�n)X��C/�7쥦!Q����_V�t�h�U���wg��J��PNL��0M ����� ��@���WE�Y�fWX���p@kd)M���� ]��[6 ���?�8���X�<U]]��E��f��6��d�[Iu�Nq�a�D�X����#�D޾�?J������7����Z�Ks�{��F�U3qU�[���~_�Q֒�mU���A)"dip���z4rV��wc�YV�Qx�YY�G!q�j� �7ơK�/~آ�'�:�!�����-9�?�o�q�7�vT�)C���4XX�F+�	����L�cVCd.X��F�N�a�l1��>ܤ�WE�}��'��b}2��1�1л���2_;�Z��B��o����հ�c��W��+I��ʰ1��₽�;=x_�ȥ�����b�am�[dK}ez6:pe�לM�-(Y֫8��f �a禎�:DE~�\=���+02�z,�7��H������Pj�G�O�0{TD���n�7-q.�kz����2Nwftȿ�}1_n�C�54�w�Pv濯/��\�O!�*�ҏТh@����Y�o��w��W���-��d��rA�ɉ��FC����6�N�ǥĐ�(V�xK6�G�����kf*Y`Q��$(��q�O?�nRG�mc-����EF�5�:[��L���n�	Ό(���~?.N`�jN�6�a�HHiu|Ӎ�U��u���=��1�"R;���CǕm��6Ԅ�)<,�ܡM�1���*<����n'�'��S�B��|���S\���4M�	�)��E$����z$>����T�^�� ����!��G�&�����<�dL�=g���pe
��`X��[v:Y��E��@�x?�w��E_���\6��*E�����M��i���T�{�1���H㡡7-��3�m��o��Cn��N���y.��$h���Yp�!��cs�a���H�2�ߤ>GH����}㩗���K;а����c�T�Ɲu�a덆P�#�Zu����æN.}���+Y�����~e�x���_�ץ�:>u ��(��o����`7bb��A�Ds[;�y��LN�����O��(9��G�0���������T�%����v���(��c�}����ހ�R����.�G��{�̟�O7W�s��L0�@��Yg@wX:(�<�qW �T�Â�3�Ty�!A�QU��$|�������	uY�o�&ɍ{+|_���X�=����ͳ;����i0#!Q/Qmj��z�����qC"e��5c�ΫƜ�����y�c9Rq����+���U>�G�e��e�����U�W�k%}}�kZ�U�c�6�x����s<7�t��r��Pc��f��ub�U3W��A���(7��V;!���~�~@�j�@�,�S���F�
?1�H�Z�!�|-���[�b�f� /�^$�芏�sT�Q�2->�zWtݯ����C�ڴ��>�z��a���z���ST)"%�7�R���V����`%7��`�D<5�(sq�[�e��`ЬM,?�[�qz�Ԩ����P2ѿ���%qg�#���g���������)�O��hF-�*�ȝ�v�~�h~^��k�c����l��uf�ת95x2��O�__Y;������RYB2-�{�G=^������h�;�2�GbZ��=Wh#��]Q�t
a���5�-ORY��n�"�K�ƛK��&��zg_)�
�2�bW��UE�;�c_���$5�v�ڕQ ��L���� ف-�3~��;g� +�[����0���}�����NR
�y1;O����8ص�;�@D������>$yv7��+���Q�8ѿ���c��u��\�� �h�`�ҳcԜ9���'l=v3��}�2��W�$�ͬ����oq0%��ZMA��3{��;F������(�d���Ӕ�W�z�����7t�t��HC�9���Z�*�C*����eS�8ٚ�lC�8d��D���iIX���(��8A�Hh9�YkJ�ek1P~��#�����ٰ�}���y���US
SY{�/L�a#&�%��i֑Ji�(�	;>~�"����;��5���OuV0c�M�7�87;-4�f]
�36x6\��@�i�p܋�fN�]F��+���ӟ��4����W���n%�V5�C�gJ=���q�.IX�-��2$��I�v�<L�73|T�k������Cw�$*:q>v�� �C]�j�ˤWD��#`*�x-5+="�Q{])�sg�����C5�������34Yx�+kY�����u�,Ji]���^���LS��kȔ�)<-�V!&9�FҞ�`����6B3�	�}��}�$���4�ӆ&v��#PgBǝS����#��˝�B����~BǑ�\�W�o��ԒL�姖Vs��$�Vd� ��Z�O*?  �	�a�������@!�0�;K��d`�� �X��5E��L�KS/,'G1KL�2ydt}�N'!ƀ �<�x�r6!�٘]�;����R.��8�4��U`�!3��gs���3�3=� S�댼����^3-mB֟��N˼Up���QA� ��`�d�pq�QӀk0D{��Ƶ<������*"�sn@���-4�pT �� h�x<�F[v��?_�jK�R �n��H`�fq[�rЂa	L��t���0o��7J���(�޺�T݉�W6�Z"H�F>��7�V=��U;���<W�6#�V��b"�Gu����q���GoE��}\�cA�UC��*��߁K� ,/*�k|�Q{��?�Z�n3Α�U�K�"�$/��M���&CH��!x7Y�퇄�Y�{'(Zg�UT��(�4�k̈�/a��Fa�UA3���d� ;do�?�[FAa�o����k����i���@�4�v;i�)J�R�67��\L���p��Mt
l��3��9��D�7��V�l��N�I.��c���� 8u��g�lM%��X�s+��N~�
{�k{�Y���kN41.F����O�WNӂj�˿g�}�4�{�=_hW�
�;*TV�S�sHRIY魽WWb(�Bd������Q�6H���_ɾ���ȥ+����(\)�g<a��U�2�A� v���)�dU�&�� �(���@�|"�ud��w�f�� ��r�?��WK��4��p`��y�� ��s�Z[�Q+�<�˖gs�~����!Q�ԚTx�ꖍJ&#�WCS�mo��P�mT��L)�@hGܲڲ��ԭ�w�G\�'��1�i,r�/�J2�/~K�%찄FH,��:WݬD�#쯼h�E�?^�$��^�Ȕqڝ!a�D��GӉ����M�#U�!r�|�=~v������HV%��r#1���~	��ݜ������34����K#�����G¢�֥�o���c�|�&6�ä	Ō���﵆���B��v[�EO����������m�+���y��1���K�b%+ʚ���*%�L�f�%���F��6���5ɸ0��!je{
+n�	~�~�(�Y�5۠H�a���(�wzh�<^Ң�b�.�k$�������&�!���l�z�-Y[20�X��"j���2t��Z��T�nq��T��eD�}Gb�
��}?n�/�����h���J�a�0����'��ÊXt"��c�O����)W�91<~�	�|��1]ʘjET�eQ҄=@����888���b�t�t|޺������man�z�I�g�56�E+����u�䃿<�Ekͭ� +��;os�� ��1��s.h��}���I �0){m%�YU6pSy��H�ް��r&M|^�53�O;�*��������ڇ5!o��hj�8�M����g�0�N��g�^G0��X�c���� �F���:�AaO��*?U^	v�xeu�Eni�����o,wDu��Wl�`Fy�5G+?�&���s.��(;�*XAđ�A��.�---��2�T���,��,��� -w��,�6
���A&q��t`B,����~V{�h=���'���#9QSs��� L��#g���	͇eUW�7�1���f��(�''�%^�-���_̷���3eB���1d.��-f
t�-�H~B�����b�/�O�%��w�Wը�����wR냛���]����?�щ�J��N.�����"9�9�7���6J��ܷ�\^�c2�x+���H���۲Y�C�������nN������yۦE����ks5��,��I�Kf�b_��	�i���km�AA�������p�)b/�Ӎ�烤����@{?��]��L2\ .ӏb�@�,~l$�݁x��Ts��S� |yW����G�J3"!w��T"�st�+�霁����ۆ��J��%�p���\/�j�hʞb���l���{+zwɥ[����RE�[v
vN-���k�����1 �7UK����r��;�|\�B���?�Ѝ���9|K�&�\xJ,7Jw9c%������)�)C�U���ܿ.�����!mx?̍��Zȗ~���b���R����	&����GJ�I�r"�2Cv�I>�5|R-n��P-�����?\�¬��2�:���m�buxL[�ڞ���>|C$7B�e ���1�4Qb��;A�V��������Pj���_��z���|�)s�����'<��߬,UT U��$�d���ϳ�&��!��`) q�E�ɕ�;}⨢�M�F��
@�����^���CH��d�O�Z|�J�V��-��M	��Rg5J�t��q_�k�B������K�����;��o*��97؄����AS)�Qh���֙���D��W��A(������g�wb�yY�@���U�žvv�5a4�����P|>�7D�E:mtI����WŹ�%<�H�n�e{�b"ô0�{s$[<��G�"���J��o�X	sH�l�S��ߏ�\�!�����?Z)w����fl������yet���Z�-ʷ�/뗊\�oQm�:�c=	�!��KT�ȱ�&t],r!b�X߫UP�	�5*�qvw��b�cH�3�颛(a!L�;�����WV`�0g���� �<��3L`�ɗ�u�iu7����
��}�r�W��t�+���(ߓWo�$b��'�W����4�4G1�Yr�j
><A�xU��F��FISZS�ض�q.ܖo&;3�w=�(&���Z������T����0a�H���Km�y���I
G{>�7Hnc�%����f�S; _4���M3]�D� ��T���]��+[���	��_I�q&����b�#zU�������*�ĠP���*�Q�2A��������vQp�G���ǿ��5$��t!1�p�G�'ur�y�#6�r�b���¿Kʀ���a��݆h����Bq���5����>�M�6��z�����w�z�އ�*4V�R�,[�W��a:�������:Ϧ�BroV"7���}��~�L�?�%�gK��žo�<��v|��n��#[5}���X���O����lr�↻�)oT>��ݗB"7q�g��w�	�~���_-���<�|#��-H &�)4䲽(B\Z�.w_3�҃3�&s��s(���l�͚�1U��(vܜ�Q3T��NB���(�^�������q�JWYe`g�HYo��-{��j���{{���2t��ɚV(~U.�D�)0�?S�Q����|�i��e.Fc���q��gVO�B���C�_�?��-�Ϯ�8�7�� �9��%:��1|��6.콒	|�zVﶬ��\�^�n-���=/7'��>��j-\� �H��p��2VG�?�b��~�/��ސ�^�̭p�?������'��Ji�c�x�_8mfDr�T>&����a�d�M�<�B�S�Ո�Գ*��M#�������_�<:�6?^_/�\=�r!�v�>�.��W���u{5Ɛ^�b}[��Hf�ݾ�*�lLe��"\'*�iK�}�< ���2�BU|k.�0\�g@&�gԻYS�0�����3��ό8�9��|->/`��85����	���т��"*�UՑ�Ew��\+ o��L��)�4�NhҼ7�T&n�k��-�F	��l*�1@�����QE�����WMdѨz#�j�m'�h�N��x/�H���]�p+`��k��s����}J<5�YE�*�2(��ڭkN��O�[P�c��aO+�%�wh��5��#>�D6_�y�ڻ�[��St�����jQ�-����������47�%\����uo<F[�*�{ ���b�TkZ�?�����}g,���Ճ/Q���%��������jԺ�#���k�oh#K�N�~�hz^< �:.�4�,����Z�G�c�A䠬JA�@��MV���z���g�����7��ZirJ_��T��p��M4u;�U-_s-U�*EJ����
��±�6���=3Ȋ�ʿ�4ⱂ�����K:M%+��7�ݏdD�Ќc���e���e���m
��n�Z�{6K�- uTf3{�U ����==��ƴ�}�u� ����U�p� ચ<�͖H}B�s�'�F��C��+�+js=��Pn���AG�n��f�ƾ[9���� �s�N����9�KF��=�-wB��c�{D����'�\j4�+9`|�����`5.Ԉ������\�Y��9Q&���B�`m�&��%�Kl�q��#v����yUi�fF�"w��-��f��k����J�P�&���	|-�<�j�W0��Y��U(p�En�~�@�����G�XR�x`����>
���X�8�<�Ւ��v��,����5��r���c�|2ʨI]kI�䟨��43�m�9$2���]Ŗ���d��n@*�\+��%���V�u!��0��Z6�r�0_�����+t0�� �zJ�2e�/����2��\��;Ю�p���(MI�tȚcط���Qc�x�r����a%3_b�遡��t������D`�[��!~2����^�T�H�3=�>_=`pT
(�Z���`u7�|�����"�ȶ�+��k���@4Q�޴s~[�6�1�ʕ�G~o��d0�~���u��(յ�ݰ`��D.�f�A\��z֙)ơw��6�+?�X����w��ǯ�Q
��ﺭWlQ���P����q`��u{kd�k1�Woo��1?˹�����9U� O�d�	0M�>�Ъ�ճ´�0�]C-x��ՙ|��E�T�,
�z-��5���|yE�taN�]� ��P���s�<��O�1�+I��O�[���M�bȥ��;�Hif��D��WdI�՟�s~�D*/����6�8�r�( ��Vb-���Fvf�?�� �|��U�w�		�k3��9�
��Ga'��[���=�ԥ�9���-�-s3
�YS��F��RK�a��tCfl��@���F�@�B��P��C��쯔L-bs'� NKd���c�� ��z"'l�~v�)v���鞓{�Q�x��T���6lQX���T<� �L���(��(�q'���~�_-ޏkD�����c"'�����m�0�L�N"D �EK�����	-�D�g㭾q�2�/�_���Lw9�U�*>Ń�� �&���&���b����1yru�5NH�uZ���?���� �MaQ�t�Y�J`wڹ"���,�hB^��%�^��,�c!��Rv��:�l%9Dd���5����ch1MN���X݄��U�$�M��"f�f��Q��]�)�\l칰�c�YЏ3hP;!}n�(�W��(�J���f��Qm���#�?��D>c}��8򣋥U~!ؾb�&�BE7��6,���
��Yb�������W]�`�;�`p�R"���RuaNF=��+��*�8WB�s�)���E0g;�-�����.�Ev�u����P&Z�s}��R~�n�F�N���!�1�YX�1u:�i����9�S�|@�u�q;-Sa	L[Ǎ�f�1�/ w��ZLU�C�`��'�0�م��@_��s��_x�da�W�x�e	$[��1�|8y��KLb�����S�90O@��TyV�k��.��v�� Dx�o7Y�v���/m�K�&W�G4�xGڶ.�OQ/�[�E��Ro��b��Vs�ݻۄ��;#M�ثm*����-{�R����0<�c~)�)}��a`��AÀ�+Q�$h(��(��h]�r\�*'�5@6� a@#~_>P��~�O1�5ťb������|eWy3�'I���c
�,��Sn��zf��[AF���,�ɽ��i��eM�E=�rgP�g`���l��X�1�`�cK�S�ӪF��(����R=�%={�, P�Ⱨ]�O6��hے�~�����-&�Cш�����w�ł�ȞF�io�̪���g��1QXp����_�(Qͩ�������ir���D|��U�0(�q�h MM���߄�{6M
����2X��"F����f	3ߦ��xk%���?ʔ�,�#Kh�u���s:1����!3��xHgH��{��+��nk��ܬ�?Q�:��R5IǢ/����5/6G�Dr)J�~��l�h�U��E6Pѵ�$���Y�d���A_Z��+oO��|Yc	nߘ�ߨ~bz���r@���D�:ͷ�!*�Dx"~SӸoVI�;�H���|��X�c{�}��0]b~6�EC������{e~�?q?v����1ă��������3A�]Y����;��?�?$<�.�;�a(V���n�����ri��5t�Fp �HS��4����.�$49����:D�	%t�ψX��6����N��?"&� -�-�#k�U�u���a�~xu�Z 4�F@���ƽ��� \�G	K:�ܽU�=�H�Lqn1�s�<�sL����v�3 {��_y���o_AH}am������A) ��m��s!\&���ȉE����X8��/��L��&�j2B삨t�1�\�k��)@u��B\<2�eP�K �.��D&ғ�53� ��һ3t1�.��z��:v@�b�>���D	N�Nr@	3a17�/��Uꥲ��b���z��.	�|:�Y��u����">;��'��������:��1���n�CJ@����W5�ձ�!V�D��-��hyJ�p�:�b�:3�C���Yj\��7�oK-k��v�M����'ns���mw�ֻ��	R�t�ktՊ�>������l�󪙠��i4F�m�?�����F_i�+@)�m`�{o�	$�{�DG��C�K�h.��^~S!v���hDh}��FL��d+�M� a|���6?�ۦ�T�*@{�(��z��DL���Cʱ��f��/�B$8�ՌCK.���5'��#뎈i�o�d7gz��ł�|!���j����6����a�~ 
�!���3f&�P|�V��"�JY���h8��w��I��V����z4>*Q��O��7V��]�p��N�3wJl�!� L�[�@�����k�@�*`\�� %Z���p5������V��H���͂�N7x
�8.`�E}�/�J,n�_��&�y,7���,�m��i/@�)��Θ�g���?�S�\�n)a�U��ښt2��`�|6�*Q&���i��Tq�AM��%�z���
��f���6t��Ȟ/ta�e�����T|U%� xm��c��!�ǿ;c3�X�ꁺ�'1�(>(7RD����]	�n#`�7bn�*�	��9��ש��T�B�Q�w^f�R�F����/��IeB�]\ח\P9���F�è��:B��$U��bP3�5v��O�.4~��J�CW�����E4ȱ�B�f����K3�sWcm�§�>���)���5�LU��"�
��Y�V��XZJS�-�[�>�L*�̆����i����Ikͫ۔`(���R��kzK\<�e�m�=�hf�D��l����X����B�~nB�D	g�uJF�+(_^�N��*����'�I����g�ї0�	�l��Q|Xϼ0��!I��ֈi������+Q�Ǯd���O+�&xX��hX��F9�G�tfg;����U�j�����;r,��v�:J',�g���}�����pl�7%�_��`Z�����_�4�9x�f1��H/�M��b(N��Lz?��>I%6,�J�W��W�Q&y񣂎��K�ҥ���V��TjD~�tH<-��?�V���Rm�f�F����V̭��fn$enu�wֳ��(��*1 (ses�vy��N9Ԡ�-z��{����I��8��,;�X�{m�C8u�5���~O9韂t�\�5ێ��X��߄���a._�O�&G��1������,2͚q]CZ�)���_��C?���C�����u��j���3z
�2�_E@���著��2�w_��2�@�[��^y�	�k��<Y9*��h
��Ż��P�/����]�Ε�=�~X��%��W�'w���f�
�~��ZSU��~;����Hh�DdB��UM�6��1W��|�ƋJmA��Έ���z�����7*5k@�˽gR��U�oa������9D�D�\�
N��2Ј�Kk�4��%X ?�Q�����X�}�qf�9�y�e@B$�w�r0Ǫ�6'6 3a�	o�U��Y���;�^� ^�-�ۊ`�?r�=��탖蛌e1޶I�o�"�HZ��_�%P,��<�GR�+�Q3 ��-�n�nK]4f)��$�U#Wx�7��> �Rd�`���|R�R�����ES腸��̊��%!���s&��,��=�Ҳx��)�9��_�Po~�D�}�K�@�p�t.+�2��n����:N��miM }u{�C��� �$���q:���\?n�8��3܌��gZ�Z���2����z����R�7�PP� �3�ig�-��u�I�"�A#�;M�gѻT&|y��/:C���A�SP�oq�z�i�<d��D��0�a�]N��D)�����ُ�B�ƪ/��*�,�57 ���SUNx=�>[ӠT�1���P�-o�΋J�K�����4����,�n�#����0���q�9g�)�_���!<5��5(�,B���n ��jm�kA�{�Hz�����Ac�ȃ�:�&������)Ǽ7�k.?_��t�\̓���ܚ˞�tR3Q�������Ju/�Ԣ7s��>�\ ��z 炆+89��[���6��A���u#����5��k:����D�P���6 a�If��5؝�!�	�a�:;�:���G�* ���)�LN�'yF�h(B��g�2hv�G�U#��e{��j34���vpl����\N ?f���	}�M�@- k 
��c,�p�]���L�^CQ�ܻFq�{��Γ,��hN-�o}�>�m9$6�����I�Ҟ��m��2��.�7�zW�u�H�c�z�������!]�8��;:ip�Pڎ��}^��l�rx�����Ip�#g�~��ո�HQt�*3����&���H(�Y_���^[��HRa��E�rB1% 3S?��%�0�?������Щ؈�����>���-2jO~�шC5y �l}�B �{&�����,e�M9<����"�� �kO���ˋ�]ȸ�3`��R�:)R�|�SV9�o�/�VY@���*0����p�4�ʳ�3ۻcq� &�[��o�%�,���k�%�87"����@�t��'��a�_�G��s7�I�#v ��\r4�����@+�P����v���!kۡ�#�(��T)�{�Աi�rg`�b������Ae`���ݬ��$T7��KϾe�u�OkV���.#����2�B~��Z?�2ָ���F���&f�6�1$��vF���`�$C�/;�Hp�w��, ���ҏ�k����'���웃z�&��2��|����8�/Z�db$���<�U��ת�-�wH� =A��v�V�\�ūA��޵͞�8󕭲=�Wo�}xk#�A��o�֒�!:r�Rtk�^�u��Bj[+�I������0D�Xp#������y|��(J��?,�>�Dh��c��c'��%BPG�6���@��bO��Wg�e���W6pl����?����������>�ÿ��!Y+xEE��8�5��:;�`���k�R��P5��}e]�~"҉h���Enm��H�ڻ�@j'�CI:��`��>���N['�?!Z@N̝�Gyj ���ɔd�\�@+T+�2�#3��$ݘ.m��٬�A��p��i�!����^��]L����ca�a�iZ�4簱����QB��G����I�5�z%�b�@��. )���)��F��<s�!5)��HJڲD��|�0�*R�/�m)Q��5�L5�u7��1'lV1�J!~�p?��7#��&7zYQ�olF���6��)�ax!O1P���	�/ ���_@,H�H�L��TZ ���y���rvE1�.�;�d[L�B+ˢ��&X�5·v�n>���7�d	V�S���IjWP��V�q�y���M>��-�zտO���b�
��*�:��dw����ʠD+��\a�k�Z�@ڢ�_+	�!` "�:�'zHE4w���L7≇E(Z��Žr�3SGam�g>���FY���K#m���va
�(%{QG��Y���n�	���D3?բ�2۫�HG��-أN�x�%↽oO��Z���5M���[�6T޹���b4���זDrG�ؗ]�M���m�L�Qd?��Nt�rh��_���c<3�c�`�!�*� �iw2��Or��rd�$9�ڰ�Iu�R�<�#%��U�����6�Co/�(�%�O�xn�m(=BJ7�i�6>�m�N��؂��%7�Z~�Lr?i�x��p˙Nh��Ms��g*�:eE)(��jxĽ����.�͇M��1c@&Y쏔�o�u��33�ba�����z�+o�刺j�?e�ڪ��"g��Ax�e�U� Gz��iC�o@6�xč�/��>�����w� ���^��^�S�s���M�0�L,Հn���0��{IX8�����`��i��_x����ERL�3�V��P[�j�T���c�~��H&ct��5
��̭
�@����S�=�{���`��63
��$��]K�@$��&?����Q;�k�s�z�YH�'��*s�HNL�)������_0FG��x���&��Y|4�ݛ��(�c�Wa�h�~��y�eA�F�"��V8�щA�~���R��S؊�b�v�W�e��[<�r�g���T(��Q�~h&u�q�:Y�a��A�	�%���gvݬ�����Ч+�`J)E��,N[�R�f���_�A��^���t|�
�H�;�h?���+�#�̬@�ԛ"��B(�T�����uN���N���yRn|�ل��5�Ze��]����QsіmO$+
dd��}�?W�Ȇ������V�ˌT��K���x"R��4��c���:v����3�Y��l�2 i�o{��̼
�st�c��\����ǖ��}C>�K���i�+�)�\��*��}� �āf)W�#{M�"j����h�}J�]7�/j��Oܘ���L�N�=��P�0B�%0�uNP�*�C{�Ɗ�>�0Z+P��������c�F�!v��d�.P�6�\�x(��+T'lTEڞG����I���� �L����2�^SV�D�%�� ��~G�����z\��0zK���3r��x�DH%�D1��~�AAM'S?s�i��ٸ��_��-ܳ�L`b���p����'=UA[@�,�s�x���u���p��/��C���s�)�K,=��7'����,�e"��*���v�p(�V[� ����ȼ�vU��:~\���=��I&"-h��o;�k��YS�5��u����%g�^�$���Z����7�A�fK�1����O	��6_�o����Z����]M;8:�߲��F�$#���G�y�>qҖ���;���{�62::jd������(ze��J?��A�G�R�~EAR:V��m����/j��s�����%۽��_20n�z��H�5�%h���������H�M[����W@��5�aH�����oz'��P#D�o�|�@nB�כjNR�ko��	 ^pK8+)ě�����&EF�mwEk(�91�7��%�M������ߗ�k��&��s����mr_�
G�#K���%��x�)����𣼦6�n0z�B�@(����B+�ꙟVx|vD��ۺs����:���y���H�W��	��M1�����A,÷X�-�ԳT`Ya����8ǫߣt�i�d>	~AaZ��lF�f�E�	`t�z��$>��$\S@)��62�����
µ{<�@I�=�D�g9��=�y�[I��\+縬P����R����a���i�g���H!�4����Pt��bC��L��1D�tY�'�X��;��j?��9�r���v��8�MCM׷�Q(\Z�I�<�h<�F�[B]V�;u�E�C���0��vÞ�w*��	��K��猢�(��Y�g:��K��AI*��I�.�ЇW��>��Y���H�`_�/�|$C$�	��D����u��HY�K0�*�o����oYgy�����$���Z9�غs��� �������F��GGN���~ .��ɏ�����Bbad��
g*�>�<�{���ƛw��c}��i�Ӵ�,����K>_�C|0�^�	�3t�	B�77�ᓪjC��r	����$�j"z	�c�P-,"��G���*�?�t/E��)�z8oS����qb4��rs��ҏ�&�m���5a�޾������˄��:v'q�n�8v�HՇ�}�Q����6�%�l�z�B��^�4���J5��;�o�/�J���X����&�*�F�%�˥E�_]_S8�S��L�;7�:�����.+w�9-��Z�5~3��P)� 7N�� 	��m`6�޸�(뛁X�!683} 0&x,|�B�6��_=d�Mh�5P�ח�gDy�"��L��T��q%��/X!9�K��;eJW�##d�b�vj+�
��H:?Է�E��mnT�_w'S��X��`��^��L*�O�=gA�
b�(�- �=6승���zP󴇗H��9�`�!G},�5�mޮxɃ�/jr� � y�1 W��M�� B:Y��?$�{��Q�v��j0�f*�t]-#E�#���PI޽��<z��N��V.��i�EQ!c�3nS�^$j.i���R�w�C������Vj_��x:�M$ ���r��%�|Z��6H����#җ
����Kt%��|7�[��o��6ޣj��;K�vx���'�(f/���$S���8���� ��I����V⪪�!�^����팺�z<���Y��L���18�r��1����B\7��/EД�~�SI%K����v�CJ��_IHS�[��@r������1����Aks�����KFƆ॑4C�iN�/���C���h�M=������'QB���<��A�ON��Y?��7� �	���uy���E�H��Op�ME��a���?�4HauY�O�M��|"�!Os�a��{و������[z^�f����y��D�=t�<��=�!S:�po(���ﲢ/V�at��r���D����Hٝ�?�Ǆ�	�(��7>�14�o��5����\��X���L��#�Ұ��C����$�T�1JC��I@*<�5ėg˗�#s�f���}l�#��5���	B���W(Y���o��f���+~7K�C�Ě�V�-y�m�H����OKx���oPc�hSh(�����7�?�����������umz��h0�b3C��yj�/A:�X�u�s���t
�6Y�����<	���f�;�$�?�|{�E��O�I��u��n|Yr���&��$�^(Y�h���|2�e/k�����D0"y7��rf�����]�Yo!?+O2���r�*D����J��9�;텅"�~ǅ��6�y�~D�%(uj�T�8��Ia����7�{��q@:�4�5Sܨ+kr#��]\r�0[2�}��*�ag�0�.B��{=�����C���$$T����'�]$Ǌ�~��5ڐ��\}�ܭ��6F>[�#f��Gĭ�~:����bN�
�q�-nQ�Bم����x�,eS*�;@A��&��Z������nH �>.tov���&�<���u}��[A��H�5��#�yI���c5��:�o�R}uW��kM�e���s����+0�TE�2P�Sl=��,z�Z>b%O�us�������I�H���ޑ�˻�Cl�������ޖVзDh��b�StY��� W��;57r��vj��-a��ɷx����'0[4o��j=�0&Sk�&��O�O�R`֜]�o;�5�߯�Be���v�^o�Օ�$q
!�x�N��-'a��fFP&�%q��p�H\˟��k��C�vRɹ~S�4D3Q+{?��⑅g��Y��Y��^����?󩱵�V��X��Dy���;`7+V���3'��g�A��H�R�����Y_�n��
�-L���ה��i4!aZW]yk�&R�⊸�8�ûD�)S^�
�W�LQV/��I@�|�I� j��C���#��&��x���h��J#���B��L���H?mf��4��gx��~�go�s?���D��7-n~>��B<͹��i9
����Z�cq�z���g!cAn�G� >1��Amǘ�:ۉ/��W��c���0b �ƪ#N>2��gv��i�� ���?��ُ��T�ɡQ� �.FP� ��+x�R�>ZU^�M5�+>�c�(x�-c�O��A�73X��IN�3Y�xOC��6��P�	 &�z �yT�,�*1)�à����Z��ܙ!e8��m�&��'��8��-�Z��H�������If/xv�c9�����wd'ב��ß�zt���k�'N|;�iT�tD���wfA��	�; ߭��R.(�)0��g}�T�)�����VN�V�ᏸ˽D:�ïRdlB���l(�����=	���a~��f�ي�#�P�=�g�P�e��X���������1����S����5�wKJf�]fl���C�`:�����Ԧz+���鏆��Ti�4��s[�W"�ݎ� ����ن#r��PHX���ԗ��:e��?�~���jէ�
�;6��s<\�J �Ӥr$.}[�q��c}�g��uHM~�54���Dl�(x��Ħ/�o�a`�.:T�FE�$i�,�#��j�Ϸ�~=� ��ꞥQd;��9`���U�W~1����v������ȭ�`c��`��i����O��YoyC��/��EzN�`��)�J���>�	.dZ�˂JU�������u�q�.F]�L=Ƹ�b�P0�a$��>�>�B�� f�`QuR4hչI�p�&Yy�[�r��QS���;C�(����x=�ġ�W�Bәt���n��E�W'�.����4N���@��S'f���ǒ�k����4Z2�)^p����OC��ȶ5d�.EX7�'�-�_��Ҁ(���UQS���Q9��)9����@�ڏ��#"8���	���n��L���Y�t�Z�j�!���JJQ2�����X]�4�rh��:c���LD�rw>�_�����H4z{�r>	N3�k¡����q�/L/��8��F�[�Ͻ���Ž�7e��-�N��z`@�TQOVQ�`�R�	����x�ج9���Q�<�߃ � �sE}@-�N�و���p�#��P$ͅ����Li�ؽ8\��+V�Wm���]pʤ	p�{|c�B������k|����<�ۈE�H��I�L�G+���ɐB����?�~�X����}3 �ݜI7�w�N_�R���krpU�������
�u��Uk�Y�U��P}ڂb����js8�����k�L!�P�l�cs��]_�8a�X��_:��[�ه�i.���bd@E.x	���K�,����[eh�7��ɯ\S�?�X���c��W�R�sn9�_��x�;�<��-\�2�۠8�^�b̋y�/�>�)//kn��������j�1��1�K�[�R�4-�H������i��r��g�9f��c�M�Z�b�1b+Cf���8T3��n3u��k�V��R0~�/Ѳ�37�����.cP��h}��[�ܿ˼��sai����O��<>�*pcP�6uҳ�:ؐ)ρ<z��Ks!���M�a"�������r͡Z�hHY�1�ND�T%��Ҭ�t�<N�Ȥ_K��Uxk2���89��A���̠c�p���!|-�>�$a��;�Ys[�^�Rc���X�PMSu��~ J�	��N\�G��~�B%��\2�������$8F�8wߚ%*��������d7}ŝ��Ē�2�っ��]����f���\��Ax���Xg��W�3�������d������۱��O��h�E!fB�\�x?m�.�mLT�Z@Z��Uhk�>�D�V(��.�l�^kB������!g�Q'�
n\�� O#�(.]%�%�#9��l��q�j�G�w����-^ߩ��] ���u���%�|�2I
�o�m�vk��n2ó�x�v��~��r�,r��1�R�44��=(��#WvK	Ar�=7����6,x�n1�IW6:a2=+4��0�p��c�Ԁ~9;%\��ͰQ������$�Dg��Y�7pc�w��Z��^�Os�����!�_��4/u��b�+?Q[Sq���X9��R�:�t2sg~��H�����_Gh�D
0t"oy��V� 'u����΁U��hN�V�o��iȤ��8����ϡCCѧ3`����T�O�$N|�]���t?�:�HA߃�TP8������~�b�S�� Zë�g$�:��k���6�6<��SU�K�t�Ťv�⾋�L���u_�Jb��e��u~+�Ua��9r�Svq����K��s��Z�[i��.D{%�e+Y��Z��P��ӧ�*$��?�(^�:�AiC1p��d[{G[�=2�O���bZ�cy�
R)ڬ_�o��` ��/6/9B�WlUx�u�Hk��n�n��x���t4� ��7��4�1��ڤ��B-/%=ܡ������:J��s>=�G]d��+��{�k�%�R��D4EGIL$�|��=1�����<[�s0�g1�n� ��BԜ쯭dh���'��k��Vp�e��$غ��8�]H�t�*'�s�Wg��OyLn�?u��x!�z�2K�-Ҳ��_��)�І�Q����I�M�E/*�g���|�O��B�RZ�B[��d<��\Z�E��P��ݴ�=��M���N��n�3�H��B �d�'��EH�k�������+ ��o���)g�\o�ժ��.n|RG=^4�+���0D9�`����3���a�i_��Ge�:�q��ne�6a���6�c�򖎳�Dg刉J.^��k}x�u�Q>�Q'��_G����AZ����́��HL���i�B�ͣ��H�K��b��9tg���e��\mu�C����0 ��o���)/W��j�q=��/.;˼T�����/u�'�Qenyk�u����>�c���F���N�y�����\�5�pm����+S�1�]IHg�k�{��ZA�U"�wkP+:�z���.�@�	o7���Eh�C�;a��A_D�T�:s�q�퉅'��3{�*��+�TU����܋�O�Ǜ5��7���\M����3�������
SIU%�	�p�a ��tar���Sj�/�e#��5�(fq��
,�)}�rО�� adm��;�|A��X	)�$f.���,���6�a �Z>��+u�����Mgv�����ޜ���7�6S��1�� ��4�]A&�,������!�8�TS�>�g"����fu�#�伝�[���`w�fC��SU�����q�S��L��^�!���g���c�WH���A"�FK�����,*���;��$�-h)C-�P�-[t�L��bח|ߜHՖa����K$`H��kqڪ,�/�ţ-�o�.��la!v��\`{��a9N�i<���A,�,r
a_x�mr�N��yu�p'�XS���`^���5�,:��+��2~�	oep�d��l��L�+�L4`s���&�^4�|�p��б�O��~��z�+T�,��ncH{H���ܖTPBju���{��z�p���j�l�s��~��x	�Ѧ�&s���#i���)~Q�a���5y�`)�D˄/D��50��%�h*��ہK���S�$�!�O{�n�p2���Dfyb<G�3����q]y�)��Շ��u�����A���(�99%�FT�mx[7�4�U�a�ʸ5�fֶ;Ν�[\�i\���dJ��n؇Nw$�Fؐ�՚l%�cc��;r��s��PS�;��o�m���C��)PGj#=���<ÀZE�m@����?�*s���y��<h(tWc��3 i����mM�h̵G��@��{%I�0�+�	r�J�I4���� F8X*%!^z8c�tQ\��M�F�m�Et�	d|J=�ayf,"�|d�A�q�Ӑ]R5����t�!J��}i���܈׈�&H��o�#��6b��\(�gȌ�2��gH��_&�!�k���D'�`ԟ문� �b�08�m=e����@I�o�V�	S�]r�
\�|�=/���TL�C���HQ�LM��,�ׁCe���W<�����tT�B?���'����b������p��`�L��_�l�D2C�"�2z��^Ơ���S5!T���FbĨ�G��7�i�Y����A�h1o�/N�9!U1.�׉Y♉i����T�M���t0Hz����j@'�Ոi��Ȃ��fK�1�h���\�Ɯ�s'Cw�."�{î��|pF���ģ*���VQQ��b�a�D ����=��D·�N���QI�����u� �v}
8Ɓ���p#�|kq�D��O�Q<t�
X��h��{i4ŀ�0>�����,(����#���ӢP�Mb_��/��&�+�3�1�xb�'�؝1L��p�獉qyg�(r}0A����?��N��5�E�x3�>FM�?��0�$�c��$>�/��%�	$:{���\.}$����3��V؂�K·����'[���w�j���z�0��w�0��i�h�pg�h��m)@��T��X���~��4=N�t�ڐ�Q��tr��Dꎘh�ɐ�,�h�������<!�}I2�"��?����7���3 iĚ;]��OW���w�|���<m�m�e|<_�XY�@7s����5הٙ�!�gG�����.�ޥpg��Y��E�C.r;;ͅr���n&MG/.+�����6ሩZ�"�nơ�UXVt4�aJ��w��f��T����:�Q�1�]�2]��v�M�gn��{�̥�4|��RV'W�?�wnwzM�=�p��<���l�vui4�c���n������tY�O�Gi#l�	ӄ\��I^_�t9��>:�4	�i1��,��U��Ȅ�(N�s_��_D��U_�5�}�����Q�R�w�.	�xޥ��"XAj7t�0l��!y�A�o�'.Z[Z�eϗp�'湗�2�x3˼H��z�%����~��r#���<�?K>�s
g�1�1�x�Y@�����]H�F����!9���H���(��A^*�� �!�� ˝~��5 ���%3���޹i���y/a>����}�|��� 2a�M�̪JV���%���Y_V��^`��J	���	(�²bt�>~��Z|O��@�Im}��?M��E�2��#���3y�����r>��a͵ �bv�<R7�+d��ج!1Y��	ޅ==��C��܋P�2�(1�Nڞ�Hpti��k���$�#(�5L�+���U�}D��6���S:B9�����\��|�:��a�B��j%��c%���S���D;-;Kbj���������$��H�=����eC�n���ێUٌ�?��ws'��T�Yb-��2�����g!��!�*��m����G�Ƶ}܃�����#�3OP͌�d@R�l��Z.��� 8�L.R�!2�5��Q��ؾ��vNìC5Y�=�
��r��iӼ�ݧ2�t�-]��\lx�xN��P�)qCq�86��crx|_���u�ݬe ��^f�����?��?w�����L�B%��� 	�37߂�8*��LqR˧vnHa+�+mj����o��np\��nꮠ_���;��H�F�L�y�g�%��D�5�D��e�X�cҐ�U��
��ӺV~�Q-�ģ�(��~?���:�|P���j?�?kx����H�9B��'����+!C-q��8���acf�|�z�i2�s2�X���jWe�Y�
�Lן����) ���}�Տ�6�P|�	�����yHgd�D�7�:��{E�WLX�a䁳I�!���`إQ�VK3ɱG)�LO��]%�����yْ�`�ϩ6�>�<$����rM)�1hR�]秒-��;M��&����͙zl��.�=3���`��7�'�*��TgB�#��+�4h�9�����B��H��#|��V�5ӹFO~�?ϴ�7[�����^;�u
�[g� ����eU��+���w�3^ ��0Id�U±�(�n�U��ߖ���M*��d)�p��o}W��wXk'c!a�1Tk'��2�"�X�����<`����P�eF����g�f�2�k0@���O!�[�e��O(�����x��x��Ͷ$�_n�/���P��Pf��!�*&���ߨ�L��:����mME;�&�Bs����LJ>֣��1�M����/�9;Ģ�z�����fO��ݍe�3dE�J����$��8�k; 2'�Γ��������pph�c�X&sE�bL�,HqL�š�x=��"�i�.r?�A#c?/�I��h"���^N�U[e	]��A+$�8��(�(N�q^����E}��D��rZ��$�J.��z2uNfƿH=�x�lk��B�q2L�y"�I�!J�� @��*T!��A�}.p��=KU�o���$Cb��B���j6T͞��+d�r^�eqM����X]���Q�g8D�����q��.�=X��W�ɖ� j���wX얈��.-}�����H��^���['�~6w�JI��1� <H]O��8y��@�W"�ʢq�j�D�褐�>���g����#��sϿ B����5-�a��%���Q
 ž�Ѵ�<}c�? �d�9��r��p�qV˥�0�*]s���Yn������xv2��}���On8����7I��"�.p��F=C�,"d��.����D������s�NX/�H�%�|PD���<u��p�v�k�� ��P�<����P�d��^�G_�Qw�G=��&�1M�O�d��5�т��]f�h�0�$��7
8Fű�;M	�~�G�e��W���|����h'���l���-ƴc�G�e^`���� �A�)��M���ޔ�s<�Gp�i� �r��
؂���y�QCpծ�]Ī3v�]|7������S��hّz����|����3o�E��VAXSŚ��s����;�"�芃�\�\c�!�!e<�	��G�9$���A��e�V�Ԃ�������-aDܜ�y2�f0c�A��d6�T���ѕS����D]�	����|��>mu��3Վ�7hW�1w ������f�#�/�O�||L$��wbnC��U�H��������a�	<d8����'��h�&0��y��c����LK�Q�6���8�� @;P:r��ʼ�	i-���ͧ���[��HL5K����0��aU`������`�M���[l�>�,;�/�8G]�;=2�������e̚W-_o�Ğ�D�Vk��>}�6�5�>��a�tb��\��r��>i��Љ�0��r��@ <�W��U���/��?����#M�U5��J�{pE-�+��v������Ĝ��iqRV	:������J\fo1I�9�e����{�ܹ�Z���~�ܔ�D������yon(/vpɤ�*Z�����<�Պ�;H�Q��:��ߘ�^�tDpn�hَF]���Z�,��(/�$�M&�P�A �@��`��} kB�_g�ʁ��T�N�Ps��:��©����~�6+"����t���b���R|ю���[T�����K���O�b�K~����ݠ|��2��C����l���s5B�w�/5�s�����8�]l�����`uk����?�S �ğRIIg䟷�,m�;����MT��B��m:�J�g��BǠNh���r��ȰQ��(b t��,y�D?��0k:�<��=7!���7b�K�	�$my[� �`VO.��E9i�[� �\ںp��)ĨD�W*I�
�C]�������]yX����׼i��Mz��6ja�$D��8:��x�Gy\�����y"P���L��24�N��'g���(���~߱��Mp����Thc�J��O@q��B�I"�*����9��o�

>���dj9��ɭ7T}��b#a��@In�D$���CBB���9����L� 2���r�%��bf�Oם�0fï����4�f$7�e
�����ե��5ɂ��xK�$W<�?kѾQN|�irH(ɶ����׈B�-���|>%�@$�O��S������Λ������Rq���v�*�ii˗��~��2.�s]?m����'�Rڨ-�/�Z@��.�UJ���c:V������/���5lT��/zR��4����De��2�u�������+��Y7'���)���!:9������sᨈ�$�]^pm��]+���������ˡ�6� �ΜWR{-�F������@���JW���s��^�|�T�h��ܴ��r�)�"��� �W�s�H �,D	,a�)Z�֥V��Ycm�{�C01��� T�xy#$ԭ��r�C��!ִ5��r�E���b,p}��=P(��iX���K�o��T0���7(��f!\�\����w
�w��Z(�������͸�3ߓ;�֍�o���b��}�����=Ef�>�V9F>u{9��A!A�p��0B�Q0q���:[�z���h��$.X�aY��:�
T���>�'q
d�z��d�lV�J�~$dq2��f�*7����2��ꬆ@��]^��־:�5�x#��EI)q4ކ�_f*��5[nb��1}t;�s�JC�O=Y5�/xf�k��Q�=R�V�6��Z�F����-W�0x��s.A�?�}q�5T����3}u���m�XI�b
���nH���W8jb�������݆,��7�ޕ	�e����1������Lg�o#Y=��"5��e1��Xb��O�֕���qv���Ζ,x���Y��#�&J�2��L�[�n��.�3]�����̂!���+�Ct�ʒ0�ɼ�* �5,J4XȠ)�<�m7~��"4E*gj�u�,h,n��aњ��cV��x�&<�l�t���^X��v�=DLi�R-z�%{��M�K4�٘�n�S����/��Δ��U��Хf���'����qJ��/��΀(������وF�' a�t�?��kw��K�93:.��U��dsd06^�ˊ�߅�G�#d�m�Y�%�EE,H��+t�}ŦaU��hkd"�0RDZ2��C��O=��E���:0,�#o,�<7X9��L`�<U��{	��e��c~�.k!����12���ɧ4�`������{ϟ�a~M����8�O�~B���n٠]p��Ҽ�����&x;��q�����
�|s��j� i���S��r�I�\� �O��7Y�}�Ɣ�Ė��s [��/C�_wd�8G �2��Ŧ.�֢�@i�|a�Ӈ�&�����\qvr��9۔T��Ӵ�
g���)oc��^iY�u�K=�y�Q���|���лݷ�����!��k�@<�?�2��p)�����%�TM�]����A��l.�n���o��$�+	.j@x
��g1C�"��c����@��ts����3�i��e��G��ag��q�}�q\Ϩdv��V�\��4���6O�e��;��-c�)E7�h^c�0=���/��T�h�L	�³I�ޅJ
h�C ��m�'���1_fz����/�+�#:�f�K+"���-ٲQ�l`T>q��1�|�}�]M��w��oc�z�A�������<;�g m<$���Q �Ҽ�9np�8�M�y�Ii����D�&�q-"HK"�}�5~�����r���	<B�+�.�z��>p�-���2Ut��2�z�ln��U�	 BŨQo�(��{-��������ČNe��tx�����O�~"L�g:�a�5���A�A/�ä�����P��L���.2�Ɇ�B�X�¥p�^Cd���X������ą�G�H�B�;�]�cC�ң����m�=���e��Rý����ה����D���Px�׉��=*�)!Q�⌒.��WVf�l���@4�t���{z�/�9�&��$�h�7g-��!@��Q�&���~�>���I�zQ�w�$4�N�3*ro��!{(����KP��@�� ��ߔ;������lJU��ϪĲ)����qr��́(T�5���U��G;��&@:R��Cg8���ۺ���H�����5��/]x�ߣl-��b+�l���p���	�	O&�@��^N��@�I�D�)�������(�����}��숒��_'�/���M�f�W>�Y�q�k�jl�����r5	U�8�.�� ���6�[J��;[�$#�oP�W*�rdar����ԥ�q�D,j������ߗָ�#�$^ +���ڪ�����
;i�0���tr&'�	R�
U���Wg���3�wj{-2E��&Ph�����o_��Z��1����E��̯ʼ�vw�*���z̽�籨}3����'�ӔI	s,��,‎�����h�Tvr~:u�_K��Z3���a�	:���������F5�h�s��n>*�#�!C��5ޏ�F��7mS�Q�_T[�Ɋz��zP�S�'ò����"�nu�����Oc��~�b,�)d	�Id %gX�<JG�n�_2�fB4�\ չ�jn���j���l����Yr �N$�ڄbƯ�t��W���p3�� ��<��z`H�N!/>�ЇQS0/�|L���>i�����?h9c���Nz�KE�c�k�:���l�"�d@T�������S�}߬{"�Uy:�'ƾ!� X��$���"�n��T�W��H���c��+�ڜ���Y�[s�
�u�z�w:�<*�R���`��U���zq���&�{*�����!�?�H��&����	��Ik���y��ع�M��ZE��i��{�ׄL�� c�r��vO��w,���bd3�J"v$RXT��%j�Bjkd|R<��|c��p���g������Uoa�O#A����瑌�ԇj�J����[$F3O[��h ���>X�^%H@���YUE(d�'q��W"�F�A
���%�#I���k8C�*O���gw��}�s��`��P���u�e���Mq�Q���.͙�/d��+��K;Q6}<����K�ZՁ{U=U`p��ߋ$ldӁ����e$ۅ:rl*�X�LB��3�>�������q��&cT�"@zDg�t
�'R�:�2B�fE�X�{�Կ{�i�ȡG����"[��i�t����c�w����+9���˴��\��hC*k����li��5��!�|�R���*�f=')�=Q~���箅���6B�C�A�����u�X^C�����ioK ��J��En��[��_�cjܦ��Ӡ�)�0!�N�睋�����[W���O�����y���3r�9��X��"���ՠ]C�U�1��U9�@^�-�P!6�u7��_���{��L�޼�T�b���i���O�RzS�)��n0|I�/4�����Q�Vh��J�B��ԥ� ~/�@�4��@��nNX���vcOtU݆�X$C��~�_9�V"�죡^͋���x�)ETV �cA��Bʸ��R�<x�������� ���(�K�֤�]��WCX�B�url�� ��bTJ;'�MB*�:?I-�S|�H��0�m�;���h���`p��;����倂�Y!tDP�b�S�X��v�5�x������<ܰDh3���*��A��'� )�c�'����"* گ7[�Z����y��;~�*;iu:�;hrZ�{{�z�W�^��'��wx|�>g���|Ӑ�'�F;�3	�I��^�T�U@�s���}�&[AYá[�t�޻ËAF��)���Ί���(9��P$��i�[��ף���T�A��7W��F��3�/�^Qgh>�S���c͞�~0:nQ�-�$5) |���Ge����?tKZ*��<똛����r\2�U6��D~np��D���`>&B����*m��"��w��5�A�U ̓�D���(���������M�n���faR�B73s<[kpV-db)�E��*��[��=�#)Z�m;ۊ�췑e�<�M�ĸ!{+,w�C���������F��6*l�"�#	A�����D����K�Js:�>)t4Y��,'~���s3�%�9��Ê���*BSf"?ߥ���1�]�e	0�e;�0�b�Yp)�o�Q��^F@����s�j�l���(�������k&��OSL�(H������39Wmw�f�;���V�,+�;kq�W<��xֻ	߃s4M��F�v�л0.�x�=����ʩ�L�b*̎�<��D+k���v!0כ盈ĥ$��,��ޔ���uf�!�G�J��o}!�n��j����V$'�[�ޘ!jL����@�ϋ9ӫ��6��n��?5�3��6����K�ig�W|BO�iE�Sy�``�vBQN��lSn�fI�.p�s�x7��ug�a��XM������ѡ��>��D���z�5D�,�@+
��N*��`�sɏ�wU����RLu�0�Ex�Q�E|o�,���_I��nK�>`�;bze�}��
�/:��r'�E���пC��-��`�K#����v�X	�wn�[s�'Y�$bΰ�Ž�&��Vh��	4�/Mv>�`)�C�&pU�g���0���Ǆ9kP�Y сZw>L�lzrT~�s�<L*���!�`�Uf����sJj:!���b'(B�@�`E��`��W�T���>9!�ut���i�C�c�`�� \�_�� �V��8�v�\ʳ�j���&��-�$�U1��i�JOu㚟;�b��h�J������0j���DM���hv��,f�k�]n8�X-!�(�ҴW�X[�Ԙ����to��r閨�( �;��C�����e�^�����_iA��Q�~��$�"T/�;��!��N����"A|�+Gp�uϕZ�i��û�ۭ7�X?�r�
�j�H�6>K��6u�:Ɂ��%�x(}���r�f'te�ld>������g���ҁ��l9yA�<�I�9s
�=]K$��iG��M��>�}��E
�S�^]F��=���x;�i64΢G�X�/`��1�+������ڤ�eSմˋة6BH�we�&^x*2,���F���UW��+����yN^�o�= `�s��"=��Q
���{��@����0�����PZ��G%�D���a�D��Ļ�.��a�) V!8΀�X]Bǋ?��qX�M"W�9-%�2�!MS�kN�����>�q�/���C-�6Q͊_��u'-��(���+'���6��ֹ��[��ō�>�X'�8�Ԅ�y���:�T�"i��AP�8���	��~	'	����Sj�'�B��AN?K��u��:���v�$�����Q�a�{�?�^8K���G�$>�p����C@��x����< WӤ�G�ozzxYn�����ϫ~���>.a���l�laU��tZ����@;Ql���&ƖK!o� �7�����gJد*�O���>Dc#s��d��q�	�-��� v#"0bdQctʠ=�.:N�^'����	ɫ&�t*L�d�l�a�b��Q�� ;�/�'\���^,_F"�@DE���9�Q��齟�z3<#�=x�z���Q�Cc滆_-�^�y�J��D��ʗ߯�jz�'�C(�c徝]蓡G��@���� xI��)V	j�!�K����O�_ƘZ�m�r;�OYq��,DI�R��� �e&�{]��;B��z��?������R�mq�ذ��<������T|V���ʒ%y�Q/[��#Pa���!�(֎��:[�
��\M'v�Q�ͬ(R6����ڶ��W����Q*~[$y��/�b����RЈ߉�;��f�F���b�VYBs5��&	�Q�i�o�N.2���W��(���s���P�P$�}9P��g �.��﷘�:�X|�����6�{e���x�BZp�ʥ"f�<��^�;�-r�B���
���
U��5k�O����ִؐ��
���]�P��L�j4$���l���
	�&��������M��r3v�]x_�]�<ĦD�����TsJ:��Fn���'W��f�A���Ye�[Tb�O[@���t�@{�ϡ.�>�W�%XZ8��i��.�׊�%Q5�@_w�����M��1�Y���\��\Y�vl�#�e�l��C����~o�\�a3�JuM�����b�����{��.���Ye!��ClxF��QsQ�h
X�ږ�%��Y-9'$R�t{�&X��s��Aʰ���K$���&@W�L�+�2}M/M���y.Һ�Z./��7�>>E����`=��(��p�q;^ӻ� !y��[�5����|^t���)����N�k넠�!!y����|	$�G��|�,�)��
x���ц<Q��}�>��4Ҧ����N�l���p���
�������6d�wU�T2�˼�$1�<�g"[5��|ź%��'�J��A^��|EOzͺ{k˅���.��&��MNQ�n,����Bo�����|�Z8���c��y��Q��h���r�H{C���{K�W����8�� �[]�gXΏQ����Y�F�_�8��k�6��kQ���jJ��tj��aDJ��e�V}��3�)u�k�����B�\�1��N�2�]Bb�,�r*[�c㚒x�)�S�0�B�`&��	Z\�������´K�ϟtA��_��ic`�_T3�Et�ޞg,�T��$�Y��BC^<ǎ�Z��|ɼQWi5C�
�-���Z����b�4�$ͣ�����\P�j��t5����>}�.�!�$jq�Vw�y>d.�CVP���G1l��ΆM�1єX����)G�W�IU�p�>���j����t� A����������,�z�O����9F�"k�"����u�`�XM�ꄋ�H��e�fh$*:�@8fr°�x���#$ /C��t�τ\�����YS<�L�Qr�%�!A��ul)�
������6k0��[�G�VPJ�`�ؖ�{�/����M9�G]��7��C���pw�x%P)o<~?�n�����BUPVkj��'.y� 
k��� Ŷ�=�z7�HS]0�6�P���1�?/���{��j��ҷ*�D&�QVנ\�w��8[ 3�?^k����ΤOuQ�Q*po�˺��'�EG��(jM�?�7���|%��aL^�2��	��3��T��Mhx��4 ��ٲ���U�iw�!������������	I���#6s��^&a��#��#����8�qf�!;+����:��O�)��3��ɾK6+��o��e��)�DA�G>���^�������8dj�Q��BR1~��5 ��m���Ͻ���χ��y|m!M�j'g�l]@�3���y4Аv6Ɔ�$�Ғ=�(Y~\c�����"~�>ﾠNM���`�1��}]#6��_���0ī��N�N�#�H@�5��eN� =�4�J$�;n�I@۲xp]T�:���������]�0K�i.Ҡ=����8��� W��a�݆����\d�uY����.r��'Q��Y���Er1��f{@k�q�0�c�`��s鑕�f�zr��ؕ�R�V����]0W�N�A�_[��^r��aG��`�E��AT3���꛰�4__���}�  �(nM�A���'(�ؐlD���p�|����ޓ½�����	\���Wy�ۡ���Ծ�����R�E�s;!&��R����G/�E�,��|�ǘl�,����z2���uV��`.�>���:�*��'���⁨�g�^\?�����+�AB��r�9���0i�b�f�N����W�p�(t?8R������~�1�|\̥@�8�M����f��N�p��k���l۪��(�W�![���Z��7��A�b�=sm�4ov���_*.@�b���$�����0��r�Z@"$5��9w�O�J�f?T{��{D�Y��_w�/ZG*	��0��h�4X��M���:T.o�	{X�AS5��qc����}�$�o��f��S!����w'$	O�q"�Q�J�蚍�u]a�g3�T�Ů��ۑ!?8T�(�eK9�<�{-�K4?<�N��Ъu{��z��ݫI'�?h�򚐱P��lU�;|�n�O����M�W%���	C�\[�1c����tp�V�WI/e�+�n B��=���tX1��#��M4�׾vHhm��/�׳�V���ا��#��F��f/E�i�ﴚ�]���,AϬ���y�4y��/� �Q3�m*P1m����g����-�E,��r��c]�SL}L��3S^u��lf�B�O0}7=S뇱O���h5=H#�l*ݿMo@]�u(�@��ad�?-���`�kJ�_����eV os; t$\�8��G�z��o[�6Q]���=�׼d@�C-C��L��8 #�%v=�;�����e�����0_0/<a ������Ix	�?BO�/��B��v.��t7��Gw�}Y��)�E��c�ڐRW�Ea�ڪR��)���d(s�Ɛʪw��:��.�
�g��T	��2��L��e�K�2Fڬ��J���O0zC�e�m6L	����~KZ��O�����@��)*�	=�md���� .�,a�w2�^6$�hM����i*	�^1����j@�I�[����'�(^m� ,����]�!s�Y��)�ʻ�&tggyS������P[�"�*��>��R���7����b��z"���I5��蘸���o�e������74�@U��U�;��{�X.#�wM�AZ� ���������p�R���_��I/a�b���^�@�z���.r��h(���|Z���<p�;q��*�����TʪG�t��Y��9d���C�����6�J��@e�:���DK�&�mL3��X�p
�_�&>>�0� ����G�"Ǡ��O�Q���&�s�*���|���v�zi�4��Q�8r��\��q>���~���eF�"�����a����#T'8@��Fr�}�.x���g�;:�Zt�tUY �te�cg���=4���ظԤWd��U�9�����5Ub�Ƶ��5�lF��w�ɴyBP�Fz#P�	4��m�=.�=�C�}e��?�/������zA�r�\:2鄥��]΀ o�[6!��L�B�|Ԓ��_]�A�2�y���'и�:������`O'�]X�޸sɏ[�AX:�� ~\���,{����UM����p���X���YQ���D,z�*�(a�n��w����O�����
�6���A�i+k��_�<dd�io�6���	�a�>�7�!/�I��;��HS�#����F� [�R�[���G7�^C��(�b�L��"*�0/� LAd��R9�uL�Y~}�	nt����6;�.��ڻ(�8��[F������Cz����n���EXn<߭�G������YD]lZ�.�i+B)��ɋ@զ��O]�݇Wk�u�-�x4n�>g�n�[=�ޥ�T[K�.��`B����0f�O�<���/���A��d�C��4|�c���w7�Ԍ�+�>��^	������̚g�߬Yc��r6>�A6��]�S��ۢ䊓�@�6{�QU�@7ƣ���6��H�T ��0��-lHF�zE���-�o�>���!��×܂72��qǫ�;�,*�q�"asQ�OCWli��?��h?	ܞэZyn�Wp�k]׍We���l����hx�c}{�|?��S�`M��\�V����G�Y�̲k�;��	���S�2�/1H����� �H���~оUe�,Z8���Wq�O�X�LJ��X4�;e�|@H:&�)YO4��i_������֖2��<�i)*�S��@W@��%�������S���C;t����:����m��Y{+FV��w��E|�xƼ:��ٵI����y;J�?
�^t%�ly4�V�
�/ruy�H��q���^^�Q�U�̰�9��A����Er/zM7�F3i�T�)KP�$�]~�P�Jf�q`9�N���t�����ڽ�'c��;�-Q������}{%���;���CKH����hć<�>� p �sO�����_��r��z��V���U6ڴ頂-��N�Bh��������z��%p� �k��-l���֦���:�i�^-/���B��Db�ۀהǣT�n�AO.�������7\m8j�ѐWFS�
������x�XcXʳ�?�22��~;�y�6.��	A�0�~��֟eX\��d���)�lj�G��-1R���<����uSh��yhN ��;�mSF5o��з���xf�O����y`@D3V���/�V��U�(8>ԊL�D�-����<�H���g���)�h,���@ò��8�!�Ȩ���m�]D�s ɴ�͙;��f���5?=����6����&�c��(<'�?b�s_���l�'�/d���"#�~CT�R�M=7_�T$V�dt"�@J]������膁�|T�CD�S��Q��mH��@p�E�w?�Б`���3��-om��5�r�/{I��3����;vJ�R@$|t��(+��z�4`Ab+L��_R���l�j�V��h�8^�O�!-U�C+:���u-<��4u���ſ71�H�;����t��&�g���W�v��.c�2�J l�׌��肾E�lzС�U�}��`�5�T[#Cp˒p.U�x�oESԶ<��K`���jd��+�Z��,�*���i��
da����; #�FB�K`5��>�����C�l"jf�w�����.\���j��3(j�=OPQ�E��6O?��үq����~���BZ_��+'x�C�MW�R��O���(�Ap�u��a��9��������x
|��|Ԕ.�J�
�>i_$��a�����~1yO�N�q��]�p������]B���qBW����b�gx��ǫp~��,8V���y-X�-_U��ں�]
Pן�6�EwH��K"5�ۅ��@O�>W�"��e��%�����~��pu�� x�&d`����OxZ���C,��N02B���1��t�x��P�MVL�J�Z�j�$M옼�1��aͳ�X�&d�:�z�Q:G�s����Έ]�_��z����w�i����c2�&��\�\���Q�\�c�X���>t#���0��e��l�g}8p0�	?[�C��XL��8\��հ��<i�0�d�̳2��mQ1p�����?<�?�7"BE�e�/ȷ�]Dϛ�>�%���2���֍�6CN�UB�쌋�KU	���_]�o{@��d
̄YS<\�pA���8��`�m����w\�T��n=cV���U���� YR��),�85�6�u��y��ܪ��3$��aA׼�����B#7�\�^��@����J��BG'�����M���9�c�Qd^�����ٜol��Uܱ,���'����|�-%Z����5�����˱1�Dr�:�gay'�m�r�<��&*�']�N�.�ٗ�2�\U�z����wL�;�igsnI�K�G��/\(�¤�8���%q"�I�Y�SOUz=�]/���]\#1�Q��A�ub��T ������K�Ȕy&-eJ�'�/H��^�������0*4�N�.�#�4x�����	�%�.{�c��E7F]�v�s%e{�E?��A.�:y�5�e~w��z�T����3���ꞡ]Hu<��w���&� ��*ʋ0�}U�yp9�)}S-n}����@�9Y☬#�XT� ~H�{w�9t�̾��y��Oߜ��Y+����f��0c�~hj�>��t�_+��zc�|�z��4�3 ���r��ZW���ܛ։�R�:�Q��P�:����Z��OIK�?���+��D�*J�_�'pq��-23��#Gb�L��=��Dq�J��/U��i����lKqƊ|�����o\�Pw�%IR	
�}���S�w{n��OH׿^�ާ9b����Ɂ���}�X; ��Q���ב_�G��?�����c��d�"(2����p�@��j���ȕh��GY�a���\�I����U�#�,-Rx�ͪ�F�k���%���`N���A ~*,����4z����.r�E���k�W1� �2�K��-���@{�P� � =\���dIT;�(UReB�oeᦴ~��c��d}`Ŗ�K{�t�Lv:ۣ.��vfT{<1ra�c��;{�Q�W5چ3��%�Sk��.h�� ��I�_~����};9�T����B�����F8b�!; ���j�;��Y�sn�P���$I�:X�� i�	����+������k�4�⑞mįh��Ÿ������%�6{w���Pbt�W���l�1Px2�(�"R����a���>>����[�a�4�����(�p���?�(�>xE����k�M�f�̽N،uo����ǰ�� Q�J	�Z"�]@MP��[C�K8��AH��R�
R/��,Q�ʹ6�͟X�k�v�˿��m�$�$��V�ǜ�aY���p݈��_ځ$���ӿ���f\h�C$���6;ڮDJ�	� rǕa���7$\P:�N����e��c�	sW�vh�u\DH����Z�٬�(c��Y�L-d/aa�A�(��ԚRߗ���/���ON�64^ti�_0ii��zb�Gizn�'`�J�c�Ҷ�ț�"������j\�����w&#;Nv�����-/`L�ə-³�tP ux��Bd{d�.�����C�*��'����r�l�[�����-)+#}�	x�Ey���x�K+r�@�X���m��;��c���T�°��:p��M]�T����P7R������6��X<�������ɫg�m|4��a��> ��*��<cqP ��4�o[� gw)���GC6NQ�x�G`Q��j+��Pp�F��ƟJ@}D]j�)Wu�|.����Ӡr�KɬV����ܭ>�A �������3��lIc���@�5�кk�ńQlvR���_�<��Jl�_�W���i獤ۖ�I��-�	�t45x7��*5�q�n�9�e}-��+��ֆ�bT2��\��U�. G���zwư�d�Z0H�>�x��L>r
�O��]񞉢5R�wG��4M��rE�Zz�kj���;�N���%dE�Nl���3���܌�.w9�$����M�H>�v1 �ם���IX�x�"��������;W��Â�D4����·�ؔd��8b?��yɽ�ϫ��a��g/G�������i�ƅ�f���-�G�Z� _q�~M�:��_	0�)1{M���]c�|V1�ߖ�����EB���`#5���J�8��o\�pg[�&I6��,5�^Ṝ]�;�2��}��_�V�0��.n�=�ei�h��):�Y*RS3w�B�`3�n�Գҍ�:�|�U���p���@�N��.6���/lo�N�5@�SD�9����R�Uw��}Rr|~�%�m��wO:�Em�,��Jvi_��i�����$�z�}ڛ8�4����� �}�c4�RF��T����/��E���S�e"!�?�7G���B�������3�F�4����8f=��ֶҶ!�{�*��=^���È�0��5S��&�Y�P��C�u�v��Ţ04a��v�`�25*en��H{`h���ml��fG:��bq݆?���s� �Z������,�c=�GIN>c �K]����!62,�4���zAfq��`����c�	����MB
gf�i� �����A��}_MZ��?
Bh�������󤌅 ���uL�Ͼ��I�>Grl{�%�=�sP�>�ozB�^��Kbe�Ľ|�#"�p�hHxE�YRaH������'��^��d�x/XzփP�G��|A��"��?fW*��>o�Sqh#�孨�3G݃ʨ�/�4����ĵ��zI֝�Wa�������j"p)�Q%+�L$FI4�"������w�%؎9�ۘv���e�e�����\�0Ϥn��0%�F�;:���y0�����o�ի�	�pۨR�W�E�r�{�)\�O�_�[�4,M/-!g���P���>}ʭ,Y�͘�ki-
���Df�d%�%O��*���Gr�և��J�F�T
�|̠ODI9���"�*ÖB���+g1�F����v�8�;H����HN��Cy~A�����yBt��*��i(�� Ʈ�_��w�g}�z�8�಄A��d�7�xc�"IP5�I ql�Pg�P�=���Z��|ȥ$���$X\�l����O��V`9T����l ��)'�[p�
d���F���̣̋�-/��rdq�-��vt�L�eod��1a2�;�׾�#i�@�D�?h׍���c�:3 �!9Qߋ���u�̧#�rB�z�㪾�<��U}���S��w,R�EH*�<'r��"��9h��W�?~�C�D;�����`%Y;��9Q��&�D��=]Y�F�=�e_ �d�ℋ�ˀD�b�J ���E���4!fF�r#�	��r*?=���܆��@���6�O�G�ˀ���K$��w�Ve89���������kꙬsҴ=+���SA����K�m�%�Th��GD�3в�ċ�՘�&5hXY;T[�r�����b�?y�K�2�>�r��Mz��%�n�Γϕ.��>E���Īj]��U�(Y�<4����(j��~ٯ�ɍ��P(#��sk�}�#��z����H�P�� ũ�z�hd(�F�W�h,'�:�ó�/e	/!Yr�P�� "}�̫�n	o C�򃫶Y�}�:��쵙6b��5J��6���-�CK�D�$�.���Df-��J�AH���ڤ2�(��xݰ�V*�,Hϲ��nh��#:k�L m�6�9y
ă�7�)�XS�!?�\��^�,��W��ɖ}nC�E�7�Z�JZ�h���hc�:�����8ǁ�_ԑ�������7�B����4�m�Y����ʜ6u@j�pFi�Jg5M��'�2��^d��KB�c~��+��T���p1�Gl-�و���Z�q(����1<�$g×8�3���f�p������/��}Aе�d9d�����d�h�P�J����%�۷�\�tof�v�ͽ]k���w󆰤6n2�IȽ�oy��k�k���L�}8�5Œ�tK�\k�~��'��k�fm�;ڵ�\�\�e�3�YETS��NT�����p9���c<�!���I�OqzI���!{X��[�����\ӭ�rs��'�U5��&�b�F�g�)�)�k��!�c���1==���"*~!�=ӭ�Q;zڞ8��:���; �/�C{�A[`t�N͌EӾ����K;Q����c[S�sDG�
�;� #G�㿘G��8���y�Qf`�h�~�a��Wk�[�:�r�X&���[��������LB5D�I�x�羢�_5�FF��_x���!�B������_܃��h�^ȔCJL�*��5��[[Qȋ��{β���A��b��O�檌߬=����i�� ^�mq�#�S�IӈX����ޭ�ˊ�՜���v��B$�hV��UH;��lxoK]�#�s݋��@+P�����n��B"���ef�O ��&�ś=�5������T��vhTVL{5�����h�^g�X�:�8��D�5�K�j�%��t4�c��m��a�N0�4?Q�� ]�YMIr]�y}�G�,�~����2��[2��o���-8V�}��]�$N�o�E�(��é��j^���K�I��\b��!��a*�:>�7ks�oRЇ�x\X;D�dvR�	N@�3[ٓD�V��m.?�X��[���9I�r�)*Z������G����{�E��鍙�dY�D�Z����2��QbBu�E�;�x�4﫣>\�^(��[���H:pC�{��E��r#z�FTQ 5�)82J�+7�G� x_[����BR�"׽�$�1���o4^������E�D��j�����P�Q���1��1���#��N�4�\ �e\��c�0���d�&��ۢ� �^<mךA^�72@��j�	�����!�E|�'z�2,t��6 ���_�i���e(��e�?v���z���EFſGk��3~��;M���D �'/�U��6^�um�X���s^��0��@����Qq�%�ZT��R3���A|�M�7�.tpI/	��mpÇ�hԗ� L�TFy�H���;s=��k�2.��V�ixՏ}!
�M�ڣ���]��؛{>u�C Q��Ǵ�j�#~T���D]�s�~K�ċR?C�F�Ю$~�����k���b�@�?�f��ɀ�3gs�,����L>�zGH\��zI���R�q����*�'*	$M�^Cs�5Τ�^#�pGj��^���n�<}Jg��5�g���o�f�����^�.�pM�����}�aE~B1�J�b��#�n�r,��2k4�Ą�Y�� �A��M�Ψ�[���(c`h����Ӫ�7!��	���%W�ذ��X�k��-c���I��!h|]ۭ��(���u�؎X|�7O;��4Y��ec'Ez���c7��\GН&KT�,Ul�6�	 ��0۬��?*�R���1We|�/��d���J
�F%sV���ҟ^����J������HIM�`s��Vla��z��\'*$o������=w���@"��
^��[B7p�C�*[%9�E4N��#��ȿ�0� ����/�G��D�����1�"�������@��/�\�q�|?�K�荰g���ոDP�G_�J�9�w�FC��M�} �d�i!�}-3���lM��cJ$V�wE����y50����&n��G���3�=��f�i�t�Q�R�t�9Ga<U�#T?� ��uy�4�2*����̴�����K��hc�H�3τ8-�d5vA̮�]Am\���j@h_��4�v���R�є�9��^	S�gW��2hͬ�3]���t4'D��?��2e�ʆ�h��_������X˵%�X]<�N[��ή�ۨ�{A҇^m�R)#�F������k�~��pL?h58)�0�/-��<h"�/��D�NYH\��tr'SP5������]�������tC%���P#�\�Y��AB�&BJ�"Y`�(�5���͗�@��z��H�&�xcec����j�n����~� ��q�	�LT���?j��T��(o�媲n��U*
q��;��~�s�%��P8E��s�^	�%�M9����E�˨;y�#��Qg�đA��J��Qj�x���a/% D��n��@� 9kZ�;3[e^=:��.�@������N���)hY��>��_�.��q_暔�ia9�n��S�,vUo�[h�|`�BEͭŜۦ�����o<�?+�o�"���em��@Hm_�:�Z{�WC��3ȼ�C�_
���;݂Y�{�����ߜ�?T��y��ͼR��A��hmp;з#�o3������M���^)Ĭ��*'�l��О���&/��4]�$�S�D$�iϛ��L[��_�ґ��e��&pB�N(y  �
?FM�<]�j�t�N1�l�"�{uk~2���T�	��/?���� �G
�m�	�Y�8V��#�J�-�s8�ځ���d�ݗ�gq�V�=p�L���TZ}e�C2��&!��9���w�eT��_8v�C���'�K���n�K}�rs�9�1. }� E��pg��u}]�X���yW�v����"i���3�Yr7�&�	����͢��	�Ɲ���.e;�CŃۣ궎��T�7�Nf: �Hӊ�#H |l�|ʸ8�P�U
�UC�e���Hz�0�����,�
r�r"���t��P�N�i�6՝F)�کM5:�w�|}4�	�n�0z`�g�f��?�b�_���]�����k��n��s����)%���y�U��� N:]��]��<�$�s�~��\��(O6�M`Zs�*��mVC�AX,��pYw�}J�;ȇ��Jt�lR��c���3(3c���aDW������q�����,	� ��'�U��c�%����B����F6O���8*��ߣ�W5�wɸ;�K���8O+>�(C8�6��e�2�!4[���W��F1������f��T}��#�X~���t[^^�3��m�+��_q�+ˣY폪������q�3b���Ni���l�3W�qI$nif�����-�#�~J�=K>�,�v��
����k�l#����d}򰴦��k@>��}^�ׂg)�R؞VT��B$(��u��',T�)Q	W�>k�f^tJ��q�G�\��dN�R%�%��G?��Fa�{/����s5��*��{̪��|Sʎ�m�����=�1����zZ�ؾrB����`#.Tx���	��������	��;2 k,��;S<(-8���2jQ1�S���ihs�K��;��C}4D�b�_�w��!�jPd�V��Y[=�Ù��#�(����+��|�}�!@M�/��[���p�=��͋��;�1�W&�-�мj���ZbO1g�X)�+�$��vě�]�.�{o�<?��[�_{a_�Um/��j����Gw�+E̠u �ՅӰ�+@�L����A���,P��+��ȅ'�e���-��٤�q��6��2�n��^���	�@�gA�T�I$�WJ��nE36���>�	J���������9�P���Q� i����\�E?�[Rq��Y�x����Y�}����t+-�(!`�*�6�C�l�����@�{����sj�%Z�)l��vMʫm~i��o�g�\�Y�r��w|���ߓ��
�3P3"�"o���/,�Eߑ�S�yȬ�%z��s��U��!������ �p]���l>��J�V�}w�kZ�3����푤�7�����O�G�:jb~"�n� �&�OAa(l2�C�>�Vʢ�B�;�sU
�����H#�b�\� "e=F�)2����Ȥ�/fZ���;��T��m+ף����95MMG�i]�Vj����J�>עa��B��o~2��d|��^�t��o]���vr1$}��[Xx��q��YJ8�G��r<"`[9��q����=�׫f�������«��㨥�dcLU��jK�(P��݁���r��H�a���F�I��W9�%'㭝��1:F_.��"m��,i�Y���5�������*��(��g�H���u_�Н�Eu���������!Z����ZiM 3��P���9��e}3�`P-��}��zq̀�H4�)�d�%�|nDNj�g?z�C1&2��+�,MlS�;�o�myn���
xJ�G��s���w��K�d[9!@w����p=��Hc�ot�n'�B��c&�5��-�73VQ߂k���6���Q�b���x��ZO?ܼ)�N8�SSM�c.�IM~^�q�(�X�V�n0�楆�G��Lt�����l���w����v��_㑩7?��b����յ�+1ә���e�f�&�Ҫ!�"n��	���
B��ҥ��hCQ��r�V��x*dԝKK��Ssop���efg#լ�ߣ�`��ж���&��u{�n�W�1����%�S~��9ՓM-H ��06B��k'�!?[x�'�-ʝ�w�<y�S�#�`L�$U�J�����o+���\:3��8.�OI�ܵ��Ӿυ���	�����-���껕��-�a����6��5WW�� Zd#�1s7g{8�~�K��_;�G�wк���8T�kr�!nY��ԘMPr�e8O��� �U}�P�K�P7���L'LF��/���n�H�d�Da�Lx;��(6�����Nf��Bm�f�Pڗ���O����5 �[z��TUlk��Y��I.������f�N��d�@���5#����$B�s�s��! 0��������� #������:jWE�W�gm�)���)R�Y*ь����NQC�w!���f����С �*��@k��<�=��))���I��>E|+`�����{Q��p5Zʺ�I�6��m�`z�k
iNA�H�܊�d�]զ��-v�UG2�Pr��%�wo�̬M� F�R`�:��5|]|��յ��h��
�1��kd�d�c7�v�p�< ��n��[){�z�{B�e��Ĉ@[��5'��ׅ�7���#?|)�$�𸸃��-,=���^.�a�4@L
��>�д�j�����'�x��ȊFe;�!�*�V����G�.�Dx�h"���0��t����+�{៚{���Xq�ԃ��ME���)��Q��S�`� �O�-ou5��B�$=�ª`똕�>�u��ɕ5x�l�>�s/BA�����΢zlx��u�f�RNI+��"n{t�W��A-��RG�Nz��J�~|�� q�p~�C]�?�st`���B��u�B&�w��uل�yIIR�ܮ/�j���9�h��'؝T�ב��{b�Z�5�{[P������O�	!~�����D��߬�^�_Ƨ���H>����g�>��#a�KNo��\�i���	/`�^�P6�*��W��saX���)��
����ݹ ��|��J�BJ�����~x�Kش#�����"ݟj��<=�>?-A��_9U�h^�h���}^$p���k��*rtI��{��u#v�Ž�`i���I��8/�7�x)E|�u8���a�f.������&y޲�W�|��♵�!L���0�R��η���k7�8Z$�1;c�lFU��;^uh�ѓ>X�X��~���}Ϗz@���:^,�XD���!o��"V��Kv�L���'�&8�v��P��y1,DE�q�OcO0S���2�:��zR�cޫ���)��툕���C���p.��7�{��ǘa��u�/�t���?��{�MH�`¤;��u�F4���-�� ��6�� I�!|���h���=�����B�~�O��3��5Z}�m�y��<5�g���O�.�% ��u������a���z��#��P�����$>xe�G��`�����ƚ�	o#Z@է���U�G5���W�r^�$K����S�I[DL�*�<������E+?�S8�S��ߢ�T�&����-���t�@���ݞ< q���C���;�xq���5�}j�v�Xd���M�9��Òdpto4x����wRp�4~#�
�;����/ne>}&d�|a��2�b=�X0�"ck�����/py]�_���W�""���E"�k=�Ho��$�L�����vc@j&�}�&?�4��W�s���#�B@=\�8s�%#]n�?� Z�Neq��.ɴ��ȹ%�L�DP�=S���{ݴ�v>��.'�p��4n�4}�[?��Lh��F*�Z��XW
m��:p���ۍ�c�؂�G�N5;�e0��/]����m�bq&M\�	@��j��q�j�jd���:@F�P�5h�S?����nį��� /-/���D~����d��[U����G���	��g��*�Ն�ՓHm9�,b�`�T�����k�pR[~��� [��S�šO���i��!~�@JUӭ���\H�Prd��({_�I�`���Y�E@IL��F�q]B>f���R>J�Ŗ�J%Q��!NԠ�2�a�{~"v��"ט���ÝU�L�[$���`�JR>�^Q%�t�y#a�rք
a�ɖq��Ĥ�3��M�B�XNU�`f�8����������x�D���}r3N�t;9�!;?L��SnB� �^a�BP-�
F�wb�Ӏ�35QFN�;bz�(�����Ӧp��� �ۯ���*
,J0�T���j|�������%d"��>_���s^���OQ6k����~�ugzw�Kw��c��u�b<5p72�5E�us^ߌ���7�����x�\��߼7�8����30��"9E�}�����g%x:�K��^K0�K���Y/4c�kGR�5]&�
?��M�}/m��F.)�..���R���V(��1G) �:���n����3l9n�o岋���~=�S���?�A�x���bz�?	��aʻJ[W7�����k���U\�)_�+C p�\��@�)����>��o\<�$�d��V�7F�+��e�N��2'��*��4�=�}!q��~�;'��K~���� vw5�.�О��o;�!/��)��b���-<���òj�c���1�\�EWD�����<#8��Ŭ�m�^�Ȧ��g�ӲF��`�Q>e��#}P\�X�ww���v��$��=���83���.�jlq�C�7%d��&��=>�z!56�	����)��C�W'.����5�C|䄜�ld,�Ju��T��_�^���'ӥ�Q����\a[Up��xH4���@C*X�=˽t�c���臓�<f�@r�4���V�Z� ��l�1Uk�.p�Q�f�\+�2�� �I+;Nh�o}��{�A{�Js�q��� ��r��n�:��@E��ؕtO��B��5/|>�TT�#H���(��P��������-9<[�'Z����;�H������A4eOGߊ�sz�Jӂ+t�'#�#팉��j��J7��0]���d��>z�.��J��|�b��K���R��m����������a(����ոd�aQȦؒ��9_a�<J��M�R5�����u�Jf��V�4
���>���{�@cbi�8m:*3��=Qo�B���� :i&��� �v�_�8�G6�e�6������]������-\��A���rx�K�(~9�أ�`���,�V۷�g}#P��7{v�i��E}����R鳵v�O�'v�����Cq������VyQ����.i�$a�XQ�a+.�����������y�(I���J�,Q�� i4���4x�f�P�"����K7l����_#᳑���p��C�\��ӻ�ԭ2ll���4����߇+K��<�}��/'���IA[� ����j:$��o�#]�y9�)�sZ��7U9�R���c���A��'ݸ<�%p1�D�(�-���p�H��oُ\үi��-�����21��E@��`�2L���J|���@yg-�~�"��9��n_=�'��ךB�T�#+T3)�6�-��o[]gP��f�ӆش�p#�7M_�G�7R�?����`>#��0�E(��J���z�������x�9��K"��k]L�\�'������yU|"�p��)��2��рJ��/5̼�g�1��{FPz�$�.��+K������ޖ��ccԭg��y���L@�_O,"�G�,�|���ԁ��)�ٽ���*g�a��W��,C����Y)�hd̨i��!�������h��ߐ�Y���)�)���v�$,1���BH�uj���=��H[SmC�3�̾-��;��}κ_��b_��-	�D<���F�e�$��8
L5a������_m�f;��qŻ��*v�fp%I�r1�h�d6|��Pr<"C�m(޲сU���X:}�J�?Jr3���2O�(��\D�Τ\Y@I4#��Mɑ���� 9v/(�GԢ{g*B���_��o&��]��4�Fs��!��?}���n�Pb�:����F�\G�5Q/�v2���OQd=P�YF���fL�B/f��+��X뗇(�k�A��|g��G�G��:��:6�'KEx���	W��7�ԉ�׃G��.�虒v��j������6⡺��$},�L>q�*f�	Wy����D%�b>vbJ�O	H`n5E��-�.�����_��Ɓ,鴌�x�������5�Vb�����ܱ�[�0��Ul �c�$���(vK,W����`�e�,*`̞Q�M����7�cԫ����YvT���B�R�V�he�� ���&M�/�n�+݈��/��y�3u��fr�Xq�ݱ�nIY�t������P���pJ�5RD����جM�
:dʹ��~��=�41l��Wx;r�a��(ZƸB1+���v�%��3<�	���lej)x���h���t�X6��*��:(*c9�p�z��K��}��e2��l�U�$;�wy\j�=j��p��z�hu�3I�p�ia;݌p���jh^��a�5�u���U�7L��?�M�$�3XV��p�2vT��V��6@�ޜd5I]Y�B��^����,O�7�tG^�Aq_#|؇��(���y�P��
��g�C|��oz��pG�����>�>�X2�K~���h�^+gZ	���qLE)(u�C�a�D_����ᆑ��iOy�+߇rV��Ⱦ��w�����]�7}=��8Bc�� ���\��ڢ�����/u�>KEug�M��y�(D��ϵs�������Y*#��w�����0kt���:�'�t@�xw�%8����j\�1�0 {��(���qYK��9�M^<�%1j/_�2�=�%��#i.�����V>��H��3�FL��kW�
ġhĞ� y���r&H�a^8�>$}ŠOj@�8�����y�A2D��Q�����Y9@�"��]D�Ф���l<�09:�v����QR\T���:�o`�6����'a����:0}æ��P��� )��I��	��_��mt�ʩٝ�:ҨaMP:���4t�fmmp�5�S��s��(�<TC@�{���n�2��M]���� ��x*C������^)�C�q�_h^]%c�O��r�u��@�.�DjL�>�w��X��ϱI���	%��ku���Ç�W� 8#@�s�^X[j����?髭����4�*;>��fbnNt �	{�m�0����~ʀ��7{WLh\��oc a��&;����~�`����Fj%������&Rҥ;{���aӬ���$O�;�b�ZOǴ,����Ҍ��x?�L�3��w�Z�
����`�{�=�����J�V�OTi�˲��e��9�7��a5)4ۙ��'�Ǌ�-V��iڦR�y�,��⣆7P�i7k�ң������*�j��;�F�=�n�޽mRσ��^�Rѿ�Bi�;�RlO�H����3�T��Y�$�����g.L����LU�&L��qN�佡��^Y�����˳=�z�ݗM,pVa�G����z����/$�Nx��t-���e�����!<M�6-�8����=��Q�Tw���TC�ʳt��y\n�g��aQ�!��0x_�O�	����m�8��j՚��D_X9�����Vh��w�lZp�>�~����$�b#�1\�&�S�#� 1X3�%�R��9R3�? ���것���d�W�����k8�+�#/�.#	F�\��[	��������>g����ߪBIta�DM��W�~3ڶ�v�:�z⥓�h̐��sY��������cu�p>_��&f�Jʤ��.J� ��Zm��N�M�5�q��sw3�_�1O-a�n�K�#�D�4��[G�{�bwEQ&��
�vk'5b�j_�&Vz���(�|�B�:��%C����{r�}�����c4)�-;��ꘑpR,�8�܊r�x�^��<��V�ֱ��q�o�ԑ[+����.z=?����W��p�_���=_X��J�nի�Xufh�<`�܇�)��^q8�Ca��PrgȂ���cS.I:��~����[��i������$��{��$�7�-'�3s���C���B%��+!��p����A�;HI�龜�����H� �8t�pI"J�3�>z�8���ݑù�Wdv�A
,��ۿԮ������k6�(��M�Y��0� �e<�>�Փ#�3͒jy�����z�>���].l(T>���!nL���K�v�Q��d��|�㷞�ip��IK��n�����XS�4���sӬ����Ib�$,�k��2���ø|]?n_4�D�[�%#Z�D��)ߢ��E=���\�P��i��`���<�YG����'k����7>�6�ݩϛ�+g��0}P|\T�ո�s��H����e&���i�y^5Z�<EV,2BGq≄X����S1��[���t���9*�됯
��<f���DE�h~6�`Zd@�v�QOdS׀%Lc	l�>�י�d4�$\��p��?�wuT����/I�0e�Ԋ���*';�;����(}<�I�H޽���=�Z���Q����~z��:��. ��`��FFn�W���uј�E,H#�A�g�ug�r	��\�`�pĜ
뒛5+��EX0����jI�TLCE��ȰM�rx)�J�mg��A��	����E/�a6Lp�W*�J���`�9+?�g�޳���-I�{ �	R�ۀ�å�@���[I�Q�Z���}R��7h���]\ ��y\� 7��n����f./hK�C��O�o�A������Uח�s���Jg0���6��� ygl���H*�!=��(��iMV�i5��e����%G~�2~D�j�㪔�n�F35.NT{��A�����4���!'K�B�z�g�:�� �~HpDЪ�LR�Ϝ4|��� 9y��-#��6T0�7�L$�R�*/�Yv�U���/'�Bs
sÔ�u<At��nv.��EO�{n8�;6����Xa�����r���Y-�(R�,T���9
%=Y~��Ո���>7��(�����&&X��v����L� �b�_�ũ^DT���݊Z:ϱ=RN�Ǫ��<㫌������Clf-�y­�E��5B���V��&����P��y/8V�G��P�*R�*�c��F�5�I+�Ipm�r~u}n��p�O0d��������R�h��b�\0����CI��a1�@��hJ��'�6�ײ��}�~YSO��lP�h+T�)A����ĺ͝�	@{�\����j��Y�`)"�+�f�S�[��TQE����� ]�t�f������W�`����A� ���}�Țé���7�w���ߎTz�� �dzG�)>9w,�	u<�ߕ����JQ���!D���ӺL�%�L��
��7�A�� 1�G��H8
mZ�c.Fk��MZ�e��h �檲�U,���h�(w���^�v-���#��gV�EbԳ?�Ď�z�?���8�v�mu���L�"c.+� �<쬀�TZ�&~���l���.��>�ͮq���qW�D�Up��^����i�&�u��r<�A�{䡾��J�r�b��Q�UL���+� ��2�vC�lØ��(mc����A:P�f������>j{3��S�L5ο���C$D����\[�xr~�6W�I�^7�פ.g��ZU��+,�O.��s�qoG���!Z+hBdo�M����Q���x�$�������\B��֋�j�t��z��%��ݜ��FDa�G���2O���~�z
2U��-5.����Ѽ��js��C�Z�FJA(��ge��!U��AT;N�N�C��2�My���$�>�|A
�|kRM�ɇ� ����ڮ��؝/�"%pn��� �6ڡ��M�6�ֺ�2����~��q%lnA��&w��Hm� %w�g��� &��'u=��9�?*jLx
����Qs�o3HCM�#w{��Ǔ�JC¿ʿ|�(8�?�}����:ÆQ�Ǒ:rփ�9�y��xx�(.g�b�C!Uuǯ�/���\A�#f��q������#�� DEՔg�i�c��b�`�����Ɂ���U\f�m�I{2��t�x��r@���$�����m�9������Z����őd�����nf���l���=��߸]��(�v��)�,�hKE䦹H��V�VYy[�M�C�!�c��:���دt����N5�O/8%�^_N:�	�!~�"*� ��k��O�'���bWl�`��B�K_�ф��rQx����h܀2=�z���k���讽μ8Ϛ�$�7��J����X�-`��(���7�N����Ӟ��;��*�0�2��<��ܹ�]�@YrMVU1ѩ����e���9�~IT"9$"��c�ZK�DD)Km%,��$Ie����0iAH=N-V�O�ˉZ�P=��ݸ��C��Hf���jf3#q��L�P�tZ��;&�,�8�sH/,[AĢM��/7����h�)��]$6���P��a�Jש.G�&n�6k���D&�>�`�'��_��ȦVN���i�+�~�?U��;�A���T�3T��\N�ylo��p3x�M��*�C��X�ȡ*Q3���6�Ђ��f���e����~U���^e
Dvމ�h�l<H��� ���}�3�2sI�H���8[��=M�S�E2�Z�K����֬^��A=�ᔯ�#�C������L�v��F5�5l|i�Y��L��a0��򂘰�.:v��g�<�0��_�C�/�V��6��9c|]��ж��ߣK�_M�q����0y�К��Q���]�DZ���@E�����2͙/	�P��p1�H�B�_͟Z��� s�զBc��>kw��V�,�7BA4���Y���t�=�{���R}p������U���c�ݠ��7)<���Cp�LP>ͅ �R&�Ӎ�k�>�� ܓ�c���_�ڠ�K�p�&8�o��^�q?C����խ�3(���S?��Nլh!"W�l���2mII�`�>�^˱���!���hm�hy��9��D�Rm����^��@�q��׻*bC�]�6ƣ�Sz�;7���:9Q��R����D��r����aW���ύ��uqݵwI���LKw]c���}ڂi:+�<6�2c���mY���ґ�(��q��P��D}�H�*n� �>��L���M̹��A���b�-���
�~�-rt�=�h���hP`Ё� lp/}Z96"ޫ&ޅP�)zQ��4��Ր�nq�d$�~�1�ݎ�ˀ�E��F���KE���L��E�#fW�݉zS�m�)ӗ4�]�ϳF�"ұյ������_ـ8Bz�c׾72���f�
�`uĞ�HC�޽<?Ê3R���c��%�����Ԭd��Eʍ����{�?�^������W�ʷ���M�����V����E��w~8B&�0��UO��,�C$Y#&����BW���n�V�� D�V&��n�Kl�W	onX|�(���.�h~�H3։#cL�<٫�[��S�]b����w��tX��rx>V�3����Ar܋E��0pl��W��w��#�7�j_�%7���+�t�Ǔ�e<-Qu/m��h�Y/CwD	���x�-��e���v-�
17�M��؀��$�z`rsh3��W���0m��������E(&_i�@_s�S�h(g�rI����)7��A)󪲊0{k��p�9;|�xO��yj�Y'�c�}�K;u�ы�'�2�����o_П�R>��y�bGÞ�$�ٶ폟�^�+���B�|�C'ax��V?.��yR#Bgr�U�-N��cu�)��� �W�˃��"S?a����g)c�!`��vo]��Y|]�D�V��i�#��݊4 ���� yQٷ̀V�k�zeh���5]�/-��Se[���
*���1��UZܻ��I0��a.&��8L�3������{1����c�~�+x��."�:�J��x]��11�]K���V$�cA˽��.�#aI�j�I�F��Q���⢆���<���X�bu{���b�{F�����<��L��X�Xdb��գ�bYbj��GC��G��k�W��5�߉�����jx�xU"�}���=�D��iz�d��� �;[]�5��XF������I��b+g|�M00�rT-�Йa�;�h��*�(�ld*��Ͱ��{��Jf��@@�A:����t�����\�v��EL����R���A�	4��s4t��*4�3�>��L����Rv�$���R��5�����^�;@�Y��-��f�?V(����~�}�S��?R�s����L�4)bS�ME;�t�m�2�AUf���m�b�.����h����l����^\y�ܐ����_(�;��f�����;��&����.�L�\NK@;��6��Պ3�:C?_�=7�_�Ѣ���ځ)��To�f8g�w�������L�+���S�tU�IM���#�I:��af9`�2�֓HI�����dB�������� [�A7r����P�	�ͻ{3%+��?����`�KA�_��Y=}ġ��:V'��=]�a�1�I-+��>�R�1����%��b��o�i�����x�dJ������z��F5h�;�ʧ��kj^l_{[��#9�>
��:��Y���6��BK+�k)�����]�\���
o'JU-εH���*���0�7�e����R�,ס�$�p �c~Ifwv����0�N���j��_iH��b�{M/
��4�s�p�8r��ȧ{���T5��W/�WU�ؽR�$�vc4b��AK*�m�g��`&4������.��.�k�T9
5��
ۏw'��NgΑ%�@��T6��,.�@�=σ�7_�g�(��v&bw����0��02Z6�f�ѷ��2��Z���D�jD��Z�#�A�ύ�����'T#,	�$�������͝.��������������'D��5�'����O�B�us����{r���:~��[F�Y�$�u�.2r�w�X�S"0�w"��?�T
é�jW���]���Y����缈y?_��,��s���D-#-P��F���T7�}jc:*���}�bF=�� �m��D�%�)��Uc�eH}i3-���e�rf�_��c��/�)'6�D�D@��6�O6�N�z�ǰL� \��7�O�9Ŋp( ����Ai�g�qYq�n�m�Z���@�y
��n�����r*�A.r���冲�����RǈT{�C@����-���Ts�U�f? ���F���y���W�W�D��Q�_�ctN��FZA�]�?(���>����+��N�p^�'OԲdڢu������6�q�,]~xҌ�g��++"����T�Ԏ }���0���ߴ�� �C����'��J4?h��u-N�ha�n��3�0�ā����t-���棿�5\5�B~�NW���|���>�D&���u�y�JEg���z�l3�ē�l�|����Nܨ�bR��턇�4�e@�`4Z��a,]���y���.���%_0�xB����/�#�!�5 ���=������<�0��x/ȩrF�`.�P�-kày�G~dsa�c� �$��=��ϴ�a����!�����
��fɩS0����-�L%[�������@�K핐]vtya<�=�� 0{3�㦗fxW�<Mq�B[�!r�� A�6��6(*n/����<fWC�H���jc��<�8C���ss�諬Hތ?���<x���C)�W	��E��T�㉓ϧ�!��+���Zwuȏ�*d��B���@?�.�q@A��$���/�o�u�W��~mB���,�w��oc������|m�PX�6rHCU9���d���:�Oᚗ��V�< ���A9}�Z�����[��s�m�q�N�����p���=h��)�l�߽6j���F�����r�9D��%��Jǘp��OT�k %G�>Ya�c�՛Z���>x`����s��RqB�S��4>�ʆ�8��|225�չ��G�5�s?]��8���ox9��9y62���Zc���2������� ��(�V@��P3f׼#����?����0�5q�q4��7P��S-���/��(>a�;�J��La�S��,$��#0���55p����if�̈�6��JVg��N�&M�B�g]`�&z��0u���f�s:$�n	��(V:iñ�5���+,�`��.O������y�ۏ�Iz�tÃR���y���Iey��	�
�f��� G�@�;s&8���ٛ�P��v�>�I�x�M�d0i*y�-�,����l�&�ؓ-�C��4�r���q6��X]¸�ȣ<f�;U���s۪��Ik����%��#rD���P�BS]V�|���� ��F3Y}�_z��=]yۀ�����ǩ�t�7�]��xV�y>Jx|�#+T�c·Z)׋vJ�+L��k���mE���l��wR�|�p�d��n���/,��o�R��S���K�ܲb�����x���5���5�'.�𪗳;A�V��7���o�v�)G��f��x�����c�lόkA�B�xMP-_y�:���?�!�A�b-�#b� >�N��H��:J��4��D�Դ��F��*���?`7%M�pݡ:uG�|�lao�w��L̔KY0[a�D�D/�o7z]b#��!&sΆ�>�f#�]Q{c'@�R/l���x�[�d���΅�O��L�5���7�l	�����	]�Y����4���F퐕(D/�Q|����<%&�R+@{�����	��A�.1?��~�"F#z0��v�vJ�<Qz&��C$�����s$ub�D�t�f�*��Oz��&4���UP/��	iW���tȑr0:�RǳG��
פo&	��q����u[���b���<�er߅�[�-l���_�
8e�D�J{�b���k�:���ͳ3->+�Ь�j �[/�Zܒ*|����9װѦ2{�B���(����
D�]���` :]�yO�6KS�44P��s��JA�,�X�Q�%��ż�h�R���c�{�$�=��l[��kƞ��do?�,�E���fb��Yȅ��x�'��SI��O�m�9Q�Ұq�jdړ�3�m�Zc�k����?䡭2��w&�1�ou��_�e�+�輩���Ux��-��(!{�����ܚDY�4�f���_8{w+1{�B�T~�_�	ۮ��[��e*q.��Ir�[��ˍ���$X\��Eq� ���A���GnS?rb���j4��%��zv���uB�w�Ds��*��;�5�cҡ�;�M��[��%�8�d(��ۗ?�]T���.��jb|�%Lv��>B�]���h�SS��;i����M�H�aƛH;� �;{дI��v�Y	�x+�Ag@�G6:�V	�y����"�:�-6�<	IO��������{�ZЁ(&HS²�w_^7ӹ��k�Kj*��r9��
S/wZat�(� �h���9Ul���s���1���Fɉ��:�ӣ~[�����%E;��c�)�^F(}�M9���X�
�v��~�m�È�0T=�%ӆ��ZwТ�
/������HT�9��"���V1Cn�n��}�ȩ��f�w%]�-M��"��Δ�m��	q=�����G��6�k��#�//�#��:;q=g��cwUE�Ft:�J�V������*t�3�k�%"5p���*l���ZVc�vz*��m�i�Mp�ژn3a�3{�镛��"k�-o	N�����X_����D 
�M�r�Yȸ�_r��s�b2/4Cm� t%b�����5B�GZ�R?��wa5h��M��< u)��C����g���W�?��u)�Z`K#4<���k��Q)(��!�����¯��I��|5��-���=�n���U+������Ntܓ���&v��#ש\`[��-v�jUH�8�gI�C#hF�����s��m�\��R�y{l+�A��=''bS�U�����q	3�\���*b�҈�����bU��S���"��Oܔrt��gyED��b��"g���<v��(��).'�M	J,�����y��_[�v��r��cK�zG׋�m�������n"�?��*~�������[&շ�`�+g4ΰ=�~>_�ί̋Pَ���� ��n�#a�mM��%{C�w�� tۖ+_p~���%��@�o}Q�����0��on��z�7���)�0V��54ym0��� SE���c�7}�Ĵ�9���~����w�o�G�|�w~�S@�lr�-L�Ɵ�������8 �Up���6��]ΥQ��O�a.ve�f�rv:��EB>���>hn0��5u�-P��mx�/��IkE�Ӥ�	��gj�i��R����� ���y�W�k�j�ۧ��z����-%�����L��6e�@�n,�Ro�t>f�ۆ�Z��{�ޙ3�2��ت}�|$�]��r��#�K|F����Ô�<:0��#�1�:[pfy����F�"���bZL���K|Ӫ	$��|�L���g�T���N@B��s�a��� Zƽ=c����#Hn�&���gpw����������p�gg�1:E:x\$&�R�~G-Ǣ��n�a���JsI c���s❍'�����K翷�޲�n�M����_�aa��l@�{�����չ�GaE-8~z����	~�A"^���8u��ɱ�w5nQS�Kŀ���hKX�:EQ�N7��'�������������e��p���LKԯvK�3�l�f�=.�k���`=��aȡ���a�ב������T��:y�P'���4��
�bl�]�V\ff.T<vD�M���,l{�OZG�r'���%�S6ʣ��?C�����R,��ml�a��?��%(?���>�:K�����Lm�%�8��ĒO�/��2LvZ�ݳ�⧲Fp����_���o�y�~�ajB�4�v�I�e��r��\Aק��3��N���.�w�3:�ȵ���;l�0�`�n�p�9�@W1r�\>��C����4�jc�Ã�?F��9yZ���ZD����K���Q���,"،L��K/�f�o���p
��κ��Y�jI,�m�?���2�܊�ۆag��va�LM�⠃�v;O�W�m��Z�^���`�;]��ɚ� �ϕB��~l�rܵ�5�\?ǆ'�9te6QyKz��,�D�H��R�a�NE"G����d/�;dT�
У.��[u#>�ٛ	�R�=�)��������r��7�x���λ��E2���'�BF*��؍���8J�_�V�!W-�rQݑ<��q���Y��c��Y�މ�e���O>��ʙu\M�o8RH���'m�Q�����ҷ����y�
C+CF��Q:7�m����<xBF������4�0�Mǜ�X�p|��Y�ӂ�L�>��u0�7JkmR���e�˅�&^"��-�*��`Y�f�jS`�Ž�{��䴴 Sv��BL�>*
0F�L�j�
�+W#ב�|�3�~�]�,����se�]G���U�|ɑ��3�ic7�G;rA�I�dJ]�IM����Z�Ѓ�ǥ��mx-�n�(�<\��WX��R�wtdp��� 5/�l��:����s.�Y�%}�k���U�'����r��N��4e��ͮ�R��WE	c� 4��N�?vBߥ���:����4��`t�ۄ^$_ZB��4blj��y��봄Y5U�Nx:�����4��f]I<�&+X���2�t�<�*��lQ�[H�Q ��#�asO�0�0�����0��D��BO���#�1+)H�w�P��lНx?z��5���	
��}*l��������ZDƃĉ�b7�<�~��~~Ҟ�f0½�ِ���
�KhC��8�ty2K)�_��s��Ы��@�Uт�
�yzh��w�'�*��i�wM���x�63β����T|ݝ- gٞ��/=�z��=,˃B��(�Z��ӗ5t�X��UΖ	�wG�8l$��6Y"S%�Oa�D��_�ws'�L�( #������,��b��@���Vī�_;�z�*�[�Jddjcj�!+��]���D	���ƒ����?�ÂG*���E����n`�RѰ��3�n�,�����JJ�.�Og�&�� �d����J@)_xp�2L�Z&l�>E��@@�d���=e���U��`Zy��pN/=t���<<�a���!ض������4���ش��B��y���.���^,��V� �l�2��-1A��C�����(n�xV��V�j��!��2�t�u֫T%��J/t����j$,���:"�z�p��$mv��6_��r�=���GL!P��媓{���)c�3d|�)�ZD`�bR��8*8�1��t0i��3w*��m��^��2�����+�C�"N`��"����)4hC��Z��@�ߐ<���y �F���{@�Ӄ@g�Y7����%�wH�a�+��r7L�1$O��_=�G��>�C��T5����՘�Y��w�Y���/�]��=��hj��j3��X<z�ϳ/���;!\b�&�5�MS�߭�>���?��h]��u=���rr�z�fώ�/#���B��U.TMڼ:������OsF��߼XY�)���^HOC{g�����8n�Ҙ��՝$��< ~:�������I]E�m��`��v� p/+��u��l3��%��	�����y�"n�ԎȌDt������t�mx�&��'�xq4�H���/�7�*�%]ݫ �d�>�����V8�U����N0AR�Q �M��G�T��1���h�r}m�飥m��`G��jL ��g�]�]�*�ś� J8��aEe��t�eq�IDo�s{�Qk}<�����u�XҀ�,��.C(����=�q]��1=��	��gDXc��k�f�e�Q�Y*�.:�����������?��
�R��
�t]u�o��7`U�<!XP8�~�ЉB�g>0��:d#�~�'d��E!���c�`�P�/J&>��I�%�P�(����s �:�Yo����r6G
��kZ��GQǲ5���̤�R���%9��������8[f5+\��ʗ4�hf2X��}���g�y#�Vq��T���p�<ߟG����g�$�!"�����M|`�5�����Զ�/�E���qJ�El��]\�9Δ�\��Nx�zZ�/���f>�aӷ��$σ0�̻�n�	�5� ��� Se���cZ��:c�S,ބ�T��1�K��P�����:����ؒ�O�җW9i��Nw�;�	BY��̣f�%oe���x�?����@�W<|cM�����\����fHrPK��}=��yk��{�h���=��k~���/P7f�cyΒ����X�ŧW(�#\�=�ӧ�a(���m�/��g��nHP�F%K��d4�v���:�-ć�J���|����פN��DG����Y�@�,Vz�����U*�׏/`maQ}�9��Q�vn`��ѯ��{�K�����yT�a��7e��+Tx[hI�i�"�Ν8^��D"h��H$�iY�5�T�8PMYI�I���#�C�RE[�.:�����m���p�"�hD-2����>�gT�TL%;�&���Gs����D�0&uER`��]R�!'� �������L�/�9�������"����12�.����Rh2�w:��w�M?2A�[���m9N���o�K��f�<mp��mǛ�^h�����^�6��	 �P4(p����<ܕ�8��mp�6�]�j�ɲ+O��N���Ղ����z*��0!^�1�p%�zg����Pp8BY,���l����"�%_��94T^��H{��w��V��c��y|����h�;��4�&�偖}q����]�� �Ȣ�@��kʒ������d3�M�B�sf�(�"�)y"̚PW�
�Xx�l"NRd����6>��j�ײ|f�G�NO�q��h��dV=��m�5�~���`*?���/���r*�N�Mq��\�׷��}_l�U�BUtt�V����B&-�Ȟ� �,L�?J��G�p�����N?q��#�8ݪ�$^�"	��G4o��m"�/�fo^'4 U��,���utϯ>7��c蛙�<��6{�	���M#h�
�����!���U.Y�G�4�녾�oU� ma����E�ov�^��ܹ��OaD�\�uvr�)���D˨1�73M$n����d�*��ϴ��th"�/nk�\�VG�����)gzoݴ�A��v����h���1�ئ�<����/_a+eo{ 8��j����ӎ�T�jV��L���+�Q��;�D��):R̹8 ��'|K2�|��C@,4p����!���>�������qikD1�7~�����3����>�w3R(���/��u�mNn۶�^+F��~��<e۔��k��G�c�ݙ���b�6<*���$@��Zx�V��_	 h��
}�c�2�ɵ��w������G�~���Q��3E����O���*���~�unr��ߌ��S�(���;x���m�b����9�ԪP6]������}��$��䙜��\Z>b�H\��Ee��tH=�c����¾;�)}�ST��8\�k��~���h�ݍ�I�ң���D{<-�7��"�����ѹ�05��N�SŁ4Ა���mvM�{2�y)�!�([��8���=
��?/����Tl�;���g�Nv"Pݿ4X�h�a��X�:��Z�aS�C�� �j�q���)�.=a
�MM�����V���ed���B��kQ;!�T�[n�PR��q�SLv5>#����7��I��U�bC3%fm+�`�  �9��F��Ɓ5/ˈ��%���o�(ؓ�+M��>-����Hk�� �`WS��뙠D�
���>
�(%Wf���!X�V�c�J���~� �U�`�M�Ѩr.k�k��w�YRYw3í�Z?�[���#��+A
~���U�6��΍�����VB�dd�t����	�R�#�5��l��
����?��|P�ق�!����ߴ�s��Yz��G�=V�~qJYc\g��|���ݐ�<�ѹ��_���⎣�
�@$LĄy8U�kd��Q�����,.2�d�xH?���A��Q�?�bu}4.ؤ�������︎*�^������6�*���_߁�3�cG�IB�>���ѐ�Qng�
��o��ĕ��&`e����q@f���5<���^���t(�^�8�w�o*7���)��UI���3[)��N����)�y�,6�bREN�����	p�v�Wv�qF��rU�u������D(��I둔�*�.0��#q'� �h|s�׷��O�6��W5��(�R��G�f!�>���Ձ��B���Z�J�?�
B.m3��PM�v]>�V�7M}J�opi��:e=Ce�5�Ļ�Hg[�O�PSC����o/=��M=Wiwy��ÖC�*��G�v��E���#�A��+#��Q�����񱃉+�)�)�3(���� ����艩���o:�����
5�f�V/��U����3�:�3��~�<�lwi�ꚾu��R�s�G�*�.dwP���/d��ĩ�4{)���B��=ջ����wi
z���|Қhg���A��ʚI��gv7�v���7�K�7���Oj����8�r `����6�uc�~�%&l
`��2�p�����=|d@���e���.s��� �M�=�<2�1:Ѱ;����QƔB%7%kaN��!A��Âi�q�z�E ��;��BL���i���yCQQuh��z�E��9���L��6]`��?|��!�&�Y�c3ّx�t��T>��xK�5 ��h��^ٲy-?0#!�]]֬ZGͭ�R�7l��buE��J��Q�{N��SqN+���Y�^�Y���qdhY�l�Br��L�&�Tu�4��T+?�=� ���4�#�|si��9ӜΫ���
��>$�ҧ����	Ā`O7�h-�������í� R���6��'S�.���.?,9�Q�7��[��#��6Ьɰ�:J��!���j�g�n���� ��.๾1�DgJ��4q�^�O�Q ��zB]�ط&K4�>,����d{�,��yQ�5�(�ʕ�8�`3uT]��.�41�����$b�~�fJ�8���������3;<��I�av��׳��i��7�����V�L#����JQ�[Pͳ&���J�v� Y�L�-�����E瓭�|����Oy
��^U1�Ǭ�3x*൐���0����wߎN�PG��:��Vg�t��*��P�h�0�Ծ�u�71SɕP�^��}�X�����Tz�__�Gt���do6�Q�Ƀ�u�Zن�J?��|q�Y}���O��qj�kڍ�.���Y�0���S��Ƿ�`�!Pt���O��ye�C�C���z�������R�`�tl�w!�p��	���.X���(�-PTd
��q�aU���,�����ذt��涳o�i���D��U麿.�*�{�p�Y�%��L's�XFCw0����`�h���<��ف5�U��^�x�@��գso��L�no�m���HN�Ě��`T'��/n�QE�T����A��WeO2u,2�'N�J�"���N'��R�����j�]��V�� �ٶ�P�(����[���Bvh
�.����/'fH��9)�E�=8��=a�v�M���[p��cm�XlG7��l��$�kC�^g-ь��\:&�&л�����(�i)VMw�H�Y�t����XcO���F�T50�]��k�öf�X��*6eg0YQo�����]8�̚Q?��[�[~D[:�1��L��Q8փ���smC�.�sE�/�TS�����\�J���t�BXf|lMf�}C]��mgV�n�ȡ�H����� 0g\�֝t��*w]t1��٨�u=}{��|�x��K4��,����^�+:�����������b1����b鷆*�����Ѣ�E�N�!CE���Q���oIDb��ħt��~��)KQ����-��m�S�q ���'�Ծ�ogoa4!G1s����s���U?��T�����%aSb��q�Y���Xk#	O�)�J(�A�EB��yu�"����*��4�9r9��·	P���<9g¥Y�(b�j�?|���
�ŉ�Y���v��>�^��V=\A((���L�z�#$�8�;O��m����E~����Z\	���7�R�ZJg��h��#X&����۫�:����L	��r��vD��lɻ�g��Yz�}��u���v�]
�Qrf�����8, 4�b���4�֭���w��Y�p�],�o�k7��yM:vGx�"�B�B)/�^�k5>���4�&�Gc�+Zy�!!�����ℶ���G�U�V1�QC��%I��Y]'������omi�hޭ%�k�����+c��A
�	��0>�7������(��i��rlA!�X���C��r���|�ާ���L�?#Xe`�����	�5n���8'YA<k4�Z�m�w��}E���S��C�05��fXG����؎O�3��0%b��Є��������QȸH3F�T�};K���A[^�����C��qD"��-���\d�W�!�,�<D�K`v��_RE4pSy\�xߠ���4�:�l�-���v���S2D>��G$G<T�M���������y���@��6q��k�8�ǆ@x���	Q���}l.��r7qC�1��2���:F�#�iD�zeח��=����͆]U��:>��<���>�j/�7�}��2�h؃��X�z4oX2�L.,��ƹ},�ڦm|�F�Ο�.�5V8���۷�ܔ6{�&�������˄jz���+n��1�W�7QBz'}�V�~8D�o#<�!z�4\��2����=+ƕ_e�j�������i*��d�)���A"dJ�ou�E>_�O�!o>_k���5���U�5�#|yGw[��F�Z(��i�����s�؝�(�<[p��Zz��5$_"fo|���h	�>�������N0�Í�[ ���f�}�!�-�V�S�셕���HJ� `cx����fm�C���0�ɇ ���)Me/�y�@�V�ᣮ�H�������t�a�����|�r����2�N��4����q�IY� ��zB�TƠ��(��5��wp$I1��pU��2m�W�P@�U��L� Φz��_��s�ǻ���T�a.���]ϘC@zT���|�f^��3�%y���㟧3�����11�=��W�8t��Tզ ٢ιBd��_�nS�6Ǉ.m�-&<-��G�	�P�[h���%O3{>�84Y���U�}��@p��H���ŵ3Ė�x�w俪Vd׵����j�v�U��ż�Rg���K:�>�׳��8�ȑ�9����n�=�UX�O���@�_B_-��|��2і�*��U4�p��v���aJj�:E��E��0k����ۂ��NM����L��<� E�� ���ĺՋ�*
c>3y��/�"X�d2����gaIqEUF(-͟����a��*��F��[Λ��\�D�Ѕ�{�~[�
Xi��"q��^��r��|@�fSi,�x����D� �l�\U�c�i  ?�qd��ޞ���?�I�s ~�8�"h�s�&'{�d��Q0��f�]x�	�ƛ��^W� ��
т.���,���~������ͼ<� ��Ϭ�᩻� ����F�LP�?j��V���m�wkk�*�6}ƙD� +�JF�_X�"�����v�����s�%U[�z�u����*����k�p|(D�͝6}L����XJ� iї��i#�Zq�ì�=�ƿ��@n�6�}cM~����ϛ�S��h阥� z��b̩�"�Z-n��x��6�&:�]
Հ$��_)h���Ǿ���;#��� ��ܰ�� Z=�	>�:��Eg�-�Z�ru%ܮ,���~2YA����}��B5�0@M���`��W�(kzg�L6p(R�5��`��~ZZ�}�ۘ��`P�ڐ�;R�"�o2�x�9ˣ�E��i�`��nwB�
���ψ��<*vo.�[���+ �bE�'
�
��.���\�4��o�5��0��ߓ����]��xᢔ�(�4�FB�4�`W\3J��KXn=��(
#�/'�+�09I'�s���� �ْ�!��f�������O���lW�~��/?e|ϸ�Ӆ�A�K�n��������"���!8j�����T�*��b�H&�
��bU�/��/'��h������ڹ��<1���k��&�����&z�c6+��B���$�*��K���<g"$��8����z����BD��^���p�#��CyϏ��;�������z�n��g&�qP�esaC����Ή%~d@�6#��C6Ҳ ô<UMo�_���ى���ҷ0Ϋw��v)�,)���h�|�ԓ�	N��a�1�2�����ttjwb�n�D�p孎��y������O��95fb�O�̼��fu�Q�� Vs�C��ה����4<hzþj�>���'�6/�!�s�AP-�Z�^#�&��1I]`��ѵ�����J���K�Y��ɓ1ۆQ4�9х���Q����,�r���y�B�>҈���.�A�4`�H�ס��F�i�n����׏����m�>�Mv5�3B3��D�ه����D�!�Om���H�����Jl-·�;i.��~.��~��M�= \DH\7�:��Qݳ&���uU=�ҤN�G+���@r�/��9Q�$$d���؛ZH-[6��#����a����j��b�7f�Ol&�0��ay!{�������=�@�f�n��lLg�|B��8�%�B�+C�.�����_!!Ӻ�.91�1T�$u����F�[�
�����2�$��I_NG7s�\��7'�P���eg�ł��U��3>w�^��	�&���D�H��ad_��&�[�*����/U cnb(C.��t���}v#����G̈́i��
~�?/��C����x���)��̱��%���x�|9���H�	hE�����a�ܩ÷1�ݤ��(w�Ӛ�7��t�bI�3�������)��L$/�"l�M�Ł�X��{������|q�wK����5�þ��.�M��)��>��RKsTU�n�d��w���HN�D'�_0r��������84���>��&h#s�PFg��;|ҽ-WZ.��Uk�Ĺ*�! �O�~���Lõ����Ͳ�1]$��;�a0�G�p������y��Y/k���㈙Kj��ex2ÔP�+IQm�"���+i�����Zծ���F�O�9�fPe"?}��?���N�HV�%f���ȤT\�k��rY�͖6�`��l���ec�bB^P�����w��e-x♦����_�!��!
4�O>�*NKN6ml�z�;��Lx;$��\���`�W�((� TA��֮������]���Uٴ�ǹ�
�*D�O�=P�je�E�� 	��;�2Ė�c��2;�W�=�k~�D��U%�a�U�^_����T�������F`j�!7]��]*bU�=��&�G���2��B�����q�x%���M���3��H�E�t�\��(c�6UոU�8�T=�=�֦&"��
;.�,��40.r^��v��ڔ���G-SfCܞ&����?���y{�9��,�����Kډ�H�KBSݰ�2�����.�%>YOއV�F�2o'���}���+n1Y�B�[�즩jh���;�j��'�J��\�`�!�������-�a��9᝞Ñ�����Q޲�eu5?��������%#�-hŏ��Zk�.`�+��
n�\����V�!��-4+&U����H�n��tep�� ������՟2uW��lY1���F�2�$�/�e�b�Q�����ǰ0a\��M�0�"h?1Y2�pp�ƍIo1$�ĽO�-�B`��[��KO�XI*;�c�?=�}4w���ܕn��V5r�"���E&u�!G�^����Kḓ�T'/�L�w���t�g\�V1��:<���C�i��Z���FQ%��Tca�] [��̏7AD#.�rP��a�v��R���#��9�'�q���w����)6[�P��Kܯ-�}!�>z����iN�p����0�k^�P?���>���Mn0��\�i
���w�Q���[J��
��A����E���A��jq1���Vj�_�E���Z�X���7-���md�kk���>4��������L�-�.��L�~��]�C@�)!�%']O7��#'�~m�O��8HF����XU���W�U��$�c��rB�Ro��D};Ԝ܄�<��<Q�����H��{+Z���֢z�~�巄2p��eX��V����O܇u�#��(+�:+���0Y��I��Ci5�!ͅq	U��|�|j�_ǅR8%��Ӑ�[9Vלg�Bht��0���D�z�U)�o�~�z��-}��os�A�w�e1��7H����qjz���(-�F�e�8oVK[���v9����U�B��vi'�5���@8�,���cG�N_
|�F�̴GJ�:�	'	
|{Z�L�e���]��ȼE|i�!CWwQ�E�
�khu�l�=o�;(�y(J���bN�s�2fޛ��|W؁����ݧR��K��OL��=d��/q���>J�^�Y&@�#I�Q7҇��f��.�Z�-��F�4ƼҒH�/�#�`�-+��5�f�X����������88.n�M0C'Xb�v6��cl�~�t�ei�^�[���lx�ژ�& .J�R2ۢ|�
$��A�2�#�/�b���7'�!X�&�y�&��R����w`�ѓ��҉�U�[� y)4�8a�n��Y�E��ܜ�r�9!��_�c]�
L��քV���:q�	�]@��O��`�qP�Sy�?������֗���C-x?��A�
T���
�/�dVt�@��MDJOgy յΠ��W��o��Z�&N��VR��`�y)��˲�.v,�h�)�0�?]��XN�i�<ȨG����2Qj� ݍ��c������8��%Q�����u��p8�M�����QK���y$�*A���Y^��Y_���̗��o�wx�1=aM@�C���S9�`�'�5��*��S��؆e�|��G��p�Q#;� 5�՞lw�-�g#02ՖX�\����,�ӊ��N~ N��γ�z0 ���|��[�ߝ������RS����F�OO�)$����-p%	�0"A��Q��͸A鏛*:�V[�)oA���|Ȍ�B)u��M0�t�9\a����`P^Q�?������kt|��+`3k�F��\@Nb_���ڶb.l<�fť���~�lt��d<���]τ���I��K��x�OZ�e.#���ѧ���V�F(�rC���Q��t"N���Mp�����v�p0g��\`�)3ћ}[؎uv.��<��-������=~*���<O_P�j���A=3�t�0��vq`�?�FL�>OmW!A>��ҽjB�=h�~
�v7y�Wq�J�+�) ���g�-���Zܫ٘m"p�:�N������ˆ�z��GN�[�TXjݘ�P�*	�)j_��i�����!����(X�{ӄ^�\�7��h_��5� 鹘��1ݭY��,�nن!m6�6z�`eO�����<ݾK�:"{�L��Q��zj%jB:8mUm i썌�Ͱ��4�馂�� �(���a�/�Ξ�Wjq�?=���y�%bv%�p%�C��T�Hk�e�F��exo����n��
WDi�$!��n��\�����C��!�3�]�T�8~g���%��}c�I��99�R�y���_ &zt��}�n?�C�C�����d]����xjF���]�X}�w�KX�pɚ.�Z���n���D���9��8�i��s����Ck�����L�V[���_����My?ۡ! ���t.�����Ǿ� ��]�O=X

}xkpC6M���M84�M�&��z���>RO��>�䒳�~c�K��JP�7!�����@^p�o��|O�u�28�����,��ߪ����[TrYʡ�8��,A��"G�.Z����֘��pCU�����O �嵙I�"Ȃ�O�SQ����������ݮ�ڮ��"u�(mZ똃wk5�����#o�^���%�%�/R�n�)MW�����6��[ r�@����ݐ�e�����w�o��H�A�lڠ�����m��s.{�V��'�����g5"���Qظ};�3-ҋ�rd�88�l&����� ��٣/���l�'w�y� �dy"tj�T-?񓡐�N&�V���2��}U�g
$��Ү�-4�C˥�s�v�C�:�׿Gm3�y;�<pz+��n�w#,�s��(̇�%A��q##�(��u56KF�!vj9�%��pRt�?778_��kϺ�Bb�!�]�R;���b{ ��$�y��	�.E��D=m��)��)e2�]�
o���}-yd���O���/,0�zj���SZTB��C���Dd~m�!{"����@���� �M��9Q�M�@�&Wi(�����Z�'�]0 �!���������T�sRx���̤�s���#ʵ,(
9p!�4�ZTT�^����Uc(�ؿ��qo�l{�C��-���7�,��b�, ���a��B��R8X�z��[��ݙ׀&V���|���`+��8�a �.}����Y#�ŔuTHb�:Is� ����h.��?��}���~��)-�#�`!���d`�1ƹf�9y�K%ɗ�L�- އޱ�-5wƴi�����Wr)�����nus
��	۽����P��T���"���ښ�yj��_$M\!��b�ɡ�qUHl��D�>�5�&d�)!�6T�)���V<7i؆b�3��>�Xˢ1Cz���Ѳ�\�5��������"���یa|�C­f��{��H�O�ޏm�=t�F���)���hӘP�d�uo�"L7��>8�f��@=i��!ψ��tq�8�~��:��j(���MO�w���!s��X��5����J.0�U�����M'�m����6~W`��Y�l�/��1˨���18gn�J���t��|}��D�:��$�g�clg؆�1&kS�a�h�<����iQ�s��Ta�-o��>jnx�q�{�Ș6���K ����u U Av�4�����*�AS����Y*��>��/����drG��qTy�j�__bg%�}x#N&�������*�s�]�0�V�X�-#r1�1ٽ?�/>.�8�HCnٸ��9ɋ;��	���
Z�|$��,�y�m�S�䩄��"��4Wf�S�4`��G.dӿT��TNj]�1���cڬn����xָ��腂�1uU����^%�ٶ�n�ay� �y���G�Mb��kV���H�V?�_��c�2t(���HZ�|�f?���c�6���Q�|�W�59����-�o�Sx��=8��;�%����]׿�<B;�.`��/�l����	�7Ih��톁��~�S��E鄗�?��i�-�e���8�V�,����hH&u�}n��[�.�k���z�pn�̼85*R���S��ֺ҆F1�BR���t��%P�Jd.�v0����+<(HP� ֤(R�CA�B���y���L���a҇��nm�
�1"�������a@��%�S��=na���h�R�Br\4�3_κ�6O/:��iA����I��t*�:�qj�\�����g�fn����@.��N�"�*�����,�v$g����f�(q$�I�����G�����c��߭��Ϝ<�5�Ŀ
�]ɪ��[�&X=a�j(ZA'�me���ڰ�$�!|w�EAA��_`w�o��y*���Y�{�dY��K��q4�Ke|������\�u�Q(���EIaJ�����iȇz�x�����J��%�.�J3�J7i�F��*r$�	�&��O^V�l���)�h�R@��ȡ��Q<����\��L��W��t��n��d
Ñ>�
�ۡ�!�t���h���x ��� �	Yڄ�������H�����+���,2%� 2��/Xؗ~���E�b�LFlh�ҽ�D2Ͳ��.q:P�_�G�'�r/�<!��!T�B�!��6�ɷQ���5L-L�{�����)�KT7c� \e�^<��N�7Bd@�*��M_4����t�e$�H��|�3�$@�n��CCb2q��3zO�3�����W�cr�;EH������"�d���:M�Z�/�we�L]ޔ�A�n�$\����k������p*`��dK�Ȁ6��|���	5Ps��M�������9�U�
����ei��J�M���9o=�����Bᕀ���E���31���|8x���/y��)ÈuS�'�U)�ک�^�q/1��U�����& ����*�4J [N00� Z��Y���5-=�_���>�+"��sO���h��ZOܵ���\S���D�k���f�k�z��Ab/x��J=`������cL;T���=��2���ۑk2�FelH�f*����rv��p����g=/R���/q �VGd��N�����C�!*�y�x�"1K�H�Rz�TL�����@��oÝP���4R�'Ғ�뵂8=,�X�p־��i�1�;��:�c�s�k��I��a�K���{v㐙M�< c��Os��&�D����?d���o�h4ܧ}Ms� ��z.�c�[���)'~� :a ��b_�� �;�= �ajbj���*�	`�e�:kH�Ê�I'���/Q�A�<�*U'E����[w7��೙��s�@_g�X�+#P���Z���|�$�S�\V�[�����Q�����Y��tƔ��%6RɣE�4�����|8��&n\X�se��[ô4�N��R�Mq�z������plO%�z���-4ȟ�M�
���ˎ���հ
`�G�0��K�1���)/Gԇ��L���
�'tb���e��f�:���zH��FL�<#Ǚ;�������H[/�y{��tcH@ފ��4/�iM��	��'�������
װ��7�ˆR
��?�0�{�<�t[닏U�m�7H�v�/�:t���Ӧ�Sܕ[��ǌ禺fޖ!8q�?�C��T��q�����15B�.6�wj!���6��f`��褣��o,�u&dFe�ő0Q���0^y^yN��}���kW�}.��M�V	��I68��}qo�(�s~�2ø�Ue[�<�s�+hSv�f�jCz* ��Y�� >�P����ｮ�L������M���~Ԗm$��=-�٨mjG����q�i�ǗwII��MS̭Q�6v�r���&�$�,)T4&������nD����}�c�X�Z��
�L���@�8��<��GP����-;. �Y���������x	xo�P�7�6�ھ��)���!�֙GH;��\�^�9�-tTB�/� ��(LQ��J6�-��ې��n�_]8� w��1��k.\�#�s��E�Mz����N'[�
:����FsP�+>��~'���p ��!��Lr�L�M� OW����4L[�x{mp��%SGZ�1��un=dp�>����?Y�f{,�x���`��=�n����+�>���lH
�%���P�u�&�������E '$�;%�):vu�������/o���!�)����b.[$�}8p�^��R���$��X~�l9,ཉT'f� ���g��2֡a���-߷&�m���0��Yg`⑗Ӯj�Z�p�1f��Rt�#�%g�βc��&SBvLF{���A,��:Gn�mq�K�'7K��=�F|��YdB:�?Yj��~�wҼcyE�*�&��j,�(�����B'����Dw$i�X���X�H
�7g_xT��L�w��&L1���^j�!����`)�k(��`�F�g �4�O�n���W��1Ez�M����O����ߘ�Am�7��q��Ks����,���$ʲr�]�1�V=�L��D~"��	��F������t�����A�*���4�52�k��j��x�_�F^��E|2�����G�01=������ou@e (�a�_+To��?؅���_8GIx&�����
�,��0���C�V�����X�Lr�Y�1!p�"|5��	
/�c��?�b����b�F�2��t�����!��7uՔ�&ԭ�Y�ţ͹b'"bG�L�"�si��PٕX�S䪉����A*�)O)Q�L�Z���E�~8J�N/H�M2P8-�L��~i˝�ޫ�G�1�����q�x�m��h哿k�
�����B��g$vt���D���)�Q�{�,�Q恑�Ź4Yȵ�������Qu���t��Pl8p�NEDuV^ɲ�
��PC�^� ��_<"|`�U_c��hO��u-7�C�$�'4P���qj�/������	d�j����ߣ_h$��v������q V��4�қ�&�C������q���W���D��!Y�LNh#&dʟ�3�y=$�k��m�n�>�!{}��߃���`+�����)�9>R�+)Q�4h|�U����k<E���#����xO�E�`*[S5w��M�"N���]�8�W�`O;F��2: �NB9���)��﴿�I�H�b��kMZ�����<̴�B	)�[
��ea�&���'��g����Y��2��7�h���ط3 �1��G'`a��C!�;��|��������*�'���8�<�t*@���.��r�Wh���*>z-�F�]&L*Z0 X���M:�0MKU���Y#�� ~@f�#��|י� �&7V1�c���g�e�$Ɵ���Y�ӛgH~r8�X��F�,F���^�x�%�߽�Ɵ�PX����u7B$\�ŀ��H;3�3J������x$A�1(����(�r�H48�șz����6��(^%R��֙6��m��#��^OZf��ɡM؊E/������P�t��]S�U1w���5����B��`�a=vۙb�4��$�F�2l�"on�v[���b��2jϩ��Yؖj���c�*�t��D"c-C4L+�RO����ڒ8}{���+����]*O����66+R1�r	���	�f킇�l�`vǁ�m�<���YH�I���"r���x�x���F������{6��z�
�ݳ���<���^��1r��|��B�{���u�x�����2jh�ph��	���{@�wa����+W2���}ge��B5K>=�8����$;�Zdq_�4�Ƙp�1�ZSm�KzLZqjY	�hI���xj;V�|�m�ӀbA�@K�Z	0?��_��鞐I[l9�X �U�٘�[h *�h7�W7�-M(�J�?pL�A��0J9zMA��:�[ܜ|.KF�a�QQ9�I&-H��;˧�k�n}0M6��Q����QO�H?�8���^Mz�@�[P������S�,��VY��տ�����^�	��U0ρ�����?�M��J��~E�g{���?�]�zF�*K5F��y
���$�~g��e*#��y3�!3����pU7���aa��l0Qƻ��&���p� �۟�S�|)��im��j��zϓ.�4x��Z��!�P��z�Q^�u�;�E#�����|G� W3a�@���o�<���Z���A�M�О����q�KU6����v�=�z���va0+NWzCb�	;C��Rc̦@U~-�4
5��f��o��t��Yi��*����	�!	�<�ד�\
����;X*|�hI"�{�a��n�z=v@gYL�&�XS��1�� Ny�;-�����f�����3u>=��4͞f��?wɷ��M�����A:��.�\��gW[El��z��d����K�����S&El��\29�|����jڶ��!7��@G��r�F*�Q��c��O��+��p�o��(fd�)�q���A��O�L� K���!��Y
��C�)g�!��zU7}�sD�b(�/�԰wg�Ϯh\�͹������q����!�z!TὈ���j.ɭ��Q|g1K�{*���yF2ҵWU V���j*#̜9d�g�0|nnǅ���f|����}��-�c�T���"��v��qz[
�[2��M"w�4e���7�}r�	����HϢ	n�+����9�Cr�%UH���.�E��q�ă��s�,O�ak
�.�҅�ɀll����l?��h��r2M7Ds*~�(X�H�M��{;����E�"���h�$������mkabp�EK�G��!U�P��ߧ;�#���V�t�=�V�~
޾� <>J�<�QJ�bӪ����u�6���Ҍ�o�{��ܶ.�����J~j�7�T�y�m�N��MX�s����֌[7���Jd��(餈�=et�U��u;4��P/����-;�~���t�'���ă�B�j�TKT=F�q�������+�Q�"����p6\����",.��'N�\�/U�뗀"���CZw��&�7�|��R���܏8�tuQV�W���F��
�Mi���%>�d�W�P#��pA�]���ʤ,��F��uŌ4��@�ٿ[�cOW����W�������H�h��.56� �����՝��G�[r�"[x%�Ѕ�g���'�ݻg\�Tǯn���C��~�͖q�"\�dX������[�_(�H�&
�C��O�L�l���6A��c� �N�.��!=,C��Jňm����­u�f�}�����x�f7ևvg�r`]P�}DC�s	�M��A��h��U�'��=��v����3r�� Pg��	y1M^M\VUuY�oI�ǖ����,aWm�P��`�"��.�E<=W���w�(����dl̇�rL$$QG4k�۔���s�L�d
�"�/�?��N��oa��]uv�����ò��-��-���{����];m�]q���´W�vw-�<�F�()_���Դ��A�H���i�? ;���y狠 u���ҝx��9��N��JfN��Ǉ�K2Q�^X*�zu�$rp�W1jU-��ݽ�3] ��ۉ�ϖV�R�p�5tl��Dqz"�ٖ=�i��^�g��Wx:1Б될�ˊ���1\�����d�]A�E�+ۦ�u5��Q� V��V{�mżݞ3��v��Gӗ8������F[�"Q�(%���Fy_lA��n��-H��\+O{�eB�Y�-�Q�k��c��|a��U0@���E���>��P��5�GuL��c�J�R�4�M�4��(���N$c4���l�u<�H���*q
���; ��P��k��	�_��H9����{���q�;��Ĝ��aa� m/���>#�õ����\z�!n��`ssoD�L�k���a�}9��'��JU�m�1_�'s0�5�Pn�X���:����/n,��k#"$Ò2��ۘ v{xXuE�p����h�M�0���b*|�[V6����wwB~s@;W�js��傶���nu1TO�����xh���i�ݽV������d�,&[eLĻ,J���9���`�R�B��R����qSM+G��%��_'�o�
�VpW�uSF��������7��M�FkR�su���o|;W/��b��|Ć�(�m�+I.��=6-Μ�;G_��).�ck�턳N��X"��w��_��n�O�}��.���ͨ��m�I�=��Jz`0!,[���NJ�t�&�ĝd�S�I���3!Ry�3����H���L�#����l;������_ډ�#b� �O�#��=��I�r�1�v�%�t��rB&��q�U+���F��[�����4���8�11�����X
��R�����Z:�K���xb���A�v�H���Mpf�&󈒈]�rb��G��^ڈ���g}1�ʵ�R�x�B	>�����#�2߰�؄�8!������}�8&��%�h}Ç��VC�R�b�uufI��� 6S���T�H|���5mlT(A����ݱ�{B�n��D�ľ�kgg�#�S%ش��i-���qU�o��ed���43��kz�xwr]��XPAk��2u��
��^B�iI�e1�yfw�ɣt�T���t���~��73ݵ�(�TS��ew�B���J��P?n��ʈU^��Sq�8��>�);۔���pH	b�f#̵�[�d����P���E���u�Sk�-�J�����~�ί��iT�~�t��l���""���^[eV�U ���#�W��m��P;��[�*��=�K��/�@V'�N�y���OJ]떜������G���b6�b�#6'o�Y?3R�ڍϕ"�ؙY��6ր���?F���eܪ�k�$��}�F����>K�!lz �K�wň�O����$����04e�,�y�@�����������H������Fق�A7'/��������jȅ�Sф>�q��JE�@O�s���s*�b�#Ut�!������WÙ1�4��^���������9�THB��k�zcY����@���]�ـ���� �s��v��*���3͠��MBXda�&�{�C���I���R�i��5���.�t�9����2� "��|@���Ng`�Ĕd����a=Ɂ�'���1t��:l����w�ó�|]z�.*�m�D�&�Z�"�bg}R-����Ɛ�3�s�z��q �~��IRZW����&��C�b"� �Y4�P?W��_��s�g��{ޮܑ�����2g#�}��~8`gQ�H}.�eַ�t����Dn�@�δ#����Ȁ���`sF�������R;O���X㓫M"].�G(�Ş���G(�7�ӁU��pR{ZKa���n�9�;�`$�C��M�R�����)A�O�f5��@v����ܠJ�����?�{H�9E0��2�VI�K|v�� ��yn��	�� ����E>�FOT��,��ȫ-�����#����A�і����n�E���"�hPV?j���1�4��L��At���nR�Hs�����x��0v���)~R�e�KXɀ��0V�>�v���c������RG�E�H�޲S@S��sa����ca���4�Ѩ���a�@uY��AEU<��O��H����_����t�Z��n�s۾��IOT��	�6;���ö�)���:�����~�����U�VB��ǜ��3L������QA�H[:\{:ٚ����?L���"�+�M���M0�����~i
���M�x#�[/t~Eո��[�8%�YkUO���ahy(q�/
��
b	"�;�0�������2������LΦE'H�-���8��de���\�!c::-�8���Px�WB��J��B/S'�VZ��8���Z=4��h���jh!�!��	Jz�ޘr��ɲt��O:p1-���X?BH�{�w��Q&�Q�A>}DO��vi�/���&`��~�!�ʍ��c���	�Q��2�<
;k��>>��y;ye1J5��Q}�"1?�֢���y���|E�<4�����x��GԊ	�a�.�����!�+)���\�SK��b�Ωs��k����Ԕ��=8��]�ɯN���<f2���Qq�9ᥧ�d��^��<�^0�M!���'nY�J��C��^B8�ţJ&��T�8�g�͏�e�=���2���e���M��wW���+1*�З��d��/��H�t�;q��I��1$�;�[���DM
�j�WJ�8��c/�+�}��5;<dGP��(�z��M�y}�朠�i�Y3@�L?�F^�-k�${J#�(P�����s%���t/a�hXfb�=�tLM��*�'
%�z��F0m�$ʠ�y0�te��]��KzS��6�Tv�ڄPy/y�0�@&W*0��)�Zm�
%d���t(��p�����\�8 p��R��$��kt�)�Ή�7kt�4-D\�q .(�n�E�Ǫ�M���+���,e��Xex<�.�����-� Fm���$�r�0N%$?��nc��J@��	2����~���&�1��{�+����l�W�47�ڔ��׃��)ʫE�yζ�#��A\f�6kw��¨$��Ld��0G�����Ųau{̻i��4����S��٘�"�t�d�;��͟�����H8`�ӬV��r9��2swR� ��;u�;-�1��+��"�>�0$�B�|\�����$P��^�Ց� ��ǋN�@;��&H�׉e�gl �7_�yP�:F�mj-p>�\v��X��y�T!�B���D���t�]E��e)��j�X�5sȴ?��>���N��w��*�$`����^~�g3`�U�c	n�c���X�X/B8�`&Z�T��`=�G��1Bs��m��>e���	����2�Xq��ϭ�M)�#�l��?��~�Uύ�����n�HMF��3��lka��Ԕ�l,��M��$rd����L�אm]��������K�!�p=���if(01A���Kw,O�c;"9���6Ǵ �\���}`=�0���N��6�Ӻ~�O�u��~����Z7�0���4��9[ӈ�1�m��Q�?����������Ɣ1�K�Z]r�t��Ê��aUFܢ܎ВN�^�&�2��}��Jts4�6�s�*���)�o�1��]��\�[/�����=NJ5:�}�įv��cp�jp�'�;q+\ �bP��C�[~Z�`� �8cf���m8>����E������fŲǭ�Rڱ�َFs��Gd�-��)��P�O�J�T���F�)������_S}oǑ#��I!�7}�*�gMʚ����F/�c��?E�P�TO��y�W��?mi���� X�T�.숆�[��`�a܉�Y{�����k
�r}�k@8D�9JQ���tf�O��3,;��!sSmR
��ok���WѴ@#��(Ō�[ǀk�(�J�������DH���"�?uQ��q��ǵys�C�pH�����J���@V�V7f�Q�}���|t�DM�������L�9�yݎ�֨�FaL�D����N�~\쫎�?��"�23�3]m�e$s��v�$�~P�����Ie
OĈ��U��!(��(/�uJ����^��FU��ZQ�7�1&�̦	�ȝJ�g����,�	�}�ä�5`�h��ݫ�xB�IGe|U&�ޭI'��M0ቖ�BM��B�g�{�Q]�ڣ�B\E��T2OY��Œ�]ߨ	��I�c�q�O?��,����v�d�jW3<�I&iQm�?�zq���
��W�N!}9p	���!�y5�ر���懧��wM���S�C�m{!����t�%{�+�Ynn��9�2Cn�V�_�L��u�#>�t��˙O��tǧX����,�SW�ܥS�642�ޔ���TD��}M�����?#"�I�#���U��f$(d�,��aƣ/�`ʢ͵R<7��׈O7�cC&h����)��e4�Iw�N�$&Ñ�|e��zp�S�U��?3�?�U��|dIݧ�w&�볷�M~t�=�a���yF��<R0�G���<}(���F��M�I��=���K�Й�����ׂ}�8g�ȴdH��v��h�
C�(s��a���m�r�r�8�YJ�|�n'�>C�}��+*b9��"�`��xa�F�m
���h����--��JǦ$Ws	���|U�)�]�c?t�S勂z�B�d����F��~	�o�=�N���]��9�Ʉ��J����P��]��@�x�(��@������� ��D���_��qvb��.�3&"x��a@E�oM����c	h��h��3@/||�̪�2������|�J�sRZe+�8v��x�;"D�AX#u��K�2k,�S�l,+\��㞭o��f�8R�s\�>��+HC�I��e��4���4wx��׌�Xm������	��]P�Q7�f����ѳ��}���(���H˔�lۀ���I�ԫ�~��|m)F`�/��y��`c[�ӫ��E��E9n<g��֖3}d�*���!x��Ɛ���	&����Js=qC�|G��?F6�[�u����c�j��d!��_%,�ĤtaU���u�� ��3"���"� s�&�O�̕��<��[+�п����m�/�@��<�"�D��]{�{��:���W5�&�q�!܅�)!���[�sS ����3TO]����֛U�hF�0
�r�����[�[9r���%=!�<����<ӰV���m�;p���Ωe�O{��[�* ���s��b��I�(?IX�ڎ,8�Ŝ��
��8�~�C�-#�oq;*��u�Lq,���2���]��ͽ�C�D�Wf���ټN l�E%Z����-M�(V��V����l+,a�Ԝ���u�>�r?����h�D�Ыg,�T�^���r1_�'��q�B���y)�	TI�d;��i�F:��"��ڀ��� t�k�[<Ź��	L��D��&e��>��pm��kкgU�P*5��9�����mHQ�Ή;����]��ں���]7R�gY����)�\��U颽1+��8;�+�2KA�~�ڵ��q*Zf�jY� si��j;WB��r�����HF>�B9�V:�V�ܱź*���X*��f��ݒt�b_i@�%�Ԏ\D|��9c���:X;TY�>������i
�)�g	�Is�8n�kNv��Z8'k�%*g]qiKgo��+ k��MM�Z�326�;xy�*�Cwoe}��y28����m�!aV�<I�x��j-��e�U\��Y�w~�~�� �dE�.
�.�p4�����;A�W�ռ�����ke������Bk/x��I:v�ǓE�Q(,p��ƫ�=��B��p�W�'S��E�CG~�S�4����I^h��$s��9�#��g�l�S�tq�ډ��X��ml͸����ɰ��,�&t�
���M|�Y��:V��>��V���~8Ѵ�M���D'NL�?��k���D��_g�%R�2�Gc�/`�;c���M�����F��Qp=��u��b�_qA�
���u�GD�<04a�+m�C�dಙ �R����#2�?�1�~V�G�T�AQ�g���u��R�W@|�vf�7���7{��zSx6�]�.�Y�[����Uݦ�ş�J���N�/_�i���WQ�R(˚�zϫ] `�������hA�ڦ+\�Oj��ׅ�Bd�!=�����
���������zh�
c?̒ �W��2s����j窌!�Ɓ���5<.�M�9���4��'^���(M����$��!������ _^	�I�����`�\�Еtn���O��1K�=��$�ckĈ�u\����p�:=R�w)yR�w~-��|o�#r��B��5g\.8�e`�M�Յ����π��|C�3婜�uï�v�&ZgԘ���_T h�H��)�
���.}��F�(eiӗ�
^�p)=����$YI�d��Y�7�S�l���'�z�X��������[�؁�ڲ�����áSR��H[��$� �te+���;̠�_'H��X�G��hC�,X���d���8{�R�H�1z�ܴ��2xz���JV�$������p��̝-��A����i��N�eH?G�����1���?Bnӷ]�4��ɒo?ޖiw��J\�fQ���N��Xd��*�*!�F��d>�PV�#v�*�j���4�>�Y�X�+lF������5���p�=����U!:i�8��E���R�% ��� ��ڧC����Qď=�����8G���+"EQ��'�L
 2� �K�`-C7�����x�nr�U}�00�
8&�@���c=
��*���:E����,�Ay�ٿ��
 �p���4��6-�� $�}���Q7�0��
=�No���|+=,iY6 �Tp�B����ՏL�z9�t���ቖd7@����ډ�V>k�"i�m�	�q��! ��&�+�*NY:��L)��F�p,�Y���Y�31�:8��7K\��=�V��޲6�p+N��H��>o�Jԡ�tw�)i�*ZǛ�hx�IJ���K4ض@Li�H�ȋ�p@Cr��A�~UlS�Cj�7OV5��j������}���dۚ��ӗ�"��s��z�	e���ZI�Dg�����w������G�DY���fA�V�m*�Vj<���4��5Y�J`Gl���AH�t�yV�b����!i��@i��N����L�.�XW�u1c>�W��8fk��QcBr�Z5q��[�N� �цB	�l�ZfZ�Cê��a�����Kkm�F�ą���69�ϛ!�O�cC��S_�4�B��t`��S�^:�M��ь2���MD�Ggv� ���Ɔå;�b�l�!���<�����ónj���G���T1�-Ě� 6��U�Ư�E!rM���ɦ��ѷ�j.����������J~3��w����\�yF8�����To�.�`�?w�	�����i[��H)�_?U��O0��ꙙC����Dɢ�os�y�l	�Qa8�MЖ��� [8x��\�$��m���<���$��� �*
��Pl�O�L�?QC��4~�`��ό�ś$��N�i(Q�B	���8.v� 58�@��FRZ�{��A6�{��7e�E�3\��J��q�>T���l/O��l��ۆ���}��U���X-x.�W�#*��M���R�� Y�a����5~\�IDNr��������-�"Z���f�|��I���>�̶Ch�,Ψ�"���nŪ5�]�i�A���8�R�{�Ll�Ԑ��ܬI\p��0Y�{�+�0E7[-��+��V�s�b�֪gO�J���ul��g_�Vr�F�	��B���b�ֱ=Ag��q��@�GMOR�F�!�+�\_̺�ǵX,)��jܛ@��y4������6)$N�笥?�ԉ��tL�y�� �*��3J�c�E��g�s���=�6�h� he��J�7�Uګ�n��	�ga2"ٳ*�=9�������e��7����-vY������#���*�Z{��(�����K���d��ơ�"�u��hƻiՅt�oG��6k�8X9�k�t��h).#=Qep'��ͦ�Ӣ��1"zڅ�}�&�A3�I�*�s1�}���Ui��ﭽ�1H��@�J��I[�_�y��:�u�61��FM��TԸ ���Ewpkaz�z~�y��aZs�,��OcV7�%RH���`�&@�>� ���T=��nn�%E��o�\��v4��B�xa �ħJkkbT��:ד��6w�3���l��pp�u bF#���EP%㫮�����H�?�-i��[�����F��3���X��Upn[�Q���W���<��S��~11�x����S{BP��v�l2�\�!��'�#d<�`���
���C/=��PR�l�.��
Z��Y�թ�f:Z;1��w�wM��x��d���I��?��&��"�5Ef�6�@R�g�0pj���/��Fk^�@���0��G7~��!{����Q�V������x���t�8Tt��o�/}]� �<�V�0�<��`.?e��U����Ѫ't�}��;�����ʋ�w�J�\�!�F{���T�&�7Mt�����@�O����g��e^����N�-�y���z0ߤ?����w�;uVo�*�k�EkU��^��xo�'�i7�%c� ��j;�:MT��������dt��$�W=յI�ʬ,AfW���v���5IZ�CPm��:K�5��.�G<5
:� >az;K��u��CRk�����.�J�A%�ʌ2��Mf�<[K�x�ynj�cP����a&�J�]E.=����� ���wX!8�r]����gL?��Q5�4���t�h�E�kj���D=������N�j�J꧗vQ���v�|�F��5�Xʅ�c���_����Lp�Q�%z�6��uT.9D�a�@+!R����H��˿�晈�v����h˶ռk&�/]I��|d�/\�6f�ax�-�{m�j���lS�/f���`YX25�,.F�ͧ �X����������|�?gڡ�Zcv(�UuK1�'+��P	w��\�E�@gr��8-��)�^)6/xc�κ�E;�ћ{q���n(��=�hǶ��&����+kA{i�Iģ{�%q��ϽJ�p�������) ��8��g��w�[cx�A�|���XE P&<+}/�v S%��NpGsDV]���Fs��x�H���"D��s �Ɗb$�>;�c�fxҟC�/��e�g
k��<���y|
�$��dH��-�@:[�E#�������pڊ&67�
J|��!I&
���b>�z1W¦*�c�:`���B������+H��wLw�G"�F��^�!}+������=h殺�ܵ3����锕�X�x�#B+����.�%;����iz��.;E6��'Ȅ\z��f1$/�
'C��(��;�-g���I�-< �|��y/kR�U-�lԲd�����1�$��J�H­�^+[\*��ق��D�Ta����Ę?D�&S�ϼ�Z8�F��c7���T�|ܠxJ���ɵ�v��ɕ(iR?��%V��\\U�!�u#ׅ?�0�̼�>������d�{���b�+
 �6ѽ�s�7+����JP�#Q��m��"$�����#Qq�.��1 U�N��#	#�;w�n�/y�L[�E�FI�R�i;��&]z�f��6��Z�F�G̒��Z��W~G[��ki[l%�ѳ(2���-
K���JB�����axzR��[hL����4q&�Me:d�w��m� (�0oE�:�Jۈ�zw�`�h�e�\�#�G2Ah+9�7��F��pVt݅bܶ���;��vH16��O
�輸�0.��s���V������pD}�"��럠��&�M�3b���C����xj�Ė���Y����'�ƒ���cr扦��ĵ��ϘUn��:��R��A�'�����k��p@�f)�F=�:��?oN���G
U�x	vX�����?)���Bh���!wjr.,�ֽ��8�LH���H�:dm�4�Om.��Ţߖ3���D���0@��)Y����~�ޘ��7�L�� ]��q�5�OX��AT
	�f�O3t��1�ް��W%l��q)g�nEs�*G?�9��cw�Lb�!G����얤������W����(����3p��K�aYSho���*?�ց2���ި��P�3Y�"�P>�v��bJu:�{��洎�m�}a��+<l9YW��c;�l�D�j�b��n��|�

�+�-Jў��_4t�Aջ%��^���#� ��d(�ٷ��U�S�)/�*B�KEzF��]h�w̃Rwp�\CȺ��俍�����8�~��H72O��I�X�����s+�OO<�Q6�.X�����.c�J�������\Hݟ�gr���o��/��[�q�#q�5�q��1z"(b����ۨ�TIaǨ�}��ʾq���^5{8</��q�)�D��5����4 HM�?M��� 5���s����ڃ�i�T�����`��	.�v������D�S��p֪>���P �|�U�6��NV:�̜�Wl��^/V�@��jK*�Ldb�5Q��1�ьm>��ʳ�'R[{z'�[��6|O��	̭r�DK 2�t���{Q�b�gծ�t����G��޿���.����!������5W��!K���%P+���d�8-�en�FP�H�!�<��%���Z�$$��2p��9����
�?JN����m�X7�#�>��r�P��6Ip@�E�Cb�_�Ė:�;DF�AH�+��ŧPs��>��Q��<k%�2�+�
�FNA�V�'�e�ޅ��U�Paf���سO[<5�1N��:��S��c�>]<Y�V�VAl[���u^����b(b|�@���� �LZ�"�i�m����[#���`h��ơ�M�UPyD���e���;7�����Y�{�D���ߦ��9���F�=Z���K����Ez�WP�� ݘ@� �d�l�W   ���V*bt�����>�����]�L���rjfj6�(���{��c�hRˠ�d�a��`�e�HFM�Ք��ڪ�qO�m�)�B �ޛ�`M��U�R�f�y��{�*��*i�@��i:F�8��z����|��nU�Q��2z�T�		�����zb��(!Z�6���f	�UFZ ]��|�Y��2��!D|�/�m����W�Jbc���&���u��Ȍ�a2}f���(�f�򃙉뵬_�{7zZ�>�O3f�7F�v��M��� mw���&�w8Hn��B��s8��Emz�k��*��B�e���)7ۧ���ž���:�X��D"{�=#]��a�Iz�d6o�ǰy{ˠ�������S'󨫚#5q�Q�+��f�;q�%)#�M�w�s�������I9uǕ�^y��ȗ��%�q=(��v��P�X/H�|oW��⬂1�1�+��L�`�bl��8���\�֓bN!$\��]�s�MC�!&~��n���/�T#�z�(5�+��aw(�a{d���#���/��L鉆ɘ%�^�	���V\����J�7���;�*��̕�� WXi
��3=*T���P�-F��UA_�:p���ne��wXK�����l�tbsm�4ǜX�Z�����=!���+D�,/�gg��FE ���pgm_yڱ�B�G���"/K�z��`���PK����^�M��J��3��MH�.�T'm��MeF�ZL���G:�9ߓ�N	���&�T7�؁��ϗ�{�XKm���.6qν#�*�4w9;n»�>S+n�"���
�S�3���)��I�T�_�ᯚf�p�/~u�1�P���BC�wy�ꆡ#,����.�PC:6�F��+����B���C�Y:�VT�b���-^����̰g}�����w�.Mǲkd�%'�JA7���d�N*�!�t�)G����@Q���t�8r)$�z�����+RЖBbޣ�����嶆*����,�G=���z#��O�`{}�%sp����0��M�H0vx ��
���V.�՟4��O7���6�4J�wQ��eM��XC��:E4n̑d`�ci*jy�t�VX-ƈw~Ϩ�m��4/��{�14f�gS�Xf#�ܨ�d,���*���6��v]T:7Ce������2*��/�߇,� I�(`���
�4��M�����a�3U���A�wQ��Cy+7ʴችh�j:.�F�I���H�bh��-�R��Դ�H�a2��b!��U�T�(9�bK��9��u;���
��3(:ȣR�W�!Ҕg��:�naKjxTN�Y{,~���v|��Q��mȘ����^S�OF��{�^ҫ++��q �L�>r�:Q�m�t*�}&�p򉉹��%*��r�REO܃��Vu�(���D���Mr�y,4�cx�-���.�~�$s/8��4�f	���Vb�H<@����Z�5��c��x5�rh��o�Y32�˲)G'Cs��pI�[z`n+f��OFL�@��'w�~�T���C8�q�Lt��]��=�$��~�_�\+j�!^K����1bs���D&�v��j��9EM�		���0@�D'��n�qK��S�YK_���%b?����_tye�!���( ���	 b���<��X�cW�e�XQ��r����,�!7���bjT�q�8q�uc�P�8�,��hOj����-��Rp����2&��#~/LB$��;$6G	�*A�42ty�.���[Mg�}�@()r�����[�&J����;G!�徙����C������!d����@n/[���[;ۿ�Q7Ʀ�JsC.F'�ڟ�����ۘ0�,�Y��w�Ru[Ae�����QPv���C��	֝�_&צ��m�6� ��h�$�E�q�>3���;r�@�o<�o�!Jɱ�&�=�[�vRL���u�_N_ف{[��Y��SM������ђi�#������K����T0P�#N>�$,go����q�����۩n@o6K� 1s����+b���<<�n���Zkq|֥�C��s�����^T_��J\��� �P�g*Ŕn�����5��m��IB�{�8Ql����0-�{İA&�Hб�,��o]G�~TU�/�_���[bl�X�f'��Ѣ��� #ʑG\g"n�\*Ȃ�*��5!0Y��̴{�Y��̯�}��I��:�V:��<�r���XV�V`���C-1�4_W�듈����K�����ǚ��FjT�J�S�9�w:�L�i�AQ�����>+b�H8�}y74e�RD
����Wp"��[�a�_*HP���\LY��'��wI��}|`��D����A��������8��ڨ'�$�#������R�+{�G'�<䍈�v�4��4;e���3�Cz��0β(Z4�Hc�9$�w���&i���5G`��˯|\�]������?y��ߪ�m�{����i㚜�K����2	�ch|�0��=����a���VnG��e�P'���e!TQB��+����:��휧�����-p �o���Z"uEl�7ڏg�#X �iN)�'1���QA�5�h�d�p����G@~��) c���J����B);vV�K���, gɣ\��C�m�� ���Vw����Oa��<����jr�4�H!��n�����Hi��!<yK�5q�������^+AL���NU�l92|�����=? ��5  :�s��Ac���l�_�Ĵ���D�$մ�xJR��b�s��X3��2�rz���!m�5�c�ŮOm��U�iӃ��i�����J���7�0�r��x(uI����RqHI)�q��-\���ҕ�eiK�J��^V�D�%|c ����3�3)x�u���z��k���=���]%�[W��]K�&���禢g�:J�)Z�ޏ�m��ho����Vּ۔�fDÈTw!��u�cm�%$����� 78�[�b��%MgI���q.U<��X0�����#?Nr�qN5��$ǂzp)����Y}���k�
7UbQ�r��t�������|MB��5/4��TC�'b��!KШ����yǏP��ţ��l�܇k�����0��x*������:{���ޟ׻T���
O,j�[���6h
��$��N*�5G�B�g��!jR�]��"�9l�Jl[�x7���O��t��=%�c�x0xʖ��/��H��W�X��:����:��v��&/��{��v:����|�RN���]���ߠ��S d�pٟ�l��u�����$�k^��B~��9���읷�¢E%{qH�����_�ae<��]�b�J�=C�e"W�Dsb��w1BUK_��<�t��Ea��kSpŨ�����O11��{�T�&~�� (̠��!�}��>��ɚ�fT%0���;�iHZ�J'h�D���Vn�f��{k;>�>]/��vJ������nvU0���A;�~��o���Y\�>� ��p�5�H�W��dK�aZ�H<�A:�͎�qj["&���s�.�!�T1AM�����xy���F
 f�-C�KF ؖQ���@Dٲ�\�����g9��&Yb4~x ���A��ut���E�X��`[G��upR+�*�$��).|��xO�y�ڵ��l����I����
��*-��{KTq��F�q����:,s��+l*���1�'�9�'ɍ=�m���3���X=��u�M4W���]KA���ւ <�L�f��-X#+F!p��)/61]Jw��`���`�T�����F@���KG O@Υ�D-���/Q�[�QN	���Bh�n|��H��/�^���zZ7����Aѐ�7��K�t���XX��ڬ���)���H��!ѯ=�
�X�5F��Ƙ)a�͵�eM��:_��3B�� �^�f��CcWC�U��Y)�0�o�4f��@Z����H���}j6dK�����rkR���5�����;�D���u��u�a� ��خ7w�%Ɋ�}�WF=������զ2�A7jOs#�,� �H�����XY�iWU���@� ������Xn��B�#�S	<@�*}Ȣ����**n9���r��E��8{�^���+������W]Y2	Y�y-3B���� aG	pߪ�Pr�]icV+U�wn/*ruV�M�x�O����]�g�4�g�
��ɣ�f˼3b�E=a]��+�gW��h2�B��%=��pI���'짞�5�b�N��{r�jQ:����h7����Z�|�� �U�;Ouq�2������W���DwDk�������+�J	�.7�̦�%�:��A�>�B@���n�!�_~�q��ǐ�$]㍔��e�����g"��ư����f�g~?��=a<�7l��Q̰k.������0�3����8K`�P'��q��0�%,���W��J��0�4��u�y�]��m2+�Pk�@��ePfϕ℘N�rFG�&S�aW[�f G���u2��w��®t��e�t�ٙ�6�����h�L�4���1�_��Ϭ��ZYje	��}�X-���
ͻ���4
si�@�g%_��F���<>6���}�ʩǳlƑ	�P	��2k�h�LW������?�`�RL��1u�i7���u�������I��qG�ض�)U� ��V� ɝ� f�-[����;sqd6���̴j�E���Ay�X��ުFp�++��D���y��ʓ�~Tb���I�� 9p�%!��~H3ᴖ�k�J"T9Q���q�������O�u��85&�~�x�����0�8�ݑf�
�Z�ɿ"���er0��$tJ�EE�=��a�1^ ����DgJ�6���xHw�.��v�Q���.� h�l8�u�������i�0��h��Hb�O�{��%/��wr�0l��6P�� V�`���"�[�aV��J��
a���)q�FNN{u�Vc��z������Q|�DϦ&*]h����Z⼆'w�t�)��wު�}���Q'��F�lWGE�k.��/s�ګ!�#w��u�n]�.��yVk������!�1���n����:�j�l &�8;`���n���e��D^1ȸw&�8�Gm�aJ��#(}~�-����T5%�ؚ9����~�@?p�]���$�"��.�\��󰊽#k�6Iȵ�͠���-z8Қ�z�%��������B�`B�H����ڪ�i�on064���`~��XQr�����\�=t!�1Q����R��J
����L}
��5��a��2�DT�^��[�cwo��B��,��*�������.T)q�n��E?����.堷��)ad���IW����C>�+jL"{Z8a^��"E�����"����z���!l�+�Ł�;����t�*�*a?�Y*�/#�֗O*@���N&a�[z����2�$�an$�pF�
���f�,&��7p������ VVҕ�4�j/��ȫlA+~�W�ln(����{�R�
����t;ji3��,o�CB���L�����|u[du�%������N�?.�=�.���i�Y#��֓�!xu��܏�=ժ�a�*�GS�M��]ܤ ���}�y��_��L�T��T��B������������f什i�rU�#����V2��n��Z����_J�Q��Ȼ�+�k�-�A=uҖ�{�-b����F� J�v;��L�W,���h���>�ӆ�֓d��O�9�VN դxM��q� �3�$����B�ѺFB������W�K�Cxd����u��J���D[��_� 4Vȶ�!�h�.��F�V��c�F��B����	�9}�6���>��^�ZSj4\n�� �]��bs�#�8�{�b�߉��! �O�sn�D�t� %	�=�Upo|^j����"+['7a���te�����"�-p� +����qM����>��kPV���q��9 .<Ǆ�q*L�P�`�W�lQ�G�X���L�3##��l�=*K�ȭ�>��C��Jf�3���Gi^loS�L�[*Hi]V�O[);[Gg~~L1�]�/a������ԣ�r�J��R�i���9V!c�)\#Z���t~�Z�r�ƻ�#�2��<ĸP�r�'���k�����ގ�I����H&`	�Y=lcI�h,"	��-ʂD�бE�^�yɧH��&�d��'-Ϙ�Ay�eSYW�𲍲i?P���a�M{��fo�{{�������z�Q �
J%'yn6H&��	��/=��#H9-Sj�O{iݸ�x�a���]�~�g!�43U��Dd9�a�w��b���>y��gew��J�F@���m����Qx�2�xu��R�A�}�ǝ�n���>T�w��C�W�.2���N�����"�P���Nn>$׿��=����e�L�mԳ��?B�4��rlIE���j��ʦ��y*ҺQ23Ư���L6mt�$ɓ�*���ǁ�h/
i)*1w�5�D�;��B�m�>ͨm�H�|�Y)N���8lw��Dv�`2;� ����2lΖѱ�j���ұ]b�,L"�fG֠�L"�B�XW|�����{{��ְ�q�*}�������(����!�8�2	"��j����l�;����-An���#8���E�V�$'����b7�{�D��׺V�D��~o=��-�#<�c�>*����u!CApveƹM7����
wg��|��*��d��c�%�2�ő��ZQ�ظeG�����n*	6 ��z�R�,n�<�\a�dNa[�K\��oU��>�x���u��)g�2�j���P�P��&q�M Rmug��w����E^�N�w�_�c~$��y�~4#�8^�	hc��x��l�d75�U
L]��h4Rqy�f<Fl͇ˆ&If!�ܞ=���-퐚�xx���G�������z�"�Q�c�ւ��$g|N�Z�
�����	�7���+:g/<&����DU{3�'�Za@�W����8��4:��~�~o��~H��N棒���]p*3�}�kݒ<�P�H���H=]��u4%@�:4��7h֩)5���0d�؟�	�Vs��^���)���?)�/��Z7E8��>��>x\����y	Z7��*�&���p�
��������r���<1R�z��`'��Y�^������O�B�ba�v
Eti2Z���ڞN�n��
0��^�1�\������G�dVB�.��k�h��鮳Q�\SXvq�Џ!��6��ƨOʲ�]{�ec�6�4t?������e�3uV�L���{�T�[��\qً��S�-6I�-�V,a2y��)J�ύ�H�9��Z#_��~غR }���yH��Gw�a9�<˜f7�i�-f�J֎A�AU��1��v��ܛwtgV�ݏz�)������э-�����S��ۇr@�
8�S�S���9=�*��D"�8!nl�h�?dN�>!B��ra�nS��R��m�	s!h��_vcP!��J�m^-�^��-������p���>@H�����
@3�u�>�$<ʧ^��Y��0��B��-�Q M��Sj��_yQLh����Ϭ����C�#�L�4�2ѕ�|��R(O�R��="�(ȁ(�ϒi�3����3'^u^����E�P���On!nv�r���(U�B�_
��~�\���?x�_s�A/H?��BHk�/Ҙ#��ƨ��9+Yq}P0���E���3T�л�
s�>�r@��bF+�J,�K�Ka`�b�o*���s�̱鸄��d`�(��o�o5�̟,��бx������ycF�-�@fu>� Ē�� �
�>	f��͆o��\P��n��L2�r4k%G�D���R,v񄚱���n���R2���(6�ǇM9~	��YJ���:}�O���Z^f�'��$�2��!t
��U0��g]�0��Y�&Qg���J��9����G�ɼQ���&�]pv�[��d�Ȥ��r?`�?��]��l�r�Ѓt�W��h0[�=���hg��x�ف/� ��
M,��	�Ga��:�����e'��^]��I"^tf���½���<J2�5�jP�؏�(��KƖ�֐r�#�-Mb!��4!(}W��j�7��p��1�zyɷ�?�@��p��,`a�U)��4�>f�>7y%�UK��;W����.k!���NzV�'�_���AK��i�� c)φK��]2'Ƃ�Y��� yX��o¼__4�a7{���5f90|������6�_�zzӷ�Z�KB[��
�c�����2%b]���I�c֒����Ǳ2I��L�+6;��H}6�az��$'�����w��Dc��C��Xʖ�&�k���gj�ZT4�ߦ����weq/�?��IP��'^�&6oݰ��p����/�fj���#չ ���������v�q��;#�y�f�ǋ�?��>"k�ee
ļW��δ�~�bL�p^_��%hB�,�xDC�:�qƕ�4��Ia�45V>f�Q�%	����pu�2�~oS��%�6rN�c]`yG�SO����ΛP��o?Ū�^��6r���j�E�P0w�Mꯈ�a&Q%{�zi���C�λ�#[�ɫ��~�7ɏ��|�W	\�q��S���)1j�����k��nԫOh,*��û@��͘��A]$�u��YM�_� �~Dy���v1je.U6�K�9�O�L��t�l⏍č�ke�?V��  nR�dLx�wS\�yHD=L���a4��)���p �_8%�v+�[<��i�R�MԘ�ǲ�A�'��]}of?�ّ��oS�5���!��G�� �G}t1ԋ� ��M�:����ۤ:��22C~��OQyM�:�G��0J
^��an�_�{�1�Z�\��k=~����$F��w LT�yqh�"�+P�N&��]��(.viH��Q]t}�$X�0��\q��~�D�@ATS���o��{5����u��>Yg��j$�:���>��&I���4O~���'@P��<�Ć�=��(c�e7Gs�-��_���!�57]��`T�����N�S�Gmk|�?M/c}���U�����C��&��xB�݈�Y�;��ܰ}2`�D$�8��հ>�i���j�Yo|x!Z'��%� ����,�;Q��~��,�bV��bev���1�@%=_D?N7��X\�9|ǥ�I�OKUs~' �9N����0U�u�Fw&2� ��A>�Bg�D~ކ�U��s"���Tn&��	J�Y���Ss�S6j����P�4�����^���P�|5�4 0�@�Z��a�@>�+�e�Ix^P4�o�Ǫ?q��-���Z6� �v�]�qk�E%A2����P�R�c3� ��	��xʸ'[�¸�a����S�tz��8�Vb_T	�Pc6]6��9W��<���'Fi�t|�+���`e��P�?+4�N��(�g�Yq?�h��R���ܐ�\=�8â����"�����8�	�|#��(���m�5E\����D����Ƀ#��3����v4t��"̎�[F{�Va���1���Ծ�����j=q�6�s�����
/�x,�CR1C�_�_��dh��$����  u�U�:��%sAf�6Y�.:��@=E\ m(���s�U����Ț`���Z�<���y��*\�n����&nh�ܣv&iZX8��}a��G�l�q�+�����ΰ��w��ў��iX�Q��met�è�(e�IQ4s���D�:��8DAH�GC�Y�H7�>2�?_o}8m򲲦z��X��iD#�CC�Ni���0�v'H.냾h�H��������2N��!���X����%[v�b �� 05q��th8� _P�-Y���99rg� �mZe���h��d`u��W���=7��N�_J��Xvp��x��l��O�g���b-s}ޕy��~�2�D���|�������Cm��Ԝ���Z�I~����*hD{�9Y]%��t�j����?�*����������l_.8�i��� �⇹���<"���[.���a���+�i奈��?++�y�	�^Z�i��b'�VĤ,
���cN(�j;���X��A֫qlt/����iÖ��9C8w�C����zP�i;$��<�h��EKr�[,�y�A�\0�8��"��?#�T��koR�
���R��-�믡��U�"�?�A6':�&
�֍��;4�n�� ��\s�z���j�%F;��w�l_"���`�'X���$�j�y�j�����_A����8͇p�H���V�!�rev�TX�������@�l�rx�G5d��]_
0L���K)��$R�]n:�dg�9����"�>�v�
w�K����P���	̏'���)�����Y{}�Pc~���+u�}oGh���'	�]��`�*�\�VA�@�*�%�z�F�@�q�p��kAӀ����Q��mo�:�� ����0�F��֜A	��6}��{��>�Dd�� uO�Wq`��Cƫ��cˣ�ɳ����p��18�g@s.�Qd��Z2�%H>��@9	Z�m�Y85�~���Q����I�x�5_S׈��x v�����ʾ�)�.����-��/ĮL\�է��~�&�F��=��g�փ��"C�eu�0�G�wV�>�����
g�ŋz�X[��gdj��Ό�g蔴��8�w^oPV�|ڂ�Z=�P��#�"H����&��t��93�p�Ғu�Ĩ����R�������T�Yc��Bv�!����s�
edO�tZ��ogf���˟�U�c �p�
PE�Y�]}�靟�W�o�m~���^��c��=���m�__��L�Ei�`�2� ��YǄ��cFUU��W�B��I@��xI�s�6 8��,M�AYy���("��	��(pJ=�+�6��k�����e��6dJ��M���I�=��qI�n(���:ī"�散,�O��o2O�X+�C���2�:����L�=k#Y)$e�5�qT�8�Tnj}X�KAB�s[:=-�����Y��p�	J�nQF1���d-�L4j�i%��"��Y�FJU�Y@
����-G_��T�;ü��9Ӟ�~���#�u���em���]�̂�VG���Elu��K�uӠw>&�`Z���&Mݚ��r:�gL$pk��7���u7*�)��J
��?�b�B4��T}��vi㣴���8Hϑ�Ռ/�`K��C��.(?I�5���C82�訒]i:^�ݤD)\Л�����N�J�����D�C,�绐�w�x@m?�!���ogZ"~�_w�?��ej���RiY�T���5߃[�)uŎT ���4��z$3:.��<�+�����b���C18"jG'� ���s4Ω���؍�mT@�W���e�)�A�j�8��B�.b���g|_P�4��/`̍R���0���9�$G�eJ�L�G��}ՠ��z��᣿��x�БM���D)4pS�b8臫b!��C�q�b�D�n��CB�,�dR��8��#g�!�nR{��ͬ�?�)#͕MǚC�tO	�����T/���c��F�
b�(<�6��/3?��7�_��S��������<����q>����΢G�6,�	@�Qu�[PK�6\�ż����Ƽ~��T�͚_ҡ�	�V�[���KnJ�O~»h�甙��C�]C{νY�>�-�Q��Rǀo,k|��«��Yv� hLw�5;�!�����w�Ղ��3D 1Ѿ7�;��g-�#7�E,?��Ч�.wx�a;���{p�:3���ë��b^������1+�UސV0�+NA�w�8�7�㊒',��װv{�����`�i�/r��M�*�D����`�.�m°��*UN�לG%:T#v/-fwH�o��QCmq����>P ;�4BM���63uG�;�"��[�]�}1GU.h*m�B���3JnA	�������`�yz�u���ڷӊ�pO�Q�p�g�Z"ގ��y����ϬQ�Qc4��L��*�.mz��M��!�'��4��,����j���RS���7��YC&yD{��@�p�@F�L�%�k��� �ogs��,�>�����J�Z�D�h�Bi_ZC�W9�F|��̺�p�
����s���A�u���>���,�izc�8��uɂ���a���Z�l�T'_��ͨ, ;�~	��~�VE$�4��N3��q�WM��p ����z�sM4w�9�i��W?����*;�'&d:cM������h�A���tJ-����A���wb����C9έ��i�W�av�K����,@����>��,2t�#>�X	x����2�)}ue$(;M����PVp�i<<����z�����u�8�������//���A�O���"Q���=�ɦ�����6�q������'[/��0����F���<?�Eش2��as~I�Ʀo��"�(ɥ`�S��e�'y)So��`-]���9��5�{n���e��<W���^t�$�0����e��P��s����iw����c���,~�\�X?p�M�������lB�>��S˔�`�y�dCȬ�g�1F]��sE�y��j��x�;��w�'���P�4G�9�pJB$�v.?�.(Ζ�u�Q���Z�`@0cnSkg=����6�p������)��m,���i�]<�wR;g2��_��B}4��~�!�~X�aC�U�%��m��x"T�hX�WlXJ����GDVt�Nm��etz���%�c,�	7|I������ �&n:n[��C�f?��.=�#���?�� ��0>�DXI����I��%J��$�8.��B�\)���O_\�KH�{�B漧�hu�r� ��Ag�~�����'Ų$E�q�bH�'\ūH���Htd����Ev&�~���%�����c(��(>4�'���h+,W\~�U�8���v���C�i�K�U��#�\�_3��y�H�j敓"im�5j���W��S*4 �;Ħ�!=��b��rP��w� A�W�*����2Ĉ�7^��hծ�7Qm6fژ}��u�DrF��S�,}�$RM�sE}���ǔ�}	|p_у��@�H�e �"뀷~�{����?�lmԺ'}C\�H�F�{�o,��&��/� �{��}�R*�P7f���|g$G���}���G{���c��w]3�3��tx��\��:�vz����4�%:��Ez|nV%�`��VW/���d <lw�B%�N�p��#I#���S7�G���M�TVy�v�u�s��ɀ�ƛ,�����s���&�[�jHZ �)H�R�6�X�,�?���z�#�F���GZ6��ͫ�<��>�D��4�o�[V;�EH>I��R�w��K�J?I��1�E�߮��r��� h��ў��Ū�[��tU�,SeO���ͧ��+�"����Hg���L�2�˹���Ǟ?DD�8��P�+ 4qs�i�\�1.Tb�r�Z��8x�����O:���3J��	���9�Ľ�����#�q�W���s?�[2��Zs��`���w���-(G_�܇�55���� |^��l�:��}�G��f��D��O)�њ,콾![��u?R���W9��3���z�Y�F{Th+"3�BM"r]c���-�A�%u:�C(��A$��«��Z����������b����1�]'�Ao"�R���\�.ud�+�~"���t3H0�=(�4�hR�lG���1�I|P\�H9PsY؁�5!�����RRZ!W#h�`���Ė��ê�p�ld���y�О�zOc�Q��?T͎#���>o~O��J^Bi^�����'?�˼�efB5#�Z�Bjk�#R����4V-`~b�,�1��E�dl���[�#8%��e$�@az^��:�E�L>�#"�����7ҵ=�u!��xת�6�*�bXMK?W���V5_'b�	�m�#S���Z��=X�l:1�)nT��v	���inr)<z��]��+���s|{��~�X=՛����%X������c���UN��+{C�������h�?�5}�������y@I����w*��r-�b��~�0עRK�`-P�������j�1���'mJ!�U�k�4?�}��ym�o�P���H�k;u%��uO�>6Ľ��I4p�\k�k�r��La�!�%4�6�0�=	�Hf�i�Q����.�RB��;�䛅���u�CgW^���|���M��4 ���>k��Ed�N�H� Ǒ�rf�\D.&�a������I�e���ڽ��CUJ&p* �<P���D����i�E��jxR��3P������kY-��a�#|�aX$o��1
o�zS#H3��=����2�$�-��F4�ǌq��c��9�!u�x�j\v�\����\ƗRN^���p1�I��+�%�f�l�,TAp����.�ud?D-Lŀ{���kd���%�*+�筯��Ti�Z��fx��?�	��ٗ�M�������9.�Ȗ_���T�����s�{�yݏ;�S�M��
/kX bK�O2�<�ς_^�+e"�(�ٿTNO��0x��$:O ���s�q%����G����~�M���!�%�.��g�'z�JE�PΘo������&DX^� ��Ls"�5u�~�ʲ�;�I]������}[�~�DK���U�U!3��?�by"���?�`�E�Q�?�9V�9��ʶ���W�P>�V#9�DI��B��[�6�s��ۅ�e�z���<���Gp��Qԑt��M�25��џ'�9EGW�sp�Yc�ź����P���IP�[.�]�|�c��{<@t���z�M��}X�7���3ݶ ���3Iჭ��[ǎ&��&Y� �r\���]IZiIn�nR�����pO|�ܹ������x��9	XG��k�_�)_�%d~E���P�ԋ�]P�=")1Q�W�E�'�ֶ"�������buXԆح���iHm��]������+�_bq�Zo���p�Ƒh�o�+j����s��_�ƣ�=W�z�x�T^2�E��Z�D�>�V�U@	)�I�E�Li�Y��ǚ\�����v(�����9u�OP(����9��+�=܋��F�D�:���Wm��Uע�$;Qf��֚�P\�Z�uE�d�*�j9Q�F��W�d�$} y�Μ���Z�ظ��{&c<�5�Z"W��ɶ�� �<|�=�8~��:�K������)(�8Ie���Nx6���ɑ��`u@a��8>t��9"�'����JJ��a�×TC���ach��_Qc�Z�ѕ�K���k߆��/eÄ�+k��Φ�Pvv 1gf��<�s��TjHzzn��i9rx���:�g �Q:H��x*�OT,��;[���a�M�����)[ MwPw-�����X�uv��A�Ւ�t��4��E>"I����^��/?���/ IfX�xj�e>C���Z��O���o��K��ݮ!p��E��¨1���F�o��v�/�qi#M���g/�g��k3c��M5�[P�=�޲�E�;���~e3�SK���E[�ހ]���o�M�Z�h1g �$����`���� ��ik�қ�0�c��z;͟��S�km����q�n9����v��Q����B(3έ��~��� ��*���f�'�M��S{?5��E'd
(��� �={�^�0'����8,ae�\#�J���p��%Cr�F�����j�}�DC"Ap�F�厤��ρa�ó��'L������F�r�PH8))`�&̋<>�A``x�j���2�c��棰�N��:��!%��� }4�?)��ͨ*�M��1"\&��*�"���5-�>���(�����?:/
(�=�0�� �	�Z#DԺ������]S�@���\�?(��Ń�f���5I�B���7_�!Va@��|C�bR�	��D��1���鏎�X�,gT��D�i�fL�>���Gx��*���8�@�np}� 7�ݱR�G�:}��_��1�bB�<�9�h�鹶�a�5���~��͝�E8=�}cx�>qT[�db{��M]d�nټ^�Q��&�(���#��J����8�h@��ZܧY�nm|> W��H�F��q?�K�����u���]�֛M�u�'hʨYj��4�Nޔ&;�eE�q(�d�k\�ur��덁L� ˚{������RiBͧ��<�f���l�o�JT��F~"�l�TV��޼��X����OO��|Aʺ~�i��D�:q,�ؾ�ux��4�O
x�[=��n�:EM�]�K� ���KMEd���U�Ը���-����`�lV�t�
�^�qo��[�1!��S�H��տu��H��;�:�~ڏg���Zʅ-��������р�q���y�/�;��"dL�U�p,�+V(�O�`<�3��V4�B(�z؆j�|�[���
���6�퓣�r�RW]<''�����93`���(���孈���,� ��$�Ӎw� �f�_%��rJv���վ���g��r���w#��aGI\��Rq�k6�Jغ��R���E�������#�wɖ��|K��j��w��Y�d���}]��K�pQ�z�X�X9���v��9l<H83���f��-�tfœd�=��.祊��%y�G�$U����{�z��]���6���*`�t�Y�,���'F�u@��̐%��t�;�����Bd��{�n�d����|�u��;)��g�������$�, �7��'�3Դmy�]V�\	:&W�㦎	D}�{�.�ă{I.	����s��i l�:\�77s����mf>0�Jz�2��˸36Loumg�A�\�I�0��~��[��ֿ5�k&ck19���,�0��PQM�:������7�yo��蓤�`x։Gz�� �0p�Rq��*P&�L�ϓ0B<�E�Ζ�t ���Aa�߾j_O0�N �MI���~�Bo�A�gec�~~|�ЛO��Q�{���/�;��s�]�,K���|�(}�N��=�p�1�j��I��3����Lj����_�;�ߪ|q����_���U�uW�i���;J$ٱ�-&2@���O�ӣ$�C]���\���笕�3���5k�h1ɡ#��o�k����|5]Z�@H>ǧ���6Hm���4A��9����W�a3���ѷ���$S	�w�;���GWO�7����-���B3�Ϊ�ìh�-�l�籺�`*h���k�����I ����o�:ع�U�kix{��훑�n��~�e��d��s�1t�zh8��f�@�ڹz^D	dxp�D��H���'T�\��Wҡ�;kǄ�Ga6� saQa0	�f�K:8-�p�i�C0�R�0���Ɂ�+Q߇��������๦���@D�b�#��%�[#�1�iFQ�����m������m�U����l���3[�y-I� ���[�T��ߊ=׺���h�������%V�^�n9}����mXPN�U���k�����C�^6���Uc#�����˴�� �� �P���P2�N�W=V�MY^�rJ�Mfݚܜ��ȱW?�=z��R�<3���?��t�R\��z����
cn�5D�έ䶾�4���K�([j�v�!@�Z��!w�]�	:ɖW�M*w���Ս{��U��3Jm�R0c��/�����?���&�k�����G������hJB��'�D���tⰊ��2�d��V(2�Z��������­��dP��$ux�j���eA�����L���Ώ�N�
P��p&�s�OJl�w��jC|��Z��2���o�1 !%��$�m�̋.<���{��/o��^>��O]_���W�����ٛ~�Xm/��B�0)��ى�57q#L�g�zUmi���f�_�gT�;�&��T�@0��DE5&��qIh����Na�4	S��ǐd��Oh�>]9�k:�����D�4GCW�3�i�ζ�ً
"��t0����>�m<�0ac�*�UT�ub��e���2�m�4/��۔v~�k,��©t5����$����t9�މ�4{O0�����L���l� ������?,�S�yG�V6�	�zeq8����ڝѼH�Y"��MK5Q(�M��jK��2�
مǰ1E7�<��ߐ��gi��j�ĥ��U��QL�L����ԙ%(4O����!<bD�{g#�>I��=J���K�K���y���_
r�oV�pA�֠�&=�j%�8��P/�=��֎F��+� �0�vp���5+��{^=��ؓD�rnEoN��l]�3pC�Ǥ�1�X���d4�p�a����p�an�U�ғ����\��3l�5��!���EǙ���
�(������C�>r��`I��N�3=Œ�p�jK�
���A)�똅}Y��Ø�
�'���)����ү{���cʻi���S���?�;��N��jj��-�=l����3��if5j �S���Vr�	n��I�%��>ɧ���ax-) h"�E���B���kK�zuI�U�a<��#��r!	�8�bRi,���*u���L��FA>�d�;�|]t�g43�C��Bl���߁EA=����C�D[���1k��~X���P��ǜ��).��ĶГ�1Mǧ����C�>�
k�UkbR���t2�!I1Y�����˹��|ֽ�^�۫CݑI
6��/ك�Mz<�I%��=�B)�ѓҴw4Hx�(:��3@�^�}Th�;����+�]B-��v�w�k��h��vѫjQ����ԑ�}�q�p���'�p�eY����ٕ{:���O"UP�uޥ��܌$���қ�K99�1it��	^��}&�o�$��M/ҨO�C�ܠ^��)�����ab˷��H��V�=R���.��^�U�~?3j<
���7�ye2}��� �J���nf���8�2�G��	?�A8$�T��0�X��b�fؚHp�i����>�h&a��Ȑ�������)��B�X�0w��Qq�)\\��{P ��+������]8���8as��cx �*u������ݽ#���Kh�ȹ�S=�mj`��$�!��J�Z�ZN� �pw*B��F�x�L��A�=X�\ok�r/��tL89c��Q6�f	Y'�B�&�I��U�r�-���Y�	��5�`6�6}�my�gI�#u�\��Z9*��+�"���Xqo�oCD@آW9�����b� t��B��YL��P��,f.�[cKt��RTl^�4�`��]:��r��q�n��u��%'��PpV�05�]�|w}���3�x�ҍ���	��+����P(dt~c=a����q�)MtdvA$���������֓���P�X߯�k��<�N+���F��)�ͷ}+ �A��z���KN�"8�J����̣��3���:�g��8����q��T��N3ۤM�&�T�q�̅'���J��@�9���Z����|\��u~����� ^��WlY5�jO�E����1-M�E�<8���p�\V����"�S>�\��D�}v&|���"J��C��>�_�~�r����+ �� :,����\Aķck ���Q�W!T'^Τ�!�hXWN�;���ݟ�4h�����3�����"���h�U�.���u�$�xH~b������Vj��-�`e��;芶T}����3�,��5V�����t{��᝽�޿T�`t[� �|����
|��;���JpPߎY����ߎ��K��,l$o�;G�������F�5�g��'�t��k���;R�;����ȿ���h�.说(�}�kl�x���D�$>�A�cq�1S
&rҦ�pl�صl{���#o(O�6��ڣ��

k�%Xy)}V��n%���4P5���]��6+0,��)v�r���͌:� )����W��.#��cZHb��'H��_>m����Ɔh|�Δ������(�k��5nvI~�b]Z�k�cC��a��Y���e4������x��LV��gp�i��u��!��cU�̯�n&@+���?�lq��\�'���'L���6�k;�pw��~��~*��}8�HF�n�W?m�[3"$���4Fb��?ݩU���~�.��t��ǯ��ʴ�7k$	43��w�~D�s�W8�D��'�9&a�~S��Rk!KӬ`۽ڪ��I�jӕI�ݥ�Ϊ��,ʣ3�2^%�īF�?P�����&��U#�������I��uo�ꓞ��<Y��=v|�ܤ�C��E(�8���^�2OFǊWX9�
���*θ,޶7�����Y�f��OlA���4bx������@�=c����CC���C�/ct.��&��A�㪁t(t	��ȹj���ۧ'6�р�󻆋�����R�0���V
ѝ"�{�תNp�[�ϣ�g{��<�b�A��=�~���B�r�`"MB�r7H��[TJv��|���$֏q��j�AU�r���ς�@�+T�ό��z���e[���C8�R�wn�ٔ�'�������������>�XI�}��c��3�����������>+)rRs�Iۤfۚ��/���A]}��U�s�9��{��8�i�u~0u�W��r4
��W/#��FW�����������B��.ǉg�6?�p��"O�[e����`9?,��4RJ��7��	�-L52�j���c	�����~��t���b�8���/ӱ���犳B2F�a/�&@�ЪmJ)�0�l�E�l���(B�p��D�w֞ܯQ���'����Z��.�Jk#0 (Ŝ�G:L��pf��㓓،u5_�J��h����D(;�լM���ClOC��t��f�M��Dx�7�3ro���`�f�CBs�GVL�!q���t�ЂN�`�_?]CN��Iw�_x����=9{*܅�O�}@�]��셀)�*��r�a>:R����1 <� q�ΟW�b�f��������o��w��q*>��K11�j�d�1#R��D�R&�QO��1Kj)�k5���.˭[���'�x�,S�ٛ�Z��(QB#Sܲ��}`V�Þڐ^D�nw���-
���hm�v���)�ג���6��lv�f	���Ib�,��.7>�����l���@�� 6{q�$����B@��cX81���k��%�������:����L��d��y6��ڬ�ٟk�X�":�� �����vc��V��w}PW�wഌ5�6�ځw���BmJ�Y1��J�����V�5#z*�_G���n���Z���j�2�VD蚨� �?���}��*��S�=
��q��P��XB5
���:R�y��9]����q`����{�%�g:N�@K���s��+����бN�E��2����{�J�T�w�m
�����=��>�Gv�a�8$��Ö�>p��TLG��}r��6�EA5�>�	O�@˿&)i"�%+��N��ФpB�gY`����	��|�ֲf�8D�4#N�95قu�KVkkHi�þ��1g}>XC]���6�������ӊ�}�Gv���4K����V(;�E�C]D&�z��1��Ĭ�s4QY%��R
�P�?X�4�֬��B��ks��oՅaVz���m�4�ޥm���B]ܥ.��N���A4��٘C�F��y,J����*�@ ���Ow��=�Tŉ�ئ�u�nBqD�X׌@x����w��5IJz�K�I��O**�a�QW [w;yR~�b;ѩ	1�/��,W),Xɮ���}Om��l_���*�xs��E�1�x��
s�#Pu�Pf_�"P+_�:G���Y@�5�b�������2 �gq�&E��Hk���gǈP	:خҐ��xB5K� ���坰�e���O<��G��T�wm-+A���D��)�|9����k�v<�U�x�)tDM�x��K���	��:��E*m��\�z N��u��!k���Lj�(�Ƀև�?��>�F�x5����&��\��B�u<����C/X.cȴ��Q;��#����V���}8������WB�g�j�]�_��3�$�+�z�,����H���@,6���q�ԩ���Ԣ��L��JY*u�b�9t��S�m�fG�kZ�<kkuP�C�n�Im	iI{�-0�碕�<'�\�]V�ڏ��[����")�#�[&|��g�Pn~E�I�
�#V��9�*y��l=���s%�O��L����%�;חLU�77��~a�^6 �l�֚@��K��	���}*?X��&�*%��] ��I(\ߤ.�#��ә;��������1WU�^��E��Zk:6��mϚ)�N�~��<, �)��~���iZ�ߴi:��D��l���Z�Ӿn�����_�ldʏɯ?�mZ�'i�m��
�ǈQ�y����y�T��7/^VGf�d!�·�a>��S��{�Eڞ#�C�K{�#UG�������Gڹ�	��kE �Aλ�X����;�O�]�68<�י����iF
�ee���?����U�U���C�����DL�2��⛣��}C�����N���g�����W���jl C0�+��雸�s^8�cHo&���\)��)� 6V�S��[��o����Vh��u��U�G4ְ�Ji1@��)q�Է���w�|pb|1[R$�ߙ�K�CK�x�� �@g����4�q�OL')�'c��]g��]�S�p�ʓ�"1:�Bw/���H0:�����%T�)6��ʲ$mf�hh��/Su�2 �I*t�w*��{��PI�,ɏ;�5#�fV�B"[�v'f�-�}��Z��n���sj,��lh��ݸ��fK��#mo��zW!sxd�����2�z'�-;:o���x3g_�ĕ� B%��_�9�pHᝧ}�^U����P�A�N����o{�*/��S2�Z��U�^R
a������aY��z�w�_af\����W~b��ㅌ�!� ��4.�ohj�Mbp��C
�ޠ._��}i�4�n+}��i�64
�{��]�2���a��̖:[�`��r�}���:_V%<^	�1�b.�ӹ���|�;�#�ѷ��Ʊw��6��������a�wѫQO�匩���4��b�hU�6�c�:��9���hW}'�f�Z*ڂ�ߐ���: .��;ŝ^^����܈���9iʪw��r�F�����[�?��EX�F��x�rt��XClK��`ˁ�6Eu%#Xb5^aœ�>�ڤ����i�ut�#z���(1M�"�}�[[=�)�r�)������"z��웝׈��G����8>��9��q\�{
N�+Rz������Y���CWۿѥ�I¶+���{739���g�to�^R�����J\�	1����}J����4AY�!�n�V�5�y:-�5�y��19�6�^�߫�;K$oÏ\5t�D�*�2ן����4�n�F��+7���!K���-�W ��5g��/>��f��#�BF��"b7�C���w�ŋ����Ӵe5tǋ�[�Ϥ��|q<ڳ����V7�����r�mFx��1�O��=��H4"�W�qt��Bcݫ:"�'���H�9V�`(Ʊ>�F�<
���nC�b(�`H������Ӈ6�D������YN$T�M�a�0 �;��z_����)<dů��0��I���{'��$�/w�S�,ٟ&����� 5�ƦCZr&��]u��Xz6ݔ|� BVeQ���k�-�ta�"?������H�A&�����<?�|KL-Q�\�8�#�"�B v�.�=��[]h��m�p��%$������ݑ�Y�j�/����O�o��������> ����(ajv���	���ʸ�+��?��o������%��Q���Ac�VOHF�������	6#q���	�	#G�>@H�WY�8@4�dd4f����]РQ���Z;:��N�u �E�`=4�ZOʥ|���FC	.\X��I�U%K����)z�e�Z��I�f��mx��\T�ܔ>�Nz9fŹ�� �A��'��$�Hp�A%8x3&W"	G��V'�V�~?$�h�h>�5tw�/����g����*]��s#1�0$���l��&����g�W��浘vsǿ/i��iܝ�7TxS�O���X��eJ��.���e����FfF�ϡ�lw�=D!�o�;��i��⠲����)�6Op��P���̠�e�'��q�4{����㚒��B��H���uCC�ly(�0���0�Ô�KÝ;jO����ݞ�G�2�(���?���h#c䖑�_�rWq� $[�Ld#���G�����|<Կ-�$C���\����9�C��;�ԙ���m��wF�T��3�zW*��	VTA�:��ݤ����wI��G/���4�O=y��t����%�vd$�P�1:X�]lK��&Wwi����&J�zVo�9˪�)�r��H⌹L_hg����?�f	���Pk�c���ݹ<7k�ptT�QNc�8�3ԍ�p+{��y��/�D�FQ�\��[C�����u��J����nR<*Si��j��1�>�48
���Os���)��МSv���Y��aE��
U�/d�+�Z��o�9c�	w��d���۬��0V}]C�,���Gڠ�Z,���;��S� �J��w��^���S�@��_�E��p�&Y���շ���m4������D��>��Tq�S��v��*]@P#K��gQ�yPI6��z���ͷS���� ��{�R�i�@4>_o�e���0��2 3?��e�r�͌���?P���)��E$}����Z*ʝ�%*޿�.Ƨ�� _�yŇ��&e��c���5�[=�sU>�gfu<z)�	�^D�d�F16=p�{dB.by�a_�����LK3��&���'�����h˞�f�C��y�+o��� S�\Z�P��e��/���u��?�
�w�e����H܅R 2�6�IrFE(M��p�]��P?�����fM�i��0.���5v'rf��cQ|��u��p@j�1q���^�3�Gf�Rb��Փ�<fZ����h�e��Ϡ�=g4>(��"�0&��e+�'%�$�L�y7���[���޿oP�/�eTb����č�6�*�;�8�iKeA1�&���a���l�xt���k5��)"p'a���UjBxw#�j|���+_Xj��<�.1�ܤ�UY\y%��QOA�oʫ�N�k'�:�԰ߜiMR���tl��@[�6@�y�t�321�Yu��cPΚ����N|�i��8�t�O��_�rxi�R���X~��<@����H�'�!�Rъ��g]�*#|In�i�\���y������Pr� �0����6eK��8�����TC��1r�~¹�|if�_\�q3^�|�t���s���F�� "����v�T�m��)'L��I���|x�1��������o�C���ׁ�hQ�����`����;U��[-l�� γ��J���X� t�#�h(>�ҧ�I<pa����S�V������w�J�z� ��p�1���2���HAv��n(�a�������}�W:���qMA��,��@�}��M�~9��^�Z,�8����{����z��_s�ֲ�N� ����v��'�r�/�`�	O�?S���Z=դdg�m�Њ��db��!��3�6�񓹽�ȣ�!V�˧!�ՙ��Xx|�oy�<���c�(jn�n�-(��H������%�sO+X�C��y׏���b�U�@�j<�� ky�ԕ�_$�'B�Ԍ�9-fC�"�b�v��r���~poVsoj0�f]�=�{�?�{RS�x�"�*b�]l�B�ŏ͐ 9���+k]<����(���BP�e��eE<6�mnE��[EN���x��ܾ�?� �4�(�i�Y.u#�g���	+�n��,��u)���x�gc��rl&;)m݉���V�V�|����QņK-��t��%E�[���������,n(p<�ܷc��4�,Ofs��B�>�;��[��#�����UK/�DC�]+�p�N�)�<o{�t���k��������y}�^�QfsuyZ�O�&r�e1��bo���/����kf���mO�d�>�q�X�����[�V{HG��6*��`Ƭ/�Σ�x�>jU1�*�Pu)�:�#���g�
��Z���;c��zV�$�ϩ����q'@�N�?�5ڂ���������z�=̡�#_���:J��k��[	)��v�����,:<�7�\#���޹�9YG���1X������<e����gK᠑4�l�:LN��FHЂ��`�5��q�� 	n)�;/��ܽ'uxz/=&B9�S!�?���������n�B����W�h4M���ev�?V
���F~�=k�׳���:2{����[[D�B*�P����/���)F��|_�T=�Y��D����bp�(=6Hk�8��������TmI~�g��\"�M�X��|�}�>&^�pE!��6��eך��C�`��b.��N��4}�c)��JZ*��mkD�u^��,�/�IE,�b��Î�G�a<E8x|:wqO!�(�$��(�^Z�jo��z$!Kե
(Pوdi�{��|����P��Xz}ڃ�}���/M���@Y����+�(�И�Γk��� 7��ι�`*q]F'�j��L��:y��X쒀.q:�{.�{�0�c&)vv%�5 +��Ec]�ڋ &瞣�ޮB���ŞG�t(�٨� 1?���}�e���6�2-lk�B��9�]t�E�Fr�&T�5��@�I����B��TM2��5M ����������W����m0�����7����Li{Z~������T)���ۻ���{}����a����fR�0J�`ͪ�rK��nvC�G���Xa�C��փ,p^�T�'()�^+�}C	��Y�pﶡO���Oz�*���1�L��=WT~P�a�;a��˗˥� c��տz=��N�(s\�A���c�����,��[�@v��%@(~BS�hÊP���6
�D�%~�#Q�����z.>n�Z�4Ӵx;����L��~9 >� �v*a�>w60��rc[O�p� B�K��ڳ��L�G�/Z��j�7�VPNsȆh7�w�uw@����ׄ5?Q[�3>�5�\�]_s<Q&ȩzSe�!�P;���/1E#��.�
(4�]����������ugp?��e�(1Y�*Y�jx<�5SJ���dҁ2sl��D�<R�]�Q���m�;Alg�}SZİ�.�Lvu(�N�%��!�		 e������Y�6�I�B�N�}�@���^d���L)�ug��%`�°�+��H��%+J>���[��c�i��n�Fz%#T۲x�2S
�����V�Ȕ3�g$�y��w+[���"����� �@�D�)b_ɺ��`�š�,�q�Y�8���@G6����O	���1�~^���7r���1��,�r�� ��yp�r|*�IUf��WZН��\
7��q���<�_W�.>{c�j�ߤ&U��ҩk\���;,nz>`n��6dX��euu.�,x���F"rz%�aBF��'&6�Jwo�M�70H3B�����h��r�a�׋tiH9w߲'����૊�h�uF��,��ۛ��@�$���t� �Z �𰵴�Ү!,�R[�?9kQO���J�Q. ��U�}&/�_U&R��Ȑh�IL�����fv��7�,(� =��0��C�ts���t��AIv�n���Í�]��7]����e>����#�P�"ce�[��o)��G2&����H�����}���4�3qͷ��C��fKE"�]�ڵ�X��^�i�̛+wD]V-���V�T�S6��Q�B��KύH �Y�mI�R�s؄��vj��,����j�48������!���l��x����*���P3 �B��ۣgD�e�� �d%���)��C�6㊒�i��t�0�;QfL9Z|Z����Ih��UR����ъ!ϗ+I����,e��h������>�/����/^o�*���'��P�ZJ��Pα1QQv3�gN�L�.��'w�X�~������p�9�b�>�(s1ˎ8�����p0�RM�ȋ�[;�a�Ӯ�`S'`KZ.��J��z�k��Zi��YN���<�I�W��t���ͻ�	#3�G��0 ����`mM��Z� ��´�4�ob�$
�^ m�e������{浌��e��̘e�xY��v��y���T�^J��-�Q�O��'!�v���	(�� h-�~���X8�-h%��Q�[ɉ�h!8e��e��gd���$Fj?�څ��q�
�ƔnX�L����T{ SVe��T�r�Nt�#��y�$�����giu�V�Y^8��<7H8��]�CX��w��]���Z��}["�wfn�P"泦�V?��Bpa4�js.Z����D�7��vL���d��Tx5��#�_'�O��'Э�e�} ��ܹKi�|���\%|]9$����,S>�����Hy�Ѣ�����ƑB2���>H��.v,WK�0����B��?���?I�T^��?Z�ǒ����������z����+���G��h()�%J9�Օmʘ3�7
T�LV�Ԅ�;��P��
E����v����T|�d�Wp2W�uvn�$�����a�Ʃ[Vm0,�4��痁�w?W���ᭋ��S���S���NZ'�����
�����jp�$)���0��3��hs��6|5�F��Z�!�Ѕ�TT�uA��y�Â#~#�J��%� �������&aW��g�Z��*��^�:#A��/�AN�����"�q�L��m���F׫}��x�1zF��J_��A��
g�T5��6@�Co��_Z__��� ���4�� ��3JI�rͭl�8k�J�B�	���1a�Բ��-p{�`,���c+��T�;��5�3��ʳ?��̡�5iQ���G�\&D T��,�s�^p���IϢ#W�1�f�6��e��"A�<W��X$���~�?����E0�P��U�$�L릮c���We� 2������L~�V\X]K�u�k�{�oN�l�~�L~��8��F�B�Z��3=Ӷ���q��2�^bo`;3���������j�����愹�
 :g�l��\���Cy[��d��6��>�!K�����*�kz�Ԑ��M�&�H�|��=Y�Z��,¤HZ1Z�7KbY+��a�������;Cy���&�9@Y�4ϳ�Ϫ�{n�(׍jW�֪P���*�Nl}δ, 4��s�f����M��7�Z�P�j�c�2/�='��b�V>�Q���2����焃��理A*��G�s"E�h,�y"�?;���ʈ�d����;�"��_y�_S��^��A!*��4b�9�d�鏴nYK<.�ѽȢ�L�:9�w��0TQџ6^� D��P;��/��*��珲�g�@M���㟺��sX��%�U���[v��^u���D����h�\ٷB��Z<�2��"���A����R��u��C�@*E+��+��N��St(��p��]C��(&���Хi)������!
���۝�#> )l��Ҭ�rÈ�]��V8�vȀ���cz}pjG<�G�`M}���1'��S�'��CC/��%�*�lG�F�أj;�P���ͳ�����&�}_�,�"�!϶�>)L�=�W�(5��M#�]�N-� D�`��y��݀�(��E�gײ\(�sM6�ė q�y�f� ��� ��f�3���O��7e�Д�G/�9N"F5��?!��Y��F�3�<�ʪJ]�����$��5��w4� �Ve0��[/����n�Ld-iȞ���.9*���W�6�ȕ�%���i��R��� l�}��
b��@��ڤ^~�?��ўh��덖_�L�W�xF��O1�f]�X��87�s�#)kB��������='^��#S�&ٞ�7e�'[��hN�2$�{fЁG���2�4��>�ع��S��2J�R����TzW�c*���Ta�'b�*��ֈJ�il�8&9K�S�3����p�p# :��%���؛}��U%�.�G���6����ЊcL��-�Rwm����;�g��%�sY�5V:�m��S�����_��h�M�j�0�ՠ|���#�Ci�?@~�b����DB�>7�5bw��u�W���X}|���qܭ��4l�:b�x��퓿 ~z]�d%Fc���#R���t�*TB�dշ���n 	T��[N�	7=��&��R=���8���R�R*\�(q#B� ���������n�㒁���,���ں�|D�� 1OJxk˻3{��gO��=x�}B|eď�f�����%�7���E�K�����K�$��B�}-�Iw"��eO`C��@O�;���_��P]���0�"�ɾc
���89���n��w:*�"L⃷�z5��'OH'�������v�r��@��H�&��	�'��w�8�,ؓ ����%��4M��K��[���J[��,�����Φ��/M�����ow^b��|�4kِ�!��C�I���T��=�A9jx����)���bqy;��ۙ8�T&���=3���H����o���yx��93����33riڒ�ݸ2��/pݩgFϵF��~	� �����/U�S�0�;���V�Ϫ�!4�5���ˎ�[ �P���0�p�*��S����X⪝HU&l �[ax\T.X�,e�i���Z\:hB�����s 	�U����5�W�_8R	����+���5�ed�i}2�6x?L�XD��V*���H%����9�Ҽ{Ճ ���M�k\f���Vpڤ�o[:�߷�~k�̑+X��a���F�F��V��$�
�a�M1Ȉh��'[��ڢi�@�B�'/R]��k9�����gʄI2"�=dKa��1^�Ӡ�M��G@�@�8��6�^*��� ��)hFt_h�R��>h�Š�s����7@K-EE_�Pd��m��?i�Ғ�8�6i>b�Ȯ=&q���XX�yD�����q�G><kY��]@��������b��c�?	Vqb҅G����\�7r�42�e�*G�y^.�Z�'��d�2�����1��Y���g�Y��>J��qu���H�:�$uI��'5i�
��[�3��}:s�mk��O��|Z4L�ޟ2����)�g�.X�bl����O��:n�x��K�WH1Z�2&h�S��<�)�l��PE�c4�x�f�w_�����m7N{��.
U��A�D���Nu�Hȩ�� �Xї?���;x�~�q��l��4���6j��σ���#�@#"��-�⋘g�.�yX���,*>��Ljo� 8�5#l�ͮ���O���
h��,u#/J����f0N������ ��U��F�����'���P,�C�z��Y;M��GHۧ�����!.)��,E77K�v�j=�)��p�i��*��ӋM�Qъ�д��y�-���,���H����li�#gH�u�)���!I�e�L~��3ĶBҘ�޻m�5�VQg�j�Q9��F���r�(T.��؎/����c��2]�0�\%u�*
�,�<��;�:�<��6�Ipnh$���We��/��K%:)E�M�cj��6�5\�ٲ+�h���B�GIs�O�,W�ld?c�C	��7�����T�96L����w������͈x�٩�Vk �% r�$���.��:��X.Hۓڻ/tf��זּ'�#6���|2�DM�7���3\,du�W��O<x:�w��tg�������m����&��gf�'���4ʏ�0Q�h|��#9J���δF`Q�J�HE�̺L�m�`�ðpn��r���g�$��zL3C,�(�̈́ ���s|��O{��.�6����@*�\_<�y���Xw~�'�\a�v�B����ٶUPW�(�Q�i5�q������r\<.Ә�ì��1���x5a��e���]xc����AYK��7A��")��K^�ѯ@�}�÷;��e����*��
�L:#.W��ӚZ$(������g�~,���.Z�����{`M/�y�
my�F1 �ձ>�9 _㦑��=�E��x�
����y7YE���$Q��`7w')��F��*�����m���qY�"��Cy�X��b�	L�5֥�S��(��S�!ۤ(�٬�^��S�X�`S�	����Y)��	Dsk�yi�_2�U����Q*da���‒����
V$�){0
�E���quQ�[$�:�D����Z�z��_ ������vhZ��!�T�xW2i��%���U%uWD���aRÊm���?(�!����=�z)�z`�n� ��"�n��H����EO%U�d�G�9�z
�jD[9�LR��y�G1[v3ڇ��� ��k�+d����>q�?�sJ�|B�8!=����wUY�
� ����T�(�.��'�_K�m�=�6�6���|R/�<�;�I��/���1��j�7s�߀EVJ���6�J�r���.���U�׹u\����,���_n�b8����ph��:�a6�+a�"����%S�ޝ�p ��	z�1��]��,�v�{4۸��F���d~?�"�G�O7����+y��~�q��B��!=��w�6 <5�������8�V�f.��x�ɖ��Gh�O�4V*��H�v�A"�|TJ��+xʦk�2�B�kK#�/@�x�w��B<��&"�\�*� �!%+;vJK]������j@M@W��o�à�.��Ƨ�����,�]�� ��mWx�/1�,��:nhׇ`��q�����C���=�셆CK��/���\��>	B�����ڗ�٪��ܲ�Z�Î�0���Bs;�QJe�ǺҼ��rVSU�B���fbw5���ވl����dݑ�5E�Tɍ�y���x"%�a�I�B�d��N*�R����z�sE��e��aFS%���c�{k��e�Ϟ���4bŪ�9�'���$<X.(�x��G����a��َ+i���A�!BCKea��ٰ���㜒�!4���{;�$Fx�^��O��
���/��x�0	�=�,+�4�q�v���ٌ㼭�lϬ�k�PƧ�W�>Ƙ��O�>�t�,WC�=�8X��g��#I�dx�e�%��0{�����/1M=���4�=�=��]ƞ�D_Kuv����(���E���a�����+�Q��0j�29��ޱ��:͍^�i�(�^_"��� &�Z#hr��R�:�. s4�p'�Ri�=��2%�p���y������t8�&�Y�y��;7R���nR�ޏ~:c|��vJd���7��Zl�!�y�z�X��uj2r^��CjUxȇlG�E� dٛ�S�#9K��o�1�l�yH�_@�hsFUXw %&�"+�jF�����F����jx���܌�)�83b���: �!�C׏9`1����4�x?�+��!v�ڹ��/J������b
��"��
�  WQ?q���ΒhA� g�׃�{[g�wm� :'�;Yn��I���W��0���r%����@U�Q���i�z�d5��<�9�b���>-�@V�իv	j����j�[�YC��Hn18�iՠ�J��bhqE^&r����YjZ0=�Qp ;#8СI�nl��;Z��x��F�҅uj�܈ɚa<ؖ�y&��t��:���(~��sI<C�?}�ztn�J��B�$<�l9��h<��N�=��ǻ>_|�I�V�M]�G�P����ә?�����Nt��j>�b����W �f��8�i"jh��)���Q�r-�6s��ߣ�e�e��e�)*��������}[�+� �ULsP�`��Q�GH�:ӽF1�c�e����2���|��l����D�ʉ�?�.�f"��!f*��n�Z� b�����eT�RI���}�U��}���$`�؅��Y_E���f'��+��^��L��T��=xҳ����'M!��'�W���O�^&>@�RAA�G]� ��$M�?���j8�06�c��G`Q�~��?�=��v	�j��z�a��o��A���jmԭT)�<]�mVh�?'Y8��,�T����G���|�[vK�Q��A����J��u��4�g:{�w�:�a&t�v+[��(�E�kW�L�7w�P�[�ݽB�R(~aVP�{d�D���8� B�/#��u}�L��Mg���Į���\�G�;2�l �oR�y~\i´��X|��+�+�����a�ʭ������G�f$I�c��O.��n��F6i���+�UܑsDZ�2	�wI@lCꞁ�*�;���ǥ[* �ug�81�}I��h��Y���v��`��5ذ�Lb��,�r8&O8�m�)K���+y݃�7��z���_tD����e�>���$��髶;[|zbM���h	pJ��\�ޮ@�b�p��Qay]��������h�V��s�2��}<OncK���m������'�.w*+��
'.(����9�q�ߝ'���y{�f�c�``.��;�l�	�Lz{��SFP��-�'�#ݦ�Xt�!��(���V�&R�ȿu�:���Eװ�qM�Z�%��/x�5��ZY�k� ��ɗ�/x׳��/z[�'nV��T���Q�K٧���Q\���|M�B�|��m|(p�� �4�CvܣQB���`�u�DՐ\W�8��ʺ�6��d��>���$��ۣ=�6�0�D�|ю ,�7��$�i��r;!ꠎ�p�@¦��-�M�HNh,�P73�Z�<U���?���dc�r�C��E��#���j��Y�W��j���+�pmJ1ӽc�S�S8[GO���2bt�sqޅ-ɧd�F2���^F�r��"��%Bd�lɼ^�%a*��:��`kh8�Jg	!���0��QEWQ��e�f�2��,�X��v ������|@%X��ϳy���'�lC��v���JF�H�G ��1z��͍A4���So�V�� �y��׸�)��_:��&m`<d�E/8�a��|σ�-k]>g�o=�����5����%w����8��CZ��(\�|�M�)�C�Aq��$io8�:/6��Cơv�4m8�߯D�ȼ 1ib�n�pyB�d�4B`@i�_��G���g=4��l��77x8�,���(Xyد-l{ىY�� �r���t~yK��ˣI����.�P��J�Y\�X�};��� ��x�KJX���bUYG��q����K��&��"�>M�gv�ʑe�!��i�u�7�~}D"���^�)㰆Woo�G��ӗRfv�����fe9�3���^0��rN���������L[�L	��Vze� �R�߁Հ�0���8u��h���L����q*�l��y� �ۛ��O#�M���/s�W=6����WQC&h鮶;佊h�c����������?(�"j�j�`15�V<�g�;	�2���� �dKe�0HOh1{����%x)�I�R����7%N���\�{�q?G�#c��'�j ֭�_��_y�Q<2����	2
b��ՌhQl�Ŕs�e�q��e�@��.o`��7O�����-��_ZM��>�����:���xJ��=�_�����\\)&����5Z�Y�O`X͖���cRyýS�{�2�#���'!D	�F��Y*��ew�����5$mQ#u�?�U�yy���X��<�b�h��¶�Q�jX�w)
���x�vz�@UVc�%�HD ��ϵ�2 qP�Ӷ�����F�!�I���G$�÷��]���\Xˏ�q�L�$�?YHn����.'S)�M��ӱR�ǐ~�v|%�Z:�X�3H��ʤtޤ��2���z^�_3�W�U�Pl�E�_�(�)6��f4�5
Zq[y���L��f8�wK��1�b_�I/�Y��bZ�$�%޷H9-��|��(�d�u���].� �>/��������\(���8$<Y�����Ylt�{SV��^S	E�͓_���� ���=���.~�r���v�C#�r���_�|��Kp����_�C����?9��mx~8�����@g��V���Qٓz|�d�#8���C�vp=c������N�,���e�2�{&�o��%)>(�4+�\ �|�>D]�F�r������U	�����+u��@���^�.��̧�4�`Î_��L��Umɥ����o8� �'����(|�wR$��&�D�e{�F~�&���4��f�<#���k���Ŗm�8#/���[)��n��9�af�b�kV�b>3�[�,� ���B���{:�����u�Ec�T��%Af���x�+��W(��g��@���g���z:��袁K�[\��&�ft-�>\�备Wa�ϙ!/���`�j:���������3��`(�.���|R竑[@�|�F�τy�|�=��fp,Z�����A;�k�c�l6j���E����"I�p��i2ͼG]�i�cש�x};*���`�L�tW|)��B,Bu�R�!#�6<~�|ƴT��,��q�L�%�9�h��9�������'�mZ�̃�h	V�#�:����K�0��J�(�&� �b����W�{Q��EJ��A�m��4QW/��O�4Rm3Q�)D�^A���;����<����r��Ǝ�0_�nm�}r�(h�����o#�e�w��u!3��h��wq�b����ыܧ9?Ӻ|�J�R���{�=���s����jq�W�@��2'��=z���!v�j� ��}J�N
R��֫"Y��Ƃ,C{��[#��i�>zYOj��.�b�����Ŵ8�C�2���JK}���A����2�ioC�|BpxPw��E9����؆�`2E�����ל9�l1��wM��'�p���K����w�wL����+���xl���0���q���Q|���)K��*�bH�Zc���Z����Dc9t��پexOI�"'���60��*��ƒqH*��!�88�VN�"ֈ��#����r��4ZN�@��Pa�����3�e��"��Q�|��b3��!�ߋ�n����Մ��gaQx� �J�[u�w��g�������ڷ�F�v,`�L�[<�B�����9��.2b�:+~rR$P�n��2������x��;"o�zH*��o�3�^}�\��)m�J@\~�C����J~��q�鴂I�� mR�lo�q��Z�Ii��/���	j. 7L�e����/<�4L�<H�wI�sr����yLc�?j�m� ��W��r_�h&��"@T����.n����-R� �8$�[�|�sP�h�/P�l���ê)1XbQd�~ �5Ͼ��9����d���uۀk������U̟�&' �@��{dQ�[[փ���*�SN٥n81ڔ��S|ӤdZ������$��i�zV��_��.�x
e��p&<���g,���I��m���Ց����U�H���p���U��\�}-2w��
��&XF$n{�9�x�nҫN�B)�̙U�պ��R��;�'���@��FY�[<���RE�	?/Gh�Gu߶���TJ�h6�e��Z݁°�����y&��������˵�b�/�P��+<+PP��㿰O,ŋ(b4��c���6J&Ɋ���n� K����{�+S�b�-���>��Y�xvO��1��C�#�<#�#�Kq�a*�N�$|��=��5H+y����&9�������?�ea����f��T�_%��������e�@]�:H�sx%���=��$�ъf<�#(�^J�k%'�j�=nk�t�w�G>�����{}U�t1�V���L<Y?)jN��0��Ų��"���	�b�üY'ɪ���-k9��gq�6{��`5�fˉE�R������v���A����c��rTm�?4L����U����!q�1�Zn��vD7yP�)�:�Be�U�F�_�_+�ԏt�CyS+w3堷RkR�Һ��G�t$T��8����%�B$�;�G��TU�خ5��
Cj�^#i�j�Z��<9X�u�_Y%�]��0��$��|���|M�[�VKA���ɬ�>�ik�|�}33�@y��I�뤊5�ș�dE�7�Ʒ�C2��j������/���%�Ҟ�R��>B����`Nҳ��b�*�L���Y������Oؔ� ��W4Qg�n;e�?)��R�	�
�|�˽7���(��[�]X��ҊkU�7ۘ}���i���C���ŽX��5GB�:ˉ����9��o�D��O��}�f��L�s/��A����e(
�*q�'�ɺ�/��!@U�\�n��n�9�����l�h�>`�1W3�}(��T36�\>0�L�iĶ�~,U��	�ϡ%g�!����*#���5K�VУclWB�=��r���z��C��ξv �V����#�F��hd���{Ń5@�]Og���9���e�1�y�q,�~�{�U9���Y>-�^�/��zP.��P�0F��RH�܌�7���%OiTy��$B� ��tl+��_@�� ��wb���e��}(�a���(UmOZ��B��@-w0�����d��>�^ՙ1P���rX��/w��\�w�T8�@v�Z��nW�6���Y����M���H���u
S�nx��k�f��7�|�6��0gU�#�b���2��O�z+&yU�f0Tɇ��@�������VHa��=�C�{�����?��/��c~/i��v�a��J�g0[�[Sf�`�����Xa1J1]ۗ���dh�}�l;=T̟I�׶=���w����*5��"7�7�>������^�A�����5c��#S�W㢂�CH��	�W$�
&U�F$�sUH�\����7br)�N���j.�-�w�H�yH�+<	oe�zA���vS�9�)�L�#o$gH�Т�UF^������
�����݋v���Jf�"�/¶����RdAR�Eb�l���A^(�&#��@O$��OEk?�0�Z����i�h�]�s����\��jiĳ�[~��?)+<�~���W�ׇ�+5O�0Ζt�c�J_;'>0K�F4`�cr"�Ty��1�m�y�޻$1�X�|�g�4��|����rG�|T'���A��W+�\��-$�,�]Ab>���<�tP�3Ե�is^�/�&����su���&�v�"<�;S$�,pL�R~l��o��U�,p�/����^�[g�LAjd��#�	��a��3m
��q9�	y��i��l	n�]7vX��i#����01˅��������9RL_iɕ�:C��3t����V���HL!�����0J�_L(�X7;<�g�m7�z�E�^���&H1�������e[�����MA� hCR�,��L@%��S�ғ]V�zs�>1�����JY~��0��q3�	�$|����jy3#��A�t�R[.�2���)Ea�f��J)�Y\�#Ι�g�fc�*��4u�T���"}F��Q����H;9/��.+/`�Wi;�yѲ7Es�=9K`� �J����8�Ue���(V��
q��,�\�[�Yv��R�%�B���{�"�j�υ�A�7ǳ�Z���A�<�F�}�y�E�ΘY������$�n)ũ���d�f�Vܜ~<J� �#�2,elU�&6��9Qޛ��JQ@�;!����؞ݩ��j
�;�1�B�����i�h��c�+�����U��R�w*�R�����L�6I�]�L)�j��q�H�3l�=�G)�f��]��!Z
�vH5��� ˼_�b�*��+�olXHm�^�[����j����
�lm�~�aw>�zl:V����I��.^.�!�u�F�c��m���Φ�0�'nx!���K㞦���._W3��Āg��Ԡ��9K.r��M���)�X�ղj�.��n�|4�1\��nC�>�$7�,҂��7�-:M��Yv��l�R���A.�~�m���\�,��@���s����+Z��5�����ȉڠ\TI��L�p�n�K��o1���'=�5�u�l��kHƅ��wVX��� �����v;'Y�'@�����c:�u؃?��Tْ4!7y`)3����R�E����1t�,�6�LӨ�kq�x9L�+�B��Y&f��4��1�D��s�Zj8����	���$��j��[�=`O�[9J��֏��ܣk]�gnD<��q��}�1;�Q)�o,�6��벇��]Uݵ�r�� R��(��{�d�"�f5t��§�z��8�6	I�D4��z��΃�=ZZ�"����;r1#���YRő�.l��?>*)e�0���RY���h[b<�:��Ϯ�����/<	q��/��=���Y&���Ty|���
�Z��<�����g��X�r��m�LӸ, h�o�$m��Sm��m+��tS�;�U&',�P<�������!Ͻ��I�nwyal�#u5\�R��Np����ٲz�A>��j.E,�7��ꎺ����6��$kU��:�	ȟ�w)<�BSS����f^�-M����b��u̧�崼;h��dL�	�S�u$;b�:^�QZ��l|��p�d�i��k���,k���7F;+��s��9�����"�R�NV�ӗUa��v.�|� ���#�\%-�v\�j^f��2�k�3e�ny� �Rή���I?���hrk|�W%f�ЎI�ߧ�[�f�l�o1(G��
�����W63o�ca��ml@ ��cH���l\�L3��	�ϥi1����ʞ����u�pb�-%[�~��}y�Z����m0�{|$����!x�H?�B`���O�_�$��$��*��fl�i��0�q�"���*H����x��ןHym��٨�^*�̠��m���G�(\��F��s&��!�@G����G�;a6H3�()��E3���r}��!��DM떖h�9�%m!�D��~��_�Y��'5|���Π� r�˘�Q�V�)|���mBK���N3��r5ފLj���z�
B?�{���� <aσ�a4����a�v�8m}��c�O�L'8�9︪�N��u4�蛰�E50v�-B���
	i,̞����5+���@0ss�ꁇ����7��	����K�x�ȱ�nf��/�Ԥt�hs6c���x�X{=N�t&�v- iK1F�Ĩ����j����;K����?����zq��/Nb�p=6��.`8�D�M�Th"��=�L�Ģ��z�]`�ċr!ƺd�삅��`�CGlV�&X;�z[j�>��(�/Z�:\NrN�R`5��d�����Kv4A����R*�����6��b#>��X�PQS���m\���$'B��z9\ �F��uAǖ�S/ߝ���0Ê#5iy��:�,VQQ�}��a�k� T����s\�WTu�7���"�q��1�4L�5���u]��\��^d�T�}�k������-��յ�@5/�vz�z��|���/ك%D�c/U�o��,�~f����Պ�_6��U$��n.3a@�O�c� ��!�]`Ri|A	
4�~Z�mBJ�O�_.�)hjf�[?mt��3W���t�6Z��`@� }��t����j+���~Ѳ�����	1$�p{�}/�J<��9v�5�H�!gNt�p.Q3�B�d��\�So�Gu��_��EB�}W���${u�{�gy�o�`������u+B��G~`y��"�����s��s�Y\�|Ҕ!8�5�(!V��G�qD=fز�W������A&;+���l��mF?��h�_͕�]�)�_q:L�V����˲������ h:)�J�B^(��Wz���Gr���27��yU;�g������ƺp��t�$�I��?���3��\|��\c��`�jODC�����Vs�q�1t���DE��i�������D���@�Ntś�\myP�ɾU��,5'��d���D���5`V�qλ?� .v!����Z%�%�i�3�����T��Lj"�4X�Ŵ�B���gӟ�D$y%���?�J���D"hpv;2��\J��a��FK��7@�s�Y{���'�V&��2��X��^���x��*�i}lĨC}�_����1N�;z��V�Ѕo`{�j�Ry$��3-��gnn�6��M&��1�	a�8IXدu7FLU�/��W�?Nߑk8�G'�#9����:�v��K�w��ui� o������5|�X�7<���הzU~P:����w��n0��C�`;�d�� #��Rѧl�]� �F�z���CWL���~]���<���&?�S�<t	2W�|dqb��/& ���x��Cp%H8q3��"��QӞcԔ�ːx�_Ք[\v��k2+Z�L+>'�& y{�RQ#��P`�i��E��8?�`7�#��3�U��R�z�ċ4}���)f���?9}q�n�8%�G�Ԅ��f���Nk��Y�޹j�,�.�c���S,�:Zh���� :�k;�!�-`>D\��+�{\�<��A �X�w�pIV��tˬG�+�ٵBL�)����q� �c����g��w	��Ǧ�5/F����"�'QȰ,�ħ�)��z��Ջ×��|��<�Gv?��S�z��FG��azΑ��贠����:_���zJ?�[�'uQYLU�u)9"-Ul�3�l.`×��^���C�1tM#w�V��I }c�f�"�5O٢���1�jN�9?Uw"��r�l'�y��d���H�̤��r���!}.�*��:Fڑ�iQ΄C�L��*��S쐹
�Lb��H�9(��B�Ԇ�n �>�A�Oi��zc��g��EnDR�,EԚa��>w��ړ[Z�H��6��s�"�{e�EpV���N�.�čt�'��9v���H��1�@}���>�t��?�g��]�ɹzqĚpg���c��z���E�h.�.���5�m�����I�_�H�����Zf�Q�%�8�ܯt�穾�����"tWp]���C��(�^x�gA�`�+���-�F��-��1W�Zu���Qe�f�Plx�=�eM�bŅ��=iv�DT��m��i�R��v���P��*�عQ�z��84��k�3k�����F���!ӧg��ŇJ�F/Ac�
��Ef��ș�+I,��5����b�9t���>~g=ٟ�9�e4#��~����b�։lw��\b�N�(���p8��w���e�إ��D�ayє墱�$�	�v?����C�b?����rg��=�i���cB��3�B�9��åBj�~��|���LB�c�zG��͑���Ț�]]��I���������YJ45�ۛ��aW�"�DX)fJS���~��;�G�I"�0@HHD^H�
e����>B(�.)��g&�LS;T�P�/�m4a|��i���p^<��kj����W6���K�e���S�"Ʃ$�X�/S���HG?�*`��7� ~Qe�=�T�]2GF���x$p��!��l#�)WuZlu�c�����Ռ3��Φ��؛��-�`E�'fB�ci��q�\�_S%�3���O�Uիv��<���M� @�@�+�g�y��D^�T��&��+s�N�R��4wD��V�߲��Î��=c6�Κ�_C7E����C�(�+$�*8����_�dV����>� ��n�L@�p	��4������w��T�Rc67�7�h���I��4�o�ʖ�	��2�z)��8X= ����q���C5)=O�����8X����I[&	�rs`��sO NB�7�������H.1t�$;taF%�گ%It�S�}���j6B��9��������0#R�.F��q/H����zY�����hz,�*�NU_�i�HW��P-����!�h���}��
�����p<p�z�~�5��m=�g[������V=S��6.\�u8�(����^#�FV���Fz�����dB�w�ԟO�p���dMT�a�D�M�d�Q�"�������%�K]�q�����7� �u��z�+��6Mﺝ�f"�|&t.�Q����z���k�إ�Z�@�UsH�B�,��|�{� 5]>όF"�WH��3�b��In830���5�s�y?M���pׅ�����I�����Q*9��d����(3�x���M��[�ٌ��[�s���fɒu��lq�N����U��"�+�c6֟-ra�o��!�Q�~�=���
�b�����	`���`���w���p	n��IQ�'f1�W������ل���f%����&e��^}[�u8L��߱�=��}cLz����)��
3�����I����e�F��U,7��(w�|�H�����X��Fe4���.�h���'��nf�����ݰ�Q|��f9�']d{ck���� �o|z����vo
p��H�ψ'�0�XfUB�{%� ���C�D�a[4�\eT�ʒ0���!���#�Մ}�LJke�C���c7�� �b
7qX�'�Ü-l�iP#�d���q�yd�?Ӛ�(����[g8�)��Ꟍ
Ay�N�����������*��:f���]���p#Bm��_�D�����Q��8���y�`��I �&��v@�V��R*�³yw�F���絘�o�P�i؄5�B"�T��5y6��p-}�Ή�+��D)���S�[���Ā`��4�0�fk�F��=�TU<I5Ѫ�!�����hj|���涁"���a̳����g�eŔbu�B�9�kS��Q��+�pER�T�=!��?A�����3���.�ef_d��{�\Z����BICa��q}n�(��}���	����c��;ŢI.�O��m����|eCU�Y�&�q�J�?��rNB�=��(-��/F��-N����ʹB���Q�"c<�8���x�Fݲ�ݨm����]���^yI�bh��aS��p�kg��'����7���}��������;&7۬I�<n���%�;y�&T��A����s�p6t������ 4����[c�2��4��e���5WR��~W�7[O�M^��dz|.�o��ԋ�*��lxfr��)0���SZ��*- 0p���]�ؒP�@��3x ͟2�%�V�-Tu� b�n
�9�iV��_A)�}jv����`a���xP~ ɑ��Q������w68�ˆ�H��@N��@i�i�&�k�F�2��7�/"�uy�W�����6��4�6>��N�ޯJ0��V�]H���o�uw+b���!T�g��	4Àl�+ٙ�^F"lБcN�f�ɿFo-%0��%wb�v#�k�J��)�w�Nr��E^��S:����	s����#
i�J0���yg`�[B �J�H�iE{���W# ��K��&t�)	��ҝ[��2
��y=䤜f���:||�����M���܆H��{�I�Vx@ �`�H~?yPs���
,��.4��=Nu�7�v���,�ܒ>�j���H�l2�6
�)�6�����|�"���h�%�ύ+��m������fa��)���������p�t�k�����PmzR���qa�H#&���w
m��	ǟd�ѳ�RĄw\��:M����8ˑ�i�=O7D�*��?��+�g�/9���ԘQ���[�@�~��J(g1ϩ�|�ou9֚�	=k"��:���mYa� -��v��3U��͊F��7l��_�<�s����`�S�z��N~Gi������7eM����q��2���X�6�3%v_�*pnn���3vN����Դ������u7jw�� V3I8�tgGIB"xƿ�q������̯�Z�8;��!-W���'Hz�^b1H?����og<�#�m�G�q�=xQ�DR1a6��<1�l� $%�Hn2פ�sm�:L$s<!G�42�/΋E��|Wp�^���-�G ݫ^���7���$��
��7���A��r+U�|�-bѮ�kz�>��%�mǳG��HS��Q���j��Tn1�#xm�kq��ҩ\uwLE�Η��{���1,�O��R�����~8j��A/��*���M�f�} ��C�Fπق�z��E]6��ikJėJg�Ϩ�ñ��LJ��T�)J^Y9�x
���{�bt����R\���^ٮ5d%N��w#���@�
0��u������������Q�����CLCp�������FOvяv�����1��/& >��9��/v�<�g�҃�~�f�)��٢<�r�fa�x^�U�riń  ���0(�g����}��y�,��a�Lu��I��#��6���Zd�T�/G%5��v�Ml-\_:I.��mh�.0/�#��ⴑL��D�9X�����%�E�`A��]�Z�m�.�����e0:80�9���a�ԾG�jfo��U��h� #�F�E�Hp��Z"�:�J~ӭu!kR���ǵh}���UQ&�Έ�������$ǅ3�:[�&�C�����A�n��,+����㚘�vCL�?z�a�����5l��zb �`A��R|stid�#����[�_:�((8�Fńy_�&=��q+*��@��nѪ�w�k�#S�<���C���|�b���ƌ�S��VfJ��1�W�d��3�w�ӕ�?{�n�WORJ��T<{PB@�B�>�OGw�H�ǽ�*i�S}FA/A����='�NQ{k�jX���f�:��ҵ\	�*��O�y�3���odʦ�k�al.I��&hgi+��a7\�M�<u�;�k�~4�9�v�y���BV���Js�'y0��~��+Ե7�R^�`V���H�_�0b%�]!��n9�xQ��,_�Կ���I��
d{�q>sz�nfI"�gq�O6{t�D% Yg�҇�Ϝp�x�(�+N����1pZ�Z�(r�M=;��A
]��ԓ����n���D�n��)�0Ae������������DC���V���KoPJ,��	�q1CԪ~U�`��^G<�H,߷���B �}��@́x�EPl�'KT�F�XZ/W+�,'7ABD>��x��&��Ӳ�C~d?hxv��L��qbA�� �(˒�uS�Wj�/�
�z	�&�X�@��R*z�C>�&/8�g�n ���3	�~��fv:�A�O���4^����n��l�;,�Yk�1��.�'����J�4���myV�߮
��XU�,�Q�.�C�f�7�#%�@"�z�Df���Y3��˂�l�d<:�zZ��\��%�l�B�uәP�	�*Z�V밁��?8�������(��V�B�4�N�ł����rẙ�/���s�tZx;��.���oX��R/ ���;3�:^���	�ry�D�:�h���Vم��V�1Y�<U� a����DA�k.r��������s��]�ǜw3j9�01����A�"���G ��!�6N���C͟���:`@�~��3���33�	Q���w̵_d�*נ]��Ǚ��?��I_��pt|���R�"�
(�G%��߉�������ځ$u�#�-u��|*�mSԸ|[U�Ѣ}|ik+̋ɹ�5�������%U�B�yy�+
��O��/[����V[
O��9D�ŬJ�8��wY|tߠ��4��� �b��-#��+���!ڇ����H�&��R#)��{�#,f]����S��0��\wɨ�[��NF	FU>rDD<kp�&Μ�.*�%i.s9����3�7B�F��: ����9Y�*W�ݨ��J��:��?��hA��܏����a^�3��Ӿ�B�j8wg%3������vRL�@��E�]�P��`��������P�%$6�h���o'H�w�Z<�
�
7>���4L@�:�|����H�O�<n3������%8����*���U�������0���ciL~��C:��0S3� d��9�b�Ւ�Ƒ�9�|�"r���T�GG�X(!SN̄_$�1�և"�>9#��L�
����U?}��ݓ���$�^�)z�2Jp�e(``Jh��͂�E��g�D����Nf���J�>�La�lc��\�~��~M��>���<�3շ�"�������w�.S�����X.�,s�V���#�3�L
�9��uP_�k��Z��c;�vF��!=c�s�nv���j������ ���~�zWo��h[�1��~*n�z�|���0ٽ�6>4�f��*\b���G�m(`$]|��]��Y$͹��d|tZ��.���'�;� PL�T�m�o�g���L�h"��P�Ȼ���m��u'��ft�G,8���-�`�d3�>ap"# F����>��)`�7���.SE%@gs��-��<5�4���~��#֪�%�>%`�6���,�����۟ZΫ1�Qs8��c:��S��[]��=�a|�8^�gOpVs���������~qen��8��&��PI�}�_����5g��ĳN����{�%)͂�ާ�I�w�f���;C�plA�����y,�C�ʳ���Hm��Z��>�`v�ow��܁��i%��$RFEY�n�{a���^4;oZ�Isx���JpUHn���~���v�L�c_,� T*Z��H}����n��h�~�bNԡ�o��T���$�fSx8���}D#y��;�<P���yq��#:�j�{�z���5�����1y	԰�������nF|���C�T���,<���ə��#0�&��Q���	��ȵM�Y��o�%�Zt�A��(\4z��O%uUo)���	���"q.�#�L�x�F|��E	��u�Ձ��Jp;�G�l�4 m�LR���᢫LÁwa0� C�`Vz��,�	�bN2�,^z��f����,{O!�~[�ɀ�y�����Ǳ��J�^��t��2K�\����=�p�C��CF���^`ȝ\?�p��\���;�'���� �829�%r.Q?l*����0��c9|�h��^vUH�|�P�odl���V�M�P�fdW�ņ&=��s�7�a��0nZ
�b����{�f��Ԣ���K�+��a��(��oE�n�7/��'� �&�PoE��Tf�m�o�*�v�oi}e�Kz��jja|b�mn7"I�6�;!�w���9ŴvQO��bT��U���� �
Z�bŻ�B(1m�`9ga�����^I��b���x�ت�\}.�V�O6"������Z}�k	���L����9�Wf��۶dFW��>>v��Ģ_�0r�E�HQ�������_���r����|�o�/P�O;q%���Ĉ�u�Ls�g8[�3����P���3f���qo:��5?�����<���?�G=��=	 �n���Zٯ'�.s=����y��1�y����E�6��CmW�
UVX ,)\�[����(�Ld_�ʮ`k�:]��JO�6Jε�G�Z:W���&^��W��_V�����ҳw�78�e7�ډA/�������k��6�@�_�ˏ�6%�k����74{���ʙ]*�Ro[@� ���g��O���4�Rk2�TjT\�:����� !c˔�%��,�9m���{��@$�a�>�<6AG2�F����mq`�\tZ��в�LѽD[��}�P�(�x׭ԯ�e8݄����I�<z��YG���U���L)�'S��i���J�Rb�#R�;=�On�K0��-� 8�j,��n��+�>e�|�L�}�j5����x�L�];��g���L�"�N�!�-
���}j�@m.u��P3Bw�]��E�x���ā��Ҁ������!�I���F�B�=9|��wQ�� 64~�xg��o+�b�$7ə�3����CDħ�c���O��s1+��Yƀ�k��aoh+����IM�;�/1?��ȩΆH�;ȣ�<2O���\�f�?�d;e8[���
˩9_Q�r�ֺ��%z��静��Ϛ����D�-��Oh0.w�e�e�x��s�[��xc*m���JA�CS���'�Y����F�����ZxGP�I��j]l!|��W�XŶ��n�?)��F�,I�
�����{y�\HW��`�0I������䧱+�5O����^%�e56��1N����Ԣ=���<;r��i��c+�e������v}P��h�wǝ
������*�f��dȺ�	�
�4]&.gp�u�E���f�SC��7rKAƙ@8~+����׌)�M}g�H��~B;%�o�Dx��)U5�,m���2V'l����{�w��c�1�[��6��Y�F��*c:�3]�JV�����إ�#����lȲ��_t�!�����?x�_ݧ�yH_�:A����t�Ww��/gi������_�WgQt��p�E��䪻;��@�6w�>s��#w�h�?�ũ�Nz�]R���oe���%�I�2/n��py8�cOf�;��C,�*�d�i��G�}��yQ�ƓNa�͠�4.�sZ!����<o�w�k��)Jp�P�.j�<��.M��c����¯)�b^��á����0���Ik�����2ĵ'F�_����]$~�j�_~0����֣��:jSrj�.[GC�"Ű*s\nn<߮�foQ��s�]T�Q��@eV��QJ�h�57�Ix�=���`w*;4[�J�)w֧����1��>%Oz�a2h��Hl7� ;�s�As�#͕��7�X�y�W
u�E�$h;	�]+h�3�>�p�a���3�9u�ۧ�Q����y��ǻ�K ��=�G,�ڣ�P��N� �r��5�������s{ f�k�@?��x���9类|Ty���؍Q O!E�fL(��f�#g�S��*��_���M��[H;���
a@��6��ES�C��*�U�{|,��u�(&��͌Τ���ʙ�=���E�����@D�=G
#���2�e��~�^�V�Ӭ5�H��~/8���~�;��c�'�a�%��s@�������s���-б��!1�ock�RZl��d�.Y�h)F���� ����K�c�x��;�aPKod8�d���[S(6Ḅ�����I&�(�8
g���/���JD�-�q��iq4��D��4�߯��JO�����چ�g�j�'N��Y4�#h4z��/��W;.�z�T\<�i�,�B���I5�lO�tPd� �1��6���+�G�B��g]Ru�:'7)ϱeD�k�=�f�;c\+�-��dM��'��

����P�?��"`w��ں��M(Q��냊��'���tg��*=�;��BT��g����t���~P�Ф�yR�K�����`ǂ���NQ�6T�yh.�U?p���F8����2��EPn�S�����Pׇ��iIh>�,n�)�
���ߵ���8��?nH�;� _y�okXA���<E��zk/?�P?�j�O��=8FҠ�G���M}�����X�g'��OSg��f��iq�$��g���9cB��2��"��A�/� b�a�z���T`T��!�[�]���}��w|����\��1Y}|QU��;����1 ϕ���:�<�>��-ɡ�Hܤ���|e�����7&ݱ3#X6%�(�ay��Si�;q�3�]�����Q����`��
�3T"��|Q��Zn0ҪWu��T(���o����M[�p��c2W�o�~�"�̕x���1M�M>n��Gx�ܩ��-n���.'��2�M%��P#����;�Y��OY��%��fs�u�4-�E��ݽ���"������Y�&I�Ƿ�f�>+��+<(��ƎtØ�!`�$�t���is�.�iM~>X`����}�j��.0󡣈	#��n?T`K�ʑ�޿�ǆ]Q�8�6n���\�)���
h�~�J9"(CL�~�/$h�M���=I�S��R�$��*�L (ڏEJ~����:?�*.�S3s:� ��*�3�<Q����ة`1҆7�V��+H�Ѩ`.|��R:�o+7j}�d�}�	x��Ь�R��F�xkb!`�����] ����x�
��xH����2�3`��~��c�T�R�&�.4N"��P(���wmE���Z���oC��T������W
�|�DTOl01���@��Mʔ{jO<;�'�����@�ӧ�D�-x�R�aA����e�Ì�N�ٯM�Qx�4q#wN���_0�c��(��6$|c�wBP��S���MǱ6�/�����XNW>�S�CaRxʷ/)��ާ��>O�"�I����Ą��@8�+������pI�~H=?���q#$�a[OSiǋm���h@�d�M���~���|Ƙ�9S��@/��T�|~�X�=�DC���Az��+�X��ш���Z9Rs�ǈ3��ORZ{�I�T�\�Y8�*����|^����z.>�P�3N~Ҿë�d6��X;4@�O��z$��l�?JnBI�]��x�s�5x&��f]�
�Z���,|t�?�EԪ�q�k�wE�����TJzl6V�eG8/ŸS�tq�3"h��㌏��i{R~k2pX��6V"R>g3ܬՉ3��I*AՍ�%Trͭ[.�<1A+�2�-Bܠ�=[��n��?�����Yuu�̥�e&��sW����m|i�G� ��w	/ڕ��.�3�T2E�ڳ͑Y�o�<�I���r[�F��Ϙ��Q�Ky%LYA���x�C\���9���5��\��0)��f4"��RE��?�(��Iv��0Ws�A�4E�$~!�s�-����޳���$3����O�y��Ҙ�l΃�������r����6o9(6�d�߾��־"#��ܲvO_hKkb�����6[�[�5Jr5��r�o���^9��PF�fU�c�2�����0�<��m3&xgq�"�,���#:�)��,�W�ĐK�X��F�y��l�4���~u��U1w��<�S��+g��W(���_}�=+6��X�@���F�\&�tO&g*������lS��:�v�7�j"`���t�h�#�JƵ�Q�ѱ�w�����F��[R�1��'W�G�Ճ��>���I�d{�j�OK�Z��L��7]�X�|Uo�`ǔzP'��}/G� A�[�� ��e,#,{��l����ώ�CIR�"���*�jh�pN�6���ƘaP��9����C�L��Ϲ�-�����`�/J�=(5�{����L�c�$˔�U�aۋ+��u������ͧ�\\�i�n�Y]}��LDK���d�hRէ�O%�����1T�t��������dRfTcou����l0	Oյ<�u3����L5��I�0Y��c���=���*�kP$s�ca�Ĕ٢���Y�V�����(�+vo?n��&"j�߀���m��n{(�d�8����KM16,Sc��\v�YC�1�f���6�#�	����L��Q�P��@ɨq�ҴEo�Mٳx���cl�t�'&�v���ϝ�B)Qv�oG���|L����G��c� ��Ԓ����{��1"	d7�҇��<��m��ހ��k}g����'2=gTW�@u�KX�hfOT^�� 7z�F�vWa�����hv;���/��3﫾@�fA�c��|T�c�-�7���U������w�`�e0#xq>a;�>���֬>��4�4�Lp�̋\�+�q$�L��
�O�����u���vE5:��G�����p�'����1-��;0�*�o�����MF����,��=��i���r]mԡ �iY/�.�X�D,�d
k�����}3L?�p~���X����h��$�K6j��-�@�xw�b��!����x�Gh~��E�5iG}:��� ����.6��C?�R����@�(����d��lò,A`C����;�u?�su�Ʉ?Ӹ�6�@;g�gn�i�A��pi^���ԧw�Ǉ�Gh�v��K���I[����1_�"������( )23t�z
��;�p;sJ�sSG��	��k$tv�M<x�eA
~f:��:듪̱ �;>QB�ֿ�<+lȷU2��)/D-�}$�"��c��������e�ûnM5�SL؊��AtD��oD�?P�6����m&:�IEH��M�%&ֆ����0��	H�y���m�g�� Y�whe�p��JL�6tT90�pb&����Y���E����_E���Qt�_H�(IR�-
h=*����a�@�d�\�r��VD����lwS�s�}RDgc� �[�������v���3z[Ug���u�������~[���XPJ�rM>̫B���]֣ܡ{���8#2���ֆH_Mbp�ln��L�D	�Q&2]=�������`ոi�i�,���)&Z����Y�|���]���p��(?���,����?v�$	�j�F]�K��d��'���W����b)�gHxA�0��cx�;l��O���-�&��G�I�T[����\FQ�����4+_�/��ĩ�d��>R��S!����,� J��$�	�)���+b Hq�]vM�e!��Y��޸A�i����.J�x�ht�$0�V�M<��x)y�2uzE���[���-�u����Z��^7x�m:���Iz��q/Em�&�ɗ�hj`O��8��}k��䗘���nFK%�x�xɭ�{JK��v��)И��B�w�M�
,,�%Z�L6@_����	�?%�sG���.9*��|@ȓj�W���
�V�C9z- \��5�|����b���$���(9��=Nci�Y׬�خ��lU>��K��fe$�H��j�vcKIW��5�dU�(�O20=£(�=N���� ����V�-��K1���P���"��;�%�Y�⪰!��7G��nz�>��Sz;�B���s�g�%��҉�A�Ws�ɑx�$�5�4�؀w^�B8�+��{����J��q�Q6��0�G|�t����|\Y���p�bQ`v%Vޙ��Gmb���$V�k^���c,��w�9�B�y��U7����i�H��`-��fx<0�sN���O��H�#���6�~pJ�
��*wJ��8)h��.�PI����K�V�Kz��OG<�-��w�,>�J|�hk��𝷮�N��&�����f� .��+��%p<�_I�j7F�x��+��fF	��KK��#����û��[�v�v�?�o�ɍ�)@f�>��20�T��!�L�U����!�T�5q������\��z�@��e�'s꛿����6�{�8��qz�o���؎)�_$)��~5H st�%H��ƫ�gΌ^���C���1��g���U���*���2�޴2�p_FĞ���Z;y�1Ms������yD誨[�x��|m1%<�m��(
��K��C%L�%�}��Қ���n���q5���~�=���G%��
�.�� ·�K�w���~ZVkć 6M!���Ai�DYL�D�@N8��dMrT\����8�K�t&�GN��K�)��[�Y���L�>�WП�2��l�k8�a"S�9��M�e_"	CBZ�ƌ��Y�m�R�q�x/�V���7I�t��ѕ5
b_s�\�fP�4��d���J��`�uN)��\CH�a�~6�7�[�m[`S�U��9�ٚ�2��yU`�m)K���� ���gR�[1g���|=��&葢���c��[0�[RK}%5#M���4���ōL-�^j��-���b��L�귘d�'LMCؼ�=�����Y8!�)r;��Ydc��ٳ�	��j��I'��V� '짔����	h�i�Y���r2ӻ��bɊL�L>�:���J�$^g>ݼ��v�jFˢIK�^�	g*O��Ҟr�nC�jF�je˩��*,~(�5d�<r�B��V��b�ZVH��~���צ� u��j�`��������m�!e$v4�ľLݰ��݃�z����`�X�zg#���8\%��)���[�;9��b�GQ�F�9 �ބ��Ҕ脬_�.C�!h|W�6l+�wq�U�;��z�����ܲ�/�A����j�ٖ�Z)-mf������+�Yȳ��D�cob���+���7�s���+���"��Xx����¨S�#��3����b�iF�ҹN���,>w'q�Cܛ#��N�6�$�*�?�V�� n�)cg�9�P'�l��w��dW%̗F@��v���k װ��Ꞃ���B��'>��B	欫��^�}��,�g� ��,?��~i������C�3_��GNQ�4"U^�cD�������	�|��aڃL�+��C;� �2��Y����,]���=�����L���G�#�gpS��~90H��m���ݩ~��3�bV�bMp~n"�Bq �A���PPp���NC�\f�G��gf����r�o���>=�T�x���� m��_;:�v<�~4�F0�2}U�ǡ��D���t�I
�Ȱ5�wh�[6a����Z�U����W�B����CV9'駢?�Kݥ�����E����
�Hxe�Ԕ��@{v�Y�p��7�X=v�Ip8�t$2ce5�ŭ����7�0B���Ls$~3�e�ON��~���X�2�����@�ѱ�sq��JU�����7�x��}R���\�Q~엮��OT����m��xr�S����JB8��lՔWsSW���� q�9��2�1��eq�Dn���Կ���!�r��,)�r�'����=ٖB��T=�ؓ<&�d�L� 7OI�������*�NY@���A�$����$Q�kH0k�v+?�;�0v7X�P����Y5��A32���6��W)m�ce8��x��Jn��=n��w����|n `׀G����EW	�n܎�%ϖP� z% �srp]��{�;��O��y�7W�</��}0w�AVXv����H7� w-��w�z�O˅���l�=0�=[�1�i����2�M�'�4��:b�y �=��DVT6,2Yv�R�����,M�����3��Y���F)4���Y�ӺL'�o&I�o�[�X���9����٣�u���k/(�D�
��lޭ���=Z�nHۿ�%�.h�\��4�01@暔����@,��]��_��f��������J_��d^QY�1�Ј�L��K����!U��[�	��2 �MG(R���~�n���d�IM^�z����Q���1|iA?<c���M����}C���A�>�I�+��h)�"���!!�(�m_�.ui73:��]
�p���,ؓ��?��.���!��A���䗇����w�[1�ݶ��C���6�t.�B��ۥ�'�G|���%��j�j�U>�rJ�����~���ze�%�Ǹ�Al�*�F�D�!@UF�D��/��VI�)[��ލ�ƈ� �
�\��HW4�,1�ٹ���n�$��ϙj2B�#�4%�J���䈹����uW����ϻ/��/���۞OV����_ّ�_9;Ok>�l|������Y�ݽ��<�����a$�"����fn�%1+����|�n�7��|�O���ˢ���G�xHG��������y2�%a9����n�}$8�p7یP/k�yZV���'�5�Ǩ=#x�k[���'��yU�s���%1���fC��b�7�:u�l:�ƛD0�L��E)	e7��H�wv�����:(%T�t��v����X	IV��qf�SdM���-��1_�}�2&�J�x28a��^��1���zs4T�b�~�V�_1l��*�@�!�*�=*���PJ�?P|i>��K@�n#:"`(X�薶ݟ�nX�ѩ�^��J���؛`o̲E�6&e��V�Y�r��w�������G� vWG�Lc�v����=�G�J�҂��1&5Bnǒ_j�)/�K.9^�=�^��ߔv��;_H���'�Wrj��e�DChy$:��Ո���j [�Z~_�m^4C&����.��o�-��Uo�3�����<i:�S�=�p���9�����1d [�"�����+����[�������g��Be��N�뵒f!�ʩ���hM,�8S�aЖL��@}�u*F^?T��@,�O�hȃ�$� �	jQ���+:�[e� 'I~ķIc�Ls�-8��p@�~'����g���o~�7n��@��8ƕ�h�P�~��Jr;�/�F� �t��k8��iy�ߘ����d�f�m��'���Mg�=I�Q��M�0t��2�K�U#V�µ����Y+Cr� z�r�j@ػ%l$�Z������*cR
�"�_��E�B��X��e�U����~��E&) E6@�F�Ư�뗴�0� ���>Q�V{�R��(^2�"��r�����7F��5���v���ѥ�b�����5��2Q�W��k��b��s|瘤���}�u�7� �=ٍ���z����VK=;���ߟ� V����P�z���Hz|�*�fH����rni�F�w�u�w^�{�w��;��%p�GvE'#qOY�	�1�e�dr�>A�/��$_!L%t�7��~�7���.e��#Z&�ނ�P���7��6`K���~r�oE�n}M����+�+�bz�_dƇ)��-K��� ���h*8���Q��l��8�;�G�i��*0����|����X���4�S�\b��L�� �;�B�l4_$<j���b�Dg	��O��Ρm�	?p�.յ1�)�qr�h�������|�ei8�i)�:9L�/a\�ܜ�^z�{��ދ��R�,:ݳ_s5��
�
��z��At�e<����J,<��SykT6��*����/O��M 6�$�h�r����.�l��]q�ۑzs�p�~v�D�������Պ���G/�Lc�6%��p�Y��*�9���/=A'Z���l��x[��B뜓z�?���pB5�e�Ѹ���c�м�4���J,e@�'k֖��`��>�c�s�f�`�䛍��c�рYT��)�|��eE�Q�?�$�
oM���=kPkR|r��p��h0�v�B5N����쪇6�-Q��'�[�mq�lB&ڒJ��վ���Y�g�m�TkK��_��F;�1$�>�r)����C�q�Œ}���O,�����W��g[T7b[:�;�wB�.��L���@��,����7Y�A�z$P7�ed�隿Ѩm}۳]�>.��,��0��p6���%���硶"K4����l]"���1���ˌ�]c⦆�Lƒ8�;C��٨l�q�t�MK�ټs<�sF&���%��ު�h�j�4v����3������� Pc���D�o�Lf&�`�����hA+�RE�vSQl����k��.م�z[���
�i�
�t�����F)�V��7:���!��R�~s��qq�O$�C���p������-E=�;b�����v�E���\�J���$�lF\ԉ$�f��p��Q�O�vT[/��
r]I�����@sHp��ʶ�u�,���������m!LaJ,�	�i�w4��E�8�q�-���^'������R����r������Ӳ6�	9�8`�l[���E���mX�<as~�t
�HE��ͧ��d"�b��FNй@Q�i¯9c��iU���f��U��}~���>,��������KXO����EB�P9���!F�D.���O�e��ō��L�H*(3��"��R�W�V�ʶj������H=H�3\J�̐��AZ�AE��O��]uq_�@��nh�0V��w�(� [y��������ݲ�#��f��fX\쩚wc��$�5֧
�N�}��v��i���J�ۈb�!��v��cI�e�A��=?x������g3kɮ�d@Q�Ph*Z�zJ�HP�Y%:S=��f�`�(m�#Ѝ�z0�$e�a�hM�6�{.��6��b~F.�y���N�y�q��g1$U�y����W�89�5�GS�.<��1�utv����6OSj�%�N���[v^�$�����[
_O�Gj��5�4�(��*m�'����Kɮg�R/��fѸF4��Ѥ��@��;�u�~���r�z���@+��HB�2��t��}�T���SF7�!���Y��l���X�3;�l��ry�{o�D�������˴�@��E���3J5��lO��?Ǳo�Ip�V��(?��𥏏��]>��� �XɎC�4��3'q_�E��E���fQ�J��nO^�����-z2W��\���¿D��Ȧ�2��Fh�����V۽L�"`���%�8���آᔰM����0�+�E��lR��%d�9Q���qX���B�pC�^���^-�5L�ܵ�H;�o�*�@'��&�[kW֕�P���D|Y�\^[��(#��q=�� q�_<4l!��8xۻ$;ˋ̛���6�@���s��t�U/�"�NH�:/:\s�Mz2�+�>�V��ңcKaRz%� �i�وL�.]�[!�l���uH���-��/jp�B�|
b�'W����������y��3&��ZE��l���^�c�oi3��֮0�r�S�Q)8���LZ%��pLF�ü���k��S�,��7�"�i��Pj`�'MI2��#]�߈�^�4/M^�-�eA]ߋ�3��}N�a�I�A�h�����B�共���s�H@�E���w�����1W�����C �x0 %"�;>�\w��W���>�'���W�!�5�W7�j��u#�E_5��m�M�D(Xح[Z������H]�acו<���yj~�ƒ�h�Ȏ��"B�b�ٵ-nm�����;�e�"��s��!��~[��2>T������q}���7L˽�PϞ����rU�c���虜�����8d�Q��4߰N��etVȨ,��$ul����V5s�~�mR�3P�j��)"[0;T�S���B�Ӿ�~Ҵ�@|E��()�߭�:𹀷���5�XU����8�cl3�J�C�܃(���kB���� �7Y��stҬ���"����Uɜ�7��=V�Б�^m�ߞ�`���b���7��꽹#⑝��c�P��b��fx��ME<|��!D�Up@�E��x�\�ӊ�ZN��ga�d��'�	��U�'�\��M��͊!j�q���I��}��b�����QXJ��q]r�+w���߮����	@Lk%~O~�V:jr���R��HG�ʘfጀg��$Zw�R��ӯh|v�!T{x<64�1� �{6h�LJ6�1�*O"4���*P�(=��	���G��(p���^̩�+x]��Z�-� �Gv��Gg����F�i����ɊJ���������A��իz<s��A_�<����1��s�1��¡s;7[P�7�.^�]!rؔ�f�s���i�j��V���M<��+�t_J�*�a�j���B��2���n1��Q�����L-�l�0\B1��&����WIa'�J`�5�[��m`?:�-�u��>Sg��l��[��)�1��a(f;�)m1�g
�p:K�c�ڐ��X���z�I����#�ϐ��4�#�J=�G=e���+bk�7����Hn�܈�#�$�Ǚ=*W�]�@�\��V=�Ӂ,B���͌�Gjm�$�N������RL��Qqr�E��o�#g��]�g�_� :��QB��a&CR�V���ǳ��/�j^� ޙ��$�iU�qƙCuT¼s�j�w��� ����Ѳ-�ҭ�(�7H
�
�D�6�heq����S�8�I�P��UQ���.}�p�3�.re��`�6�hZ����b��P{��́�rS�\��wyŌ��$<��Ȼ���˄�ir�cBeMBwW���K�XvtZ[��(Wޅ�+~�5ux��#aYbI��6!�^�ͦ�ʯ#_Q��U��sQ�UgT�EQա�8Ȕ�4{�
���N��Kz��M��<+�9�b��lF�C �ņ���Ѝ�@%J_`>G�G�ːҾ2Qnf˲�;=@�E`Y'�L�.�+ӭ��ڥ0��Ab<��{x��ܹ_ނ����*�R�{�D��:Vm���G_g�b�F�[�|N���h�H���@~�ڟ!O�&�B���פ�	�@Q���?�E�! �c+�FO���)�wzA3ͨM��d��4.�f�[�Xl���iU<�?)�Z]>�,�Q���Ygyz�X7w"���,�
�He=��3-@q�� �|��v���a�6w=~5��!c����ɺϹb��q�Y6�Z'�Ճ��I�W��xz�G~�6��V�͖�=S&�[g��VA�5�n9z�KaJ��J�UŠ����xD���U��뤷�%
�Df�'"@QnP�d"��-�D���Ԃ�[s/���R�q��JTsn�!�_��1ЍG1�j��FN���f�Z���w�|8��z�60��n�cRjK�'�e6M-՗+����$�.�_�*.Hc:B�����NC��
J�������8��ǖ��JK53gB(�O"�E"��O<�WHS{����������E��r�Fm�t7'���ZI�w��y��S�T�Ru��!����x��N!<���3m�!儒�������=N��q���ܵ�G���~��n���u�� 9
#�P�f���`���S��!Q\��#�7�lu���0ѫ��M���Qx��+7I�����9���/��F��Ld3���`A���c�$˹�W�.*J�q��]���T?�"t�s+�������[œ�[}�}�r�#W� ���Iѻf=P�Kӕ�ʕբ��v^�2,����s�vX'f�8����&�u6�h���)�k����W��z�G�\C�輺�z�K0���!M��<�㱠!uY!d�%մ�'�s��+6�_%�Ȃk����O��g'a|N��|0fGS�v�m�:�"ajFv+m3w�^�|�@���cl�^�h���L 6�D�#��G{$�����s���R�u�6)f���t3'/�8�=�XW�[^�i(�`�F`S9�J	f��׈��E�}��H��E���T4x4h������tٓ���e�$N2.����,7��D�;" �
"� :�۽�&Y�d�[ї�,O��++KY��Sd�&�16LW|�B).�Otf��+���>1�@ˊǖ����]lQ�&���$g�R5}�f�g��z~���Y� � x�KH�j��{W<�a�
lEYYI�n��㸗�-�(�`c��W�:��u��[ۿ�a&#�M���,���i�Z*֫_�����!����_XC�n+�ڎ�V��E<�Ҧ���G�d�w>����
���u�� ��G�*�$w�v]#E5����%D�-�7�+M��giZ�������&#*_<ѐ=��c9�fb���)��i�����،GE(t�9jnW�3�rR�T�{u5����o�����ɳt{����ft¾��NƗ-�i쇥�)���K%Z-ז��<��3�`o)�"�p:��FSL6�<�f2�F3X*^�d��+Z�o�Zj��s&�tL�7�mAm��qqr�i0z�f�����-1(\���nc���:s%>A�dA����L�͢V���z�;OI�ԚKe�YcQ~e~o�O��͎�\f����pb�������N����
�}�*\��}&O���ºN�.��T�&FQ�h�O�~�qݸ5r-�: _���f߹��_�.��!�h
�_,�h�('>�c��t#�*����-�uh��w慲�zj�*�!\���� *�7�8-���"z�)>y�&�
���t`l��ŭxR����<'��-��y�&Yv����/���e��l���{�l&q�Zn��z�	������4���m��F|xâ@��a�LʮX[��&��#㙈�[�2�C�j�������6nY3]��0|'�w���`�֣&��/,�u��Q�����PR��XRh��&��t���U��}ً�ޓ9:�UB�C�t��'v}
X!=���J٦Rc4vG�,�r8[� %�Z_��X�/'P�ɋt*�ʵ��t�1QNE�[Ш�΍R)�dN� 	�}����l��%r��
[��v8����mD0� a�$юn�2��Oe������nYVHKY��R��gM��%@(U��V�ğ���,�D{�O	ʄ���h��mb����zy��;ee	Sn����ޠ�35aѰ񂾌��ަ����-$x�+D�����Τ+AI���'xAƑ�,�N���S�kᄬ��c�P��4ځ���G�g(�R�:��������p�2�-ϩ����d&�a~��S@SY�	M��s����ܺ�n-��'�@n� a!��<�gQ�]���%me1s��z��C�sK��4?����wY��w����B�c�T�vz����(�|���X�,��,�1H�1��=�;Q3d�eL�e��ڲdծ,7�ٕ�4߳Cw�T��p��ΛVM`����x�*lW�W��@���8 ��[2���P����=�vc�Z��Y�C�)�N�U���]�������tnA�>�����O�[�It���
޵ny���)�Z������M%��N�*"Y�}������w����۶h]�WB��@�0��4��:��ѺGf�JSk`�9�3��N��3ևv��{�ش�B�Z��ᱞ1�؍c�2�3�k-�1���� ��ީ.Y�<�@��VP:7�}l���z�0��
\�Ȓ��n�i�
�LV�jL���K��o�P܎XuТƢ?���	/:F�Ǌ����>Ĕd���1!�L���7�M[j��>���Y��̑����i�lއ胗ui���m}��Nᴧ������g}�YҚJ�ͧ���i�Aev+;A\Z�-p�x���s̼��2`S�O�uM{J���(Weg�1o;�/�:/�����K<Mұ��?�����C��
���!�Z��X@����(D��o]��\�R,�dr���"9�*�K��Բ�.#���hG�b�2�0�xz���]��;b��p6���A�k�3{_�Ư��gqDW'`ZI����(��[I�&J�!�5/̂�&d�{`�ʤ�'��8��z�ʑx�o`D�nB���[:�>���Y���gý�Z
��z��>��wIZ
�L�
�AC���ܝ76ś���RK�M+�yY�/ڂe��5|��`~GĞL��wm�ܼݯ!��Ĥ���ٝRl��َα���R[�t�h��l�\k)r:گ>�:V/�{WbPUz�	������@�YAI Hi0���*����A�^�PH@W��'գi�ӈ��76S�{��n����9Վ���d\�����_(����ђ�i��V�DL<�i�M�UA�}�2�}6�_ˌߙ���^F<ײ=�]�M��}ʑb�F��:������C6������E��"
[$ɪz�6�HO�zE�	N��`���jW�%D�+���f��`���9���<��n��@�f������&o`X�I�
��kѣܰs/D�ϱQ��N�]�/+�e�>4Ni��m&�AT=Փ�p��@�Q��;7ݣGJ��bO˨}�j�8Zv�u�/\���O[��j�`�Q�bb��&���7$�6�Cws�k��N4~(��"���l0���2I�ul1�z�o a�@k���B��#�6AUq�i����.�
�����E�:�|е�?0�$�`�����%���7�0DA�D�+�� �KE纣dێ�ɬ�Y��Q�N �w�F�&�NI|T�A ����D �3��]��H�����.
��U��b|�(p�/<�?	z�S���\,1�V�b�E<%o4�-��J����=�2\i�f�U��O��)��XW�!D���J��>�*�cI��-��i�6����o�����d���������ر�u���@�IO�0�]2\��o���
W��od0� ��ha�\�k���	���n5��B]�.�f�x��tNl �'�|�C�"y����O�G��HѬ3Xf`pY{�U�AF�\ՍE���ذ��pp��(�o5��P[a����4P��}�)����_��s�m0cK��M����W�^T@6dS���P�̋�2o��;Kz,E�����u�\[�m}��%���͙����j�0j&�	Kc2�&9�E��y]qB�I!��U[̱�6�	�\�ۊ2�G2akr+y��L�(��xY�6e����#�s��1����욗��%��o�-�M�Q<����P��(.��+^�$%�ÌS�[e�o t����{e�oq���߈�u��cϝc�w�e"������S�E�a2�i�FB��3�])g5��~��kO$�&��AmpC���ӻY�dK)�k�9�&"V w2���z���L�"Ba�!4�lK'AQ�Y_�L��o��v����<Q�T�Ǧ��./P����~����r��!P��09%|��@W3�ڸ�CY�T�a�A���V�!g�u��W�HZ��C����Vb�	'q6y�=��ح����($XΨ ϛ�_���'�飦T�ِd��X��y���� ]�F�V:�uQ�dؠ��	���<*2(Sbx�sjjn�o@`K($�؆f�SSd�� ^q�Ю���� g��𭜑��>�M��m��hj*�U����W	�5�`V˭��p��j�bg��\X�2� �)���Ag'd\�V�@j�D���4pA�C:Q���/-�4h3�^T'��D�1y5q��h�&�?һ���oz�bq'Z��D�ԇE䶯��0����BVyi".�߀]�^�䐿�C����c`!�������~]$�ȧ�#�C�(d�?���BD�r`=q����DZ����LW,�&��#ǎa�r���o��*xT[1��cχ+F.3{���A�"���{s�x�|�l�]յ���o��}��Uw y(^IYo�� ˪|��_�At����0��~�
>�/�[�X3�R5ٻ��9��-*�O�;��u7G�7e�;��ŷ�*��}0�D��xS���g�����V)�:.#�l[K-��c� �{#�/ A"���]�Q�\�_U����Ǵ�\y ��B¸�_����m��m@��Q�C��4�q��~�A���t�Y�>d�`	"P�K��ŕi@ñ��'<bз�@�����N���薳�g	*wN� ow��Hҁs�^ӕ��P�4���Q5/������|���O&E+n��k(2�?2�����MUyE{�odu`��|v�R�3X�!�8��������v�T���i%W�W���X���
��ԙ�.Q�Y����,=�:�;�����B�G+y�ܚR��5�=��K��9���1HC�˵R ��J �vV�X�(�,M`��a(�,�"pl��\҈�'�6�$pI4�S�#��Х��;�H�g�'�N*M�&������1v����(�miQ�����C�_�:�j�G%x���۪,e�4 �~K��|̨V�ݭ�pw���i����k����Xw.���#{��2 
ˉ]���2[�6�;��K�Ahh�|)v�F�U���EN^�)//[�I?'
�K�xP���vxf��bg����}�[_�c]'I���IrW��������[H���8Ce��ߠ^Q�m
]�ʑ�!P��d����dD+J3ػ6�%=��bg�cw�Ŧ��u���Jb�nS�)e�C��/�Uo	Q�2 a��e���F��z�yn!�2'���&'��Ұ����Db���va�7��+���9*��I�K| 5��v �4�(��A��,P�:1�G
S�:�f<��1ohC;��XYė��k�6W���M�_ݴ�2x�����~ݓp�����m�������0�d��Ef9�J"�',=j7��}���I�����j��mi��cp����`�l�iv3���pK8���8f:��D��T'o�!3N��h��c���d	MI.�ZOm-s��مz�
w�w$��9Ʀ8
_��]؟|.������������ ��9�{�	�F�ϲ	���6���.$S����;5���0&�o��l�>Z�_���ݎ�-�i�!"��������Zq����gm{�[�+]�Р�%C�}L��M�mh��N�Ϣt����Ak�$Ιg�͖�W��0@>��=kb��7�O�"�Ȅ=���>�H�N%���Ŭ
M���۝R�5��t9��
�02_Em�A�!�1-
p�kf���5p�y�����U<B��r����<B ]��ߖ;Л���q�$�F$���nO��J��ۛ���k(���D�=U�`0g\!��z��w0����w���hX����>h�V�}��z5f��-�S����H���=J�L:�P�+R�=��i�WR8�� �|���Z��˘�G7���������/�=Ma΂W�9����I�x��f]���8|{!?�
��Z�n
���x~���v�Vm�F'.�S��ϑGqAHu�����<���U�m�YZZ]���H��؄�p��.W��d�0���fn��ԡ����>c�����F�1}��z,U�cdS��C��f�q�&��fVR����`�a������m�VS5�P������s�YH^nяV��܈%o���[�Q=�X�R�c��I��r�J��Yd�s��&]wt��Q�!�Cz�5Y��Ph
؍~��~�)���\ta��s��&�6�Rύ�fPMy�c^$���6f�U*�U�QU�U�/��IO~lD\A����1��d$�>�ɓ�$N�j��ȱ8�R��{VL[9�.Y�.�0�M�:������s�R����n�
��K� U��bt,-�6d"����ϪahS����M�>x76�@�����h[ޢ&�JZ����^vN���g3i+{�Di���J?%�v�ǟ�p�"��j��+��&g��_���2l@D��A�М����o/��om52@����|�7([D{4�`���r?�����2�H�x�gu����%���-�/�%ؕ� ��������7C/��h��9�g���k���4E�� T �$l5��z�OpT����1���6<�n$�+��Z`;��k�,$Mq�尗�$����}�	粼r�o�����n����Y�P�>Z&�,9,�`s��^혿���z�~Kf���Ѷc� �O%jo.��"pmpU!�z�ǖ�  �mh{��6l��7</q�	tI'�������0Q��<P2��Q�Q숪rz��J��Wc�.*0<�i]Gs2g� �����ϛN�ڑ�%�Lq~�V̂oC;���I=;�!*j�xCbS枼G�0�o��Í��j"�^���t��$c�$b������Ӥm:�qm�J�0���G��^�ht�f3(��<�P@�����6�ԏ�x�ܘ^���� )�����*3�#@���P��:����/����W0U��3�_p�t�d����F �=������0,l�Z�n)���Nn�]	����s�������w���=��=.H*2�ƚ����hu�����"ĺ�~_Ld4��� ���'��	������#b���|�۫�*�tIaX������edd��PU9w
!8�Ѳx*Y\K������✪--�E�Եi��F�JU~��`[��1��E��xύ�0�8�k���8ҳL���aKA�R�"��OCs��4/��Ͽ��8��MF�J�ok�mby�8�P�_E`�����vk,3O}���k̲;�����?��돩���#ݠ��D���v�}��i�SB���"�!4,��^�z�n"��ۯ�i�;�ɛ6�q .O�٘l��:x2������T�5L��k�EM����Қ�����2�;umϷ��5A�L����3^�/e�JEv������:wBX�O�7�)+�֬B�._6#�'��)��5o�KH���"M�ZM��9�x�H\nt���J�0x$�aY�=�:H�U�<�8`pS�����iF�y��Q[l��W�5T��im�� 9 kC�Yh�u4�"�o{��ϵ~��!�����M�v�AڭFK8h�c��#�9$g�E4x�­ɂ)A�!�8��Ϭ3\��j�"�3���,OB�-�o���>� 2)��vM�?��JH����c��e��Ӯ���'�Yv����D�5½)�ޜ�L�A�,�=�k��#�;��G��3q��j�����ϻ�p"w�{���v�m�OG��Cʯ"v��Q�q��ՔzZ�����a}rNѓx���eL�%�ϒ�
���-5	9d2U�p�pS����K�'}:�U�%�%�1��U��ZTM!�+>��:�nh��t�O':��&��/������J��V.�(����y�6GLO��U��p�r��q�F�������/�+T�^�v��r��i�'Z��X[$�� �]H��������VD�6c�lK�!�|�,`g8!B��-���8ǣ�ۑ2ŕCH�u6�w���J1<#]M�lu������� �wG�C�J9ȑH�O�h����7j����y��&��i����'������N)�ż ��Vp�|��RMQB�w�6Qd>��pؠxww�o�o����>w�>s�s �Uѫ�ľ���u���z�2W�e�)j���9#[U�<v@.'K�73����Ǭ+��69����h�鈦ւ�����<G> P5��Ԃ���ԝ�$䢓� TJh���
n�����;:�Es�"ܪG��E2�V/0CY�{����`�E������#6͚���T�ǧ�{s2eL��l=��a"�Bv�2#�y�&tʙB�����4��٤����N��N�D3b�����Ԕ�%~�*���i5K�K!Yɇ$�� �U�ܺ1R}�$i)�:���V훩U�T�C��7����Q��>�a��?���(�0�A�}���8ͭ&���~p5�`��|��t�b�܁����3{J�\�[8b��W84����
3[6�h�W0�������cG�,���&[v~:l�L;R"wp�&'&�A��&�P7F�zq$W)�k,&���T���f3WN�'����Z8���^J�FM��zϜ�T]�� ����=s�����.�ϔ�i�2��at�	���V���Bz����3�,/�Xނ�Uj��?�ڙ
&E��۹�^jy��0S:ȣ<ٯ��q���@��'�ٺ_��|WM(�vm�3�d�<�%���|t�jA�IL��8�Gɴ�/����bW�w�eݤjƻ�ʮ�+dz��JS�gTR����sڣz}�Y�j����+on��ʫbkXؖ��=�|_%ʮ+��D�>ޢ�q�y�R[���ad��g`^�r7^����#��b��[xc��A�>�����sQ��T��֡ؿ�e�[=��=�1�4�`�f��o�H��1dgtP��ɧN�;�������yA%R��jJ{�U�	\�	�h�m��#���`���!���g���_����I-�V�y������%>z���9'�yfN)�rfO�CJ'gΒ�-���)m+^8t�#�Vm�A��k݆}�_d�\j@�{8��x �;l?�lB�T��rW�z�j���˪�qneR�gɖ܂���OHD�S`��V�wX�+2f�ui8q��i��8(7� ���יB��I[2�4�Y�$����4d�Sx�,������_���7g���i�`[��d�|�?+>]�*���)��x�mð��<d-�襷�nH2��|��q�B�b�]^I}y_u�}�ع�^m�5=%�=���f�=q#Q���v�g�n9��,�>m�����X5M�M�Sbs]��n��W���𴨖�Hd�a�Ɏ�;�^m�&Ga"�i��g�S��;��^2��L�h�t��k�X5sE�u���������>Dؾw���d���'�t��^x�-駜S5���4�ɖB�r
F���}��1�v�fd@;q
"�1����� l�Ý6|[>�i�9Ȩr��zHN�<��_fn$M�-ׂ .���]'��7 �EZO%s���	d�ɦX�?�@�=���9�lީ
�����4�[K#�T,I�gt�.�E6�q�\v�@�X>�^7���f����a,�1��Iw��n]��¥H-����Ys^1�k��Б�?N���c�wބ���̡��p�6��?�G2_�&R���e ��x�T�"�'��O7W<h؆zx���W�u��H2�-P��p�Q�ѱi�WUw��:�.�熃�}ӘX��*dy���dW���v�5�eI���)�{ ?�La�oɶH��C���yu{Z��Йݽr)5f8���~U/��vxk+�5�-B��]�;Nۺ�_T?����2[ ^�.�"I��(w�����w���X���~*�Pf{yVO���5j�g 2.A7v�u
�Q��Ɠ�,c�?�B�Bk8w�MKA�$@mF�-�U~:g+�ګjp��f�o`C�J����3e7�h�:Fͮ��[ta���E�Ħ�%?�_�r���ŷ���[$�;��%ߡ]��j:�!�X��h��pB�g�&zfcAx�k�qH?��G������x�[Iܪ �(r��2��]���6إ�%e�N�p���ie�d0r��N��$�nc��x9T4��s�y��z
�*��GN�&fӦ�|����-��$�Ȓ�xܱ�[�0K��*V��{2Z>�?�^�Q_�g���× ��e��VlIQl�'y{x"�Ӿt�m������f�?��K��3
���4���X��6�K�~�%*���P��.����>�ʘ���nIH�X�S0]�y�Ŭ z��Py�k ��c��;���r7��;$ڪvi�Q�px�|� �M?�5�;�mҺj������+��	�r����*j���W�MmxMe�U�C:��������9�Ʋf�Bc|8��q�E����:xqO�!1�sQ��A�m ]�,b�޺ sW�d��u�6דbI���	F�G�e\�� A�Y�5Ɗ�]�r�[�RP�mh��%���1�f���G1 ��Ko~�K��*�b��馩�~*~�ǵe�$����I���b�t(Q���=В�<qGQP%�y;m̾�m�����'"'�s3����ÂV��t �X����7�g��E�1-�Ӭۭ�N�sQ��&�k"���bTw�5����B�R��338�tf �{R|Ř��.j���^�]lfg���!�zp*is��;�b7������ �	��U$�zz�0!;�\�J�J�u��� +��Ԅˡx2�8s�0�D�_k ��)��5ҏ��ҙ7-��\��i4���d��r�R.*��oY��\��(Us{�d5��zC'�-�����oalk9��iN���l7e��Q�bp8�^M�!z��ݪ�H�z&K���V�W�I�� �Ɛ�D�z;,B����7�K��H4�mrp.j��gHv`�����Kʙo�(UL�V1�O
���+�;��l9��xӌ�*�n�0_}VI���`YP����<+}3a�A�c���!
��y�=�`���i4X$���')4�"9���y��R��.��vtD:^��]y����Zs���t��0�=��;�JF�zX�5�Al��%���f&/�6��Yӣ��f^��`;�Qy��,]�i�9ϳ��N��(��/us�i��R܊�@���߭
����bN��};��|�ž�J>�r��<Ͻ���:����������Q,�!�-/҆8�q���9����xw�r�ɜ����+;�`\�2w���MT�*ۡ��/��¯]�4+<�x�~�@�wT�K����K���f�sP��L�0#�${����"���F�N��U�5n�81����Ͱ���<х߄��M�>�k���̠�s9Y��u���ӕ�gm�����Z7�f�\�!F[� ���t!���
Io�~��{ɥ���4ڦP��1\���&d���6��a�}hvy)�1������ف�B�S�g�4��0��6X~����f=Q�Gi��o�p��H�$
�ߤ�i�P�i�Oy��S�G�Em%d��^G4�x$�s&&�w�4f��{9B4]�Z��%���s~E�Se�ó&��!9j6�~�^\ g�M��VCu�%`<Q` ����� 8�z�t�Yz$�3!�0`�I`��wZ��פ����XL/�G��{�5��x����s8��b���@~�؅�Z8���U!;�U3�߀ M�ݔ 	��@�k�J��ң,�F޴g����+�{5�C-V�h�b��-�u-�>�����R�߯;Nv�����q}n�3��ީ�^��=�Ḇ^&��[\Z���D�Z��JJ���f���3lH��P�fU�Ipz��_��Lo�t������0���Ӂ���@��k��Ub�v�	;Yjn˻� �K�4b��Ҏ� �R��}��s"M{��%P��MCq���i}'��r��K^=|1.���d~��
�lamC�����3�o�fA7�k�癇���t�np�w�4��}w�=^��4.��7����7�ز�/��(?�p�f<�i����v@U�(՞�����n�\�zZ���.�*FNI^?S��"893���R����Wb��u�*�gGH]�4����M�3��f��\q�v�
.��f��~j�B�(ZE ���%����g�2EUB02!�f�?� ��%0���ΠJ+���bt���%K�EM��xN�]�E�R�+z���
/d�n���� ϚfTCp�H%a�y�c�c�T�0������X���P�?�	��7^J���g�E��t�w���8��_.�o+�T C�r���J�b�^e�������#1�j��K�o�yY��=�Q��h{�&����Ԛ�pR�5�ić�a���y�H�>�f�,��x���j�@[��a5T�=�+tr�E�̣ÑG�n�nۥäk\�Fs3�<���:L���0�Xd#2}��A �\=�7��O�sU�5�1��iX4�jy��lZS��k��,�:i��u�\z5-;�2)}�-�#�L 1�wG�==nX�J;��_	�zҨZ��M��o�b�fO�2s��##H�V�U�%d��M�e7r�Im��J
ar�m�����v�~ Y� �J�^��쳫whtK@5�K��l����R�������Ca�>�MͨkF��B�?SH�JiQa3�S��Z������F���S���A�I�1�l���-N@6�F���� ���}a��j�$%��u�s��0Q�>�챀��%���U]u��	:���<��G)����'���@l���7���֠k�`�͔؊!Q��6�����������"i��;��!%q��3Y�ޮ���Ǡj&-
\�}�L��Ղ���R;5�a��ԿB�HO����д�[��᳢�{i��Mv�^�BB|�C�@Y��*�+��hڱӌ�s���{�	V����������Ad���swh�& ��`'�b~�V��p7�4��s%����SlC�(���M{j��v<�v��!�Է��:��Y�$��'E�C(;(��x�B�6��;��XqB��0��h^�-�l3D��9J9ȫrjds�vYj?<Y�-��#�F$-�G��Ft�τ�٦��qf�ބ�8��� �u���a�c��sڮ  )��
`Y 7Aҧ��B@!,~�kz��I���J�G���[���i�'�eϜ*9��]E�N�$�y�-�큶���,����i�&A����7X����MU��rB�2m/�n���G�I?)�������s) �����OH�lovE�w`E�ԇFÉ��M����Kc7��XH�����P��a��(�~�V�v9�[�A��Q��.��U\�^����Hb4aov̴���7�$c�2S�x�|�x��3��-�J&�kd����r�WϩB�q���$~�!Hsy[��7������\�sY��Y�L�;&�z�`��w����|�b�;��<��V���I���*:B��Y�0�7k�����/J�_ ϳc*��N|�l�H�A
Si7�]�y�=N��M	Jr�v�h,uw`��vr�,m�Q��:%�B	�f�o�~8�tu��v�4l˒���H&�0���kJ�� qpw��� �5|u����,m69F�* iAJұ��O��zH��4a�����0�E���q�NF�6�}�5Pփ� ���L�Q�轵DTsIN�Ԫ�=Գe�~��o��-�Zq���3�Q�����5*u��~�/��щc�o��qmOc9/di��r��������B���V]�(9B���cU�Qq2sȊ�KLlli#�<@�]A�Τ*�P��
ٞoaA�M�����[JVєO���!�V�5�쩴�I���R2HN�	�\�o��Ԡ4����F�@;B*F�-�d���z�e(���(ı(r񮋺�H�ͅfE��2���e�9��i�X��4N����v� �M��f�b���n��Z�\��Pl1�G��/o�P=<�1oI}���-�;[#`-�O�?�6�H�m��갶A�'7U�	�1S=ʱ=��%Ԭ�x�������J����$����QE�ǳ��`���>^���M�h��R�p7�p���A��V��dܳ��BT�%�#V��u׆fd��Q��:��W&8�'j:��k,�zĦ��i�͝�R�)QQ9 �kt�B/�o�Z�4�NǧV�*��Uv�y�Ff_p����:�ꕺ��j�>?�V���<]�T"��~��������7��l��1"�Hsߙ�٢c6+mV�0n#��7-���"J�����o��aMf�p$9,��56^���}X��"����ч�g7�x:�Ի�A �R�K&,����y�z)B5��^K-:��AB]�<6H/���đ8��ZlQp ٫pэx.<�*����� �1��)�C�L�Î=ߚ$ϴX�bM<�B���؞d���x+Nt�P�k;6P��[�vj�~��Y�ͧZ��Z� ���$o���=A����I����XT�?�6 �F�&���p�+z�k��@��G�u?�G��8�ռ�t:�f�\�x��:����t���!���P�*C��uE���aZ'Ed��7XC8�Oi�2��,6���RaG��2�Ct������n�p�E��t���S5��^X�J3��sdGFK���`)KM<>�Ԯ+.7]l�xS4�5-��U�Oo��J���K$�Lf�8�����(�br�~7�9Ane�qlTV��	�� �:�(A$`K}(/Tp��q}�7k��&�qӇ/���r������Z7�����d���沨x>�������uZ�����x�8auej|�$P�j�W�L���t�.��N�|cK��])5)ɷ���m��L4�<��1YP֟`9�� �j7V�u:�8�* �s��y16X.>���nuɃ����	�Zu��y��ze�C��5V�
��}�0�k)�č���g�9T��0!#<��7��@�_�@�R3�{��v��a��h�f�%�;ġr�3j�sl��G�}�`3e�~�`�1���w_�:���.�2�'z���d����IXu�w��'������m�DW��쫏hV-�"GN����yp����b��nl�h���r쿒�Z@M��v��L��p�	�6pU�vH)�6�Fyh�ϣ�Kn���dD�K��5N���T� ��F&1K���� U��ښ����'�cD�m
�����j@�Ba~fX�E:�������A��_�̋Z��\�����H�:�T�y��P��&��L��L
��6��F^��3��>&%O�;	���S �t�f�y�gYr��;�3������Jmž�s*7=��b�Hr�iF���+�I)ƪқ��"|r/, �\Y��?�YZ��W�v�r�9v�j�Y�&t���&�_qn��l �^�.��9J���O��ٿ8�قb޷�7���T�#��޷wE\���ת��^W�$�Ʉ���uFd��o�lf1#ޕ��R�����Q�_�0EN�C �Q��W��6CP+�f0��y��@ՠX��VIl+|*��ʀ�;�+7G�\��@=Y"�F|��܆�� �d�~*X
�P���GhiW��1F�[���xzK뭡Z�����a�~�Ձ���4`�������A)?�ޠ���݂�@o�5����*A���^)Pܫ�|Yw�
Q+�7-�}fp�g�Y^�a�(&Y�E�;zI+���]�H�����3�a.M���=��ڬ�m��yߊ�X�;?����:DGG�a�&��Q�or�.V�*�~dd�Nw�pᇾS�'�h#�.�y̍�o'�
���fYKH�!{Y܍�q�ҊWi!t�d��AH���w��3���(|x'��f�_.�
��i��wAn���e��!�	�6�wM��x~�1��/8`.�'[>(C��b�N���n$��a�l+�༭)�r/�2�	8ҹO�Π��Ү�s���_���X����R0�NW���ېA&c�V}�������ڻ��<��������ҙh��s20�l2�}��o�E��qY�������t^/��R���'�!X�#�������_�F>I9'�4x�'B0H%�UZ�_~�J3�@<2���o��^�_M�d%Q�˒ؖl�#���S�l�T�8�ٷ���VKo�{��F.q���/48��[�.��m�=��@��ouG�#�!Ʃ��E���=��sэ��=�_�\}���$h���F��F~��������#�BĘeLސ�5M�'�U�A����U,��]YK�r���z�����D���r�d4�k~�����~�5u�4����gm�A�9�J�jW���F��@w�JE���>��!6]˓���2�o�Ex3Y$6I�����W����MGL$�c�Z��w�K$�	39��y/�؁	K�ڮG�w�C7�4~W��W��9���N�����tL���^YJ�6�tg�v'�(.�3@�#�6.?��#�jwY;�2Y�#�ǈn�ގ��{�M	4�|�ϧ���Ӵ����o����7�1���z��g9P�DnO�Y�	��M<țqL��<��Yxlm��[Gh����*
�Ia�~yL����I�*mG8}����p�}�@��\|=�7�,�$勦6�zA���I���� ��������K����Y���a�����n�=�|�wF7��.�_=`��(a銔g���r(EEB �p�<�5� �r㑭�e��/ń	�ha�(�]�NɯT$=V��I[�d�N��?������@F�C��#����������IӰ��1�{1��f��y�UOI�U�f�>�zƁ$��=srw��w�-4��/�,lm8=�)��崭9Iս�&��r��l(+/�D�v��Ia.�4�0`������yG͟N�����9�$Q�5��=Ξ6(�Y��_��S��~Â5,ʌ�|���Ym3>/"ZA�����{Zݟ��W&J�iX8mM|�!z8��i�w��Bq�`�]���7��`?Brc)��_�=F������'����L:d�|X��#���_*�c���YS����z h��U-��/����ۆ:�Sk䅲����ꗼ�4i��.~s�N�V�~��(�P	YY�Oy���r����:����D����q�=�^&��'�����K�p4��|E&T`���Q3"�l� ���A#A���@�8�������M(�}*{@ί��#�!��c�5�*p�X`{���:��ʏɏ����x��Z9��ݧ�݂yL����,�,�I�B�~�;�!#�Cǽ9v�2n�/�A(_��5bP�^���y��6�neZ�VZ�ʃ?�d��;��ځ�(��yt��1񏾉V���eVe�K�m�x��W"Ly��� ��f�o-�$�Q_�J!�ћ�'���[�U
�Ɋ8�J$/c[�^V"�4ZI�%�06^�o�~�ۖ#^��o�3s�Z�����RѤ^9Y.���	r�n�VjȖ�-r
�sO����o���R.
A��8�
~%Z��d�r�u?h:�}�bh�_u�B�`[?=�;�Ư�(Mpd��C�vQ�)���^�<��1�]i��`� �9�
��־��yݣb���c%q��~��t�� ��Ŕ�J2y�D
d�y%)�"&���� ��N̈́���4G�#c *j��]�ȟ�tjR"�O�.�:m���2�Ne�gN6H�(��3Pn�.��>)�	�<oT[���[g�>٫X�����~0��餮�]O6�a�+��я�g�G�E�l�Tݜ�D��l.�� 4p�u�+���1�l	��]r��-��2�Z��_��H�mcK|��Q�Um����}��QxQ9��V8���� �������<K�_�T��^b~he5Z��$�@Z��j09LA�YN���|6e;��j�F����cιG~%��|�z(���Q�9�&O��I`ߐb_��Z�RA�� �+�Q�gg�5����C����k���wg�$ā��D@��ƙ�1Pr���bM��N�����P-Kg���j�N�^�f	��1�Bw���`1K��0��Ǿ�`�7�}��Rx����<J�W ���;-}"~�m@q�m-C,vc����}&�H��8,b��L����(2��b"�=�!1��{C6��JB���]m�2
���9���;R�������؃�?��
�r.�מ�Vn7C�w~\O� ��kT���Lr@?`���+��K.���{+k�w��$l�|�+��a�l���ע�Ύ�c���l�9R47� Q�Bi������g���p�<N)�G͚����a��\��m�����	&�X�P7�Mm_6S�p�1}��� %�����+�3W�K�����l�K��
X{�*��l��f�9,\��br��2��WM�d�kd�ٻ�n�
9m�����R��M�^]QiÏ�ћt�oL��(��$��h4m�ǀ;�\����%�ty�X����ʟ��ָM%��G ��.f�;��Q�Z�cj�C�������&�P������V�g��������ۻ�Fc� �0�zI:��9�_�i�6|4���'&�v�Xt����h����"O:e@�)�v��/EH���Bz��{��'1:VJQ� 4jhN���D��s�{o����X������6d���s3���������vq��_�%q:i���2�`�,�0�9R�Z�r�c(��_��0�Y7<��UD�5�����B�]`�
B����%b��N�t9HZJ�E�
up�j��+<D��[Y�������#��}�b��}�1�5ͪ�� ��C�l�͂@s|��Z��jno�7���E6r��q��݌Z57�KP��`����l�-��ӗ��0$� ��SK����q=���[>-?��#
,}�1I�/'�@��v�n�1z�M�v��tH�J����aZ�Lu:`�c8h��AH�����}����1��[v��bi'���q�0�5�G*��3J�3��W�I����"lT�"f�[�Gށ��yM`C�8�L5G1{��blї�j�p��>�<��v�-�7+�Y2F�����f����8�~&�xM�s�(9�T��%����&1ɩ��/����#�7��V�3E��� ?X:�<��*�Dv�u��sH\���h�����ƭ��2�bK���X��AZ�0 ��^<ł�4ok��Nw��	�7��4��t�8�=��9�7�4V��&X$eG��F�� ɳ�O�%������)�������< X@��x	Q=A�����]��tp�*>l�HC��<�>�BAT��N����{�9�tz`(����q�>l��#��?�s̌̿n�ZT�x��G��1�51t#�#�e����$tAnm��^�N���e�i��m��Jl���Fh����R����&F�tP]A�����"�G�Sȶ\b�$! �t۵�ؕ�O�/e��h�b��+�����D`i�wJ�F�!]%Dbի3��V\��
�����r;i�(��;��?�-M��B<en�P�<�^/{+k��j��|z\ɴABN*���m��`����wЂ/��#��&���Ռ���ʿ���cќ+pO�9CK�j�P[bz�eK�tv��9a�Yҽ�*n?m�Ļ����I9svIMt =,i�Z�%XA�2*�ʦu@��DŰ�n^)���ͩ����km�P��oA}KUT��D�F�����1�����XS��}Uۣ���C%1���|�c;�bu��F���&�XP�Jڷ���*Y�Ŷ��qh_�+w��
����n9� >˿*t� �N8��w��nʶ��pC�`���O�׶$��T��ٍ����
�j�%��� �ũ�$,.5ϥ&��
�&C��P��A��pB���L^�y]s�Hd�>R�36���>k�0��Y'�sgLE�R�;����_��1KG�u����1���M�:���A�i��ۗ ��סt�1(�4�8&ؑ�x�z��j����a`�JA7IU�����3TQ�=Q��i�71�����.3����݇.�mHw�n�T��5�V�S�:-�po}�b��j����g�#󹱊
r���>o,�4-�q�%jS�I^�/�-mO�?�a}�� 
�Xc��;o��J���/58�VS��zlDr<���K���ۤ����vǸ!BO��	2��@���M��?���FZ܃c;N�Q��� Z�+K�s���<��Wwn�� �*�Nd��ʡa0��K5y=��Vs�F�=�k�W�0�M�9 ^�!1#�|��M2��qLs	/��ͦ����r�X�_�(��)��{Z��=i�m��l�V|;G$;Xg��cz��ЀﭽE�U�3D��>C�r�:�����X��^�~b7�1:��#��P.s���!H�QYx�e��z[����Oc�W�2�G����� ����#4���R��>)��!�޴�
c_]��8d��Z��h��.՚����_�*]�RX����
Q #���:���������,��W�M-����Ә&0.| ���`��7�G� T����]�1@�<S��P�d]���GT�e-\�a�p����d��i6a�zB�'����?O�'�A��H�wS��_�U�<ހ2�m�Qj�aA������q�Z�����q���] ̉��y�=��R4�N�΀������|� �8��ʓ��R�D��M͞ws��d���dwjTpK�};��4� gG���_i*�1�����z�kw��őޑ�#�2'7�dMQ��>35T#��%2l��UY�ho����r˻!�9�Tapj��r�3��>P���un��lpA�Ǜ���Ę�9k=+��n�]��+V4zF�g5ϯ�C���'W`�`�B �O���]��H�ɺb�C���5Z{�!��Ғ����4���\Z$�Z�r7��Y�PS�&a�h~���&p��P�/����E�U�1�- d��l�{��i��ҝ&V ��q�t6���~�Z5Ƣ=R�,�	�`k��'�����{Z��Ge�(�q)X��gT TN��:ޏ'4��e!�th��*�s��J�06,f��|n}���X��&�V=I���`�Ah����X��M=���� $ڣ�T����B�F&r�����F��K���@�i�3엻�~J�xrn����NBft�t�:V�d5EEQ����k9?�N�_���_c��G`���8����AR�v�Z?$�TwB�vk�Za���v:����&�g���˒4�̴� ��$���On�LO���_C�8�Y2$��:~�z����HɱU�k����b&�NTY�(�?F{F_���0:�h���"�A��Ym�<2QGu(�g��{e�-��ܨY:����<����Ň�c�l��l�#v�4�T�x�;���g��O����3=��|����8���̩��c���`��i>:}8��딺��aD�寄o0��>��OI�,-׎�pr�R����y���>	VPf�1�Ӷ�UM?�`l�I��A��(㡂`-4��\R_�=��̢�ȷ��3���ۺ�.�=y�ܬ�N	�2�8ᧂ��)3�v�D����W�x��m��5v�7�f��C�D�?[�UNO!G�/I[n�^PX��ή>��QЏ�I�vH0G�&��=&��J�T������
ΙRp8���*1��aB*��
 �l�$(����[�W�i�.�˥�_fV�b�~ZCޑ͵��%�T�p�1��`����a��b����*BN�dQ�4��q���)����Z���|U��ס@D��/���-E�:&ԀQ�QD ��Vy]X�5=c\B�T?�/d0�V�h���0�<�6���L��9[��w	�E�+�/����A�~c��)���Z�i��Z���պ���&�k��ɘ��_�2m����'%�f���j
�Ny���������0:ЖK��h� ��{���cȽay�0�O���R}������������oܥ������Q��#��qh��:���)�N���E����%���"�F�����Đ��!4��Y��r�!c}�&ڵ5�CUj�,jHu�#��S��.�\������EȺM�ٗ��cn��r�����V��Ө�^c'v��7�����9Kfm'U̓�;�^�̣u�� b5�#ຩM�w!y�9���
R�d���z!����ӣJ>Ib�Nx-r�Xqҧ t����9G߃�/a'H}@].'�.?*��l(1p�����6�~��e�;a5�_J���<P����,PzG���I�˗�sD����^=�~�>l'��Ӧ��Ti�;�F[>Ap���(�Q�Mb;Rn	`�Dy$�����0�53�u{9�[Іm�Yl�у`-�o0���tg�q`�U�z���O�΢y����[wmK�+��^Y��+�\,P��$���0�/X��%<���P���j���dI�h��KI���/rf���4O��a$���P�q-���o<�7E����<rh�/���
A�9 N I%���)�>�6Q�{�i�����ꎉk���V|r�6()���)�A��޸�c�pKBH���M�B�$B���C�z�~�k�׏����O�1�K
�;��4�E3�E6/�.gu���k�De�DԶ�B�m)�tj�P}o��O��Ee:�2�#���=��R��'�ْ�����(Z��D�K�����=��uO�W|���3Y"q+G�ꤗ��s�ݡ�t�0���[�<T�qŐb�R�������L���M"��|9 *���QCx��W�pL�_iJVxOH�kH�v$i޿�Z\�W�9*�l��I�ډ���Zu����
�و��;Mv��o�X
����� �C>#���˵)bShC���8�'?d5����x��m�5wl��8ai�3/~�j~A�>�N��z��-�Eg�RcztȈ'm8�`�ou��.{_c+���򾥒pc�ئ�Ԟ?}Y���^��Jj�r־�I)�P��p������G*��ܼ�&]�$�`n���UB�F��px�_ɏ{�Cq���HV=�.U����t����%I�bxr�O�<G���đ��Aź��'�x�|���1������� a�*���r�%���z��O�ZoT�nY_�&k�\@�|R<҂.?;�+��F?>���/�U1���Gje(:Uu�&�\�"'|Vʊ�v&$�/�q���=L��
Q��u&��H{G�oc�+_B�s-��BjEn0A<>�חh��]<rI[��bA �X�6�f/��W�� 3��E0��5�N��-r	��1����TҤ�W��0��68� �7Q�r�����xsM��fGԘq�q�t����۪H�uL.�u���G{�+UY�]&N{� v�������� ��nŎr��X����Rω�%7�U�O>�	`��!���!��j\6=��T�ɺ@��^��c�I�;���������I�k���1�l�ҁ'��$Z]�yk _��| �is �1�����c`��I�B��[�ϑc/y�y�Ԇ��;�}��6�*�wo�%W�rO|Е��h�}�d3π��2�)m��hC,($�hAh�F�QY��C�"A�
�Mr����]��|��	2��|��6l���O�Z��M�*ZÑˎm���3K:�1���I�Q���}}˓�[}E���Jqƍخ&8Zk��h	��}&�b_�}a����`�;H��L���É�B��rs��@rj���
������%�K;=�b&#�C�f�z�FM��U��K������Ci�[���J��JI꠾-|p�n&�-�K��p+�����jH���5��6��0����E�{��U�Z�]>Uk�<w�W�k�����D�U�6���?N0J!4�[��qÍ�W�Z�h�.��6˫]�G}%"� nqҡ�7�W��3�u
o޻�q�f�Q/pۭ�|��I�:����@r������2l|P��F��k{���WZf�z��RC�X��a�3ys�z����a�u��@xp��/N	��6�Y��c����J���k�e��p�vN���������n�R���0�b�יE.�J�6�PE{�q����ҍV(p��58_�g1)��K4�5b�/�����-�lp�-���_᭢gɨ �%�H�}���r�k� H���X���Xu���V�� �0\z��,�o)�1����>���9�e=�=�@��"��_�d�tˣ�DF�oC��X��i�����¼��
[��8��ԣ��5��7:G`�=[��}o���s�07˅�h3��XV��T6�`���"�`�nإ��uS�!�F+(-�
?���"����Ղ�M$wE�$~�!&5�iW[��6�92�i�:�,r�6�#��P���?{��X���Wʼ"!��\���+Y���/�,:�P��+�Ҟ�Pm�S;��!�t|�����bl:TS�C��2�����qd�.Ҙ"!9��R�e+���^jn���a
/i�de�&*0l}�����j�<�~�'\G����To"6(�r�Z�t�t�K�/(�?J9��*���{�K�*;r�;��XY�N��ز� T���BCYƇl,=�B�A�߉7�O�=	}u|^ ���;Os�av:_��
l�ށ��9b�Yͽ�2sW�su���G���ȭV7��]ν��� jJ��a#3��l���s���[~��#N�ssc�S�g��q�Z_FI�~~4M�[a�(H�����n@��^��:X�"�<���y������kRJ�$p	͖0�zq&Ɂ��z'��[z���[4a�x�5#��h�4��L���L��S�ů���
�T�n����s
����u��u��/N��$�K�̋$�H�=�^�����A�E�x�E�a����X~�A���i�ȕY��������ѱ�$��̿�#���Ni�_�i����2,1��3A���#>+�T���Wh�^����E���F`R'K5��O�baQ0���"nT�Ùh�����E��gc#�q`�ֲ�����p�9ߛ�N����7��.�S?�DV��73ZW�,o�:ì�^�pK{JTf-h�.u��#�:���>�D��hu��(3Ab�Ȕ(dv���K'���7!��&H��>���jFsyB>,[A���+m��D���d�s8�vLE$��p�mILVI1�$HL=F��@��pJ��w����@8�x�:�ިk�wi�	�G1̤ȥ�i풩Dv�L��b�V^3�'�I�k��k`�Z�F����ȉ���;�#*��BIEE>`D���{��bD�!�0�şg���Δ�H��d�`[Υd$���R�W�J�J��d���(�l)�,��j9z� ���C�I	禜���"&�}��k���ꡂ~=�=3���`�*��$������@�\g�:�hca��+�[7F���qhwu�y�(*�j��/�.��P��1�O�8_W��I#m���E�������xs�i�fW�-�Ȏ�iF3`�Ff�e��zu�
۵$�BY+,(��Y���9X��T���e:�A��Ո���]V#��Z�>ᒥ�.M�^��"��{vY����M�O�4A�Xt�s��dR�K�JZgKP2.��lDz��]I�o��x�!�nF����,�4�	�6
</-�c���UE�9n�����+�}H���[��Z��kXeo����%���̷e-����VMR�5c�IUjx��&�#�!�'��}Ifr��L=Ց��&F.:���-ex��<��|����>��v;�H��:!hb�{\F��h}���cT���XWPnB=�؜��*�݇ �{�s�O-������9хn���;�VL=K�	��{�!i�F<�n�ט`��`�Q�HE�.��]�`�C8Y%�@45}ɹ�X[�����K>b�hb֧�L�v�8��b�
K�����&_EnV��'�Z� �k[����p
]�5�oʓ��ѷ�D8v�������,¨��)�K����wcxȂ�F���_�d?�L�{�̬x��ɭ�g:���\S �:=�N�����$zK�Lm8�������Mո��{�μjɤ��=-'���9p􆻳.��g[�E���9���)�Q^�q���Iz����8�I�w5�B쐆5�n7Yم���L5`2baH'��ƪ�kM���r u�Iq���%��⮍��ɔt�DF�o,�!ڋ����&������\��Z�B�a�h��q�� g�=r���CY ��zi��v��)���"!e���չN��� c��X2����Nc�����Ʋ���vz�+q�:��׌+���޽'?���ua`5�w��J%�x��}t���g�/������$c<)ز�n�V�`dX�Y�<sj�vv0�x�!�6�����S��F}��%eO0u6�ڵ�΃�%!u����X!0�J�Bދ'	B��l���÷��>�gʺM��b�M&']"�m>�!$J�m�Hk������U�GS���{g��H�E��rmΊ�S�Xo�i�jd�"V� W�X���z�����}Q���#/��燫�&�n2dۘB���+|@N�2�����ڍ���TZ�׵�ʄ�)]s���+|�G�:�䬥Q���2R:��ߟ	�^��jy�Z��ފ�އt@�/M��A'�%
��h�u�,p���n3ܠ��B/��.T`��2jc0�&�<�Ej��,K�?�x��s�]���|`��D#t�ܽ-��4��*�n���E��b������&�Szf(SQ1��{�����
��G�gxF9P���zUg�R9`k�^d�m�����@�����S �7��@e>�#�Q��A�xic���X1(p��������>���/��t+S	a-���O��:DaH`��w�B��]�M��j���-��k����%D��?U����d�0�������^	�X�V_�盯w���&�E�^1~KwԱGD��i/�Qp�[�/<+�v��t��W�'�ꟽb6	�o��{�q��V�fM�#���Y�@*�Gx�y���u�@p��2Y�\[��.��y"�+\�Y���&<_�
Òz2t0X��<���H�>O�'�m5��
a=��Ȼ:��Z����-oU��1��L�Q�n,�iL�V�	i�ᣵ+��+W#�YD.��91���K�0�Ji�U��x��	M1HMr��F��hl�#�^n��MW9K�Xǡ�A�g=ۏ��C�����K.�-��s���I!d�~�R1&�z�L����+�����$&"]��jz�p%�ϓH�*-�Q�Pf[�꾽c��������\���{_^���-�S���
���R&C(^>�D8�m�����j��wƍ�d2��+�4�z��P��E�l��Ձӝ0#V؄v�f"�
x��В���޲,���{U��6��P�?��k����ړ�=��39l��4ylX��7����߭�>`UG\��"���u��4+f�ͪ�Of�1��]��F@İ�r��-����W��,���I�pD#2�����Td�T�
�$�^F���L8���	JY��	�A�(;+��h�I��L��"���������xf�?#&)f��G��U�J����A}/�Mb�6�F��!R=	�J�l�F�xɁ���{���w��x>�F~� �\�VK#�`!|�V���*�h 6b[��݃���%��M��4l=���5��;W����|Z�Dyh�[8g[�x9��$	`��kט��I����xO�=h!��Al{����~���\C���S�q��f��n�댇��`$<B
KK��N'��j!3/���]xI��i�!VD�B!Ҥ�C7��.3M�P{��'���B? 4�:�4��7���m�;��,y�WQ����Xs��iO��pW�]l/��h��x�;-2��C��Y]�Н?ya��t�h�J~~8�f�ʽ$,�,(%�%��u��k����{UߠJ�����2�OW��c��<|M_]�-����Gs �i�$�U��y��XMP�Ko�*�n���Tc�e�Ƹ�8�_�by1���ѱ~x��4���M;�O_|��Ϻ��b�̝�AV~��O�}4pYQoV��Jj9��E"��<�I��`d-�vQ�vE�c�ŜG)_��V!�1���ȋu�WFWaK��X��9Q�Yщc<�B�y�
c8z^�.��1�q�Q����2�t]��-J�S�хLy'�3���c�����Haw�0>��i�q������2֯��oX3x��ΐۉ���ղ��P�J쿪���W6zJTU���
g8H���ϯo�H�%jt?���@�*���6��,r�+Կhs��`l�X9���p��]t��^��7�����V0��V]#�>?�ݼ�|���(U���F�Jb�Rb��;������Q;2�yG�O�������T����� ����yӓؠZ�D���S9����l�33�asZ4h�"��M��PzQ�$�<�Ui�����qj#j���PN�'|h&�+��{�f�ڥJT��E>��-�*l������è�w��=8;�k9q۪I*/�����lw/��?�Ŭ� �׷�!I��o��\W~��|rCd�E��	��v��Z��o��&��9_�:�1��~�R��fV-�i#�`'c��k�f�����[(M��MRSx�`W�2q����=<�m������<V��&�V��-�b� �
�*ܿ�����L.L֗l�$������Y�/������R�?�c�7)P��&<o�@_A5����9��k�OY�=ji;DM͢O�����������A4��ySԼ��Wק�^�T�D��WJ�77Un-�ԕdj�����F"�Y�a_��y�,v
����gS!�K��[�Z9ڈ�mTT���x����יG�.�ͽ�[5rl3�>�jr�/4P
C|�3?)�g��J-ߋ����V䢳C�d�4���(��; 4_ -�P.�E������߂K�S��j+��z���S!��ELb� ��3֙��D�.����q���L�=���Ly"���"�!a?xfo����-�]:x\s�ǌx��屽�C<�t��&)C5Lo��t��cE��l�B+�5q�:������!�jY*�"����#�#�JÏ��g"E�u��:5�l�?�+���޿h�m�\v,#������Q�h�@LF�b'GGnr��81�{�0蔌d�"�җ^=>��)�Al:S�?%![Q����o�4�-Z�����3�g���K�N����]��[�Lo��mro�n���^�H����K�P���sA)f1yћ�c�9�S��γ�YE����~���q�;�m���ܐ"Z;<o8�˃��O��&h���ȮM�̍�e|룸Dn_9j�{X�%vE���a#^h����T�F��\?4D.���7O�����ḍ��d�F�B���F�aa�e7+�9B�����D/��J~q�S�lQ)ԛ̵J����]=�����S�7�It ^v�J�cX1�ٿ�I镁�����;ng�F�`�����M��g�2 B/���}�S+��dN%p�X�ha*5�r	4��8��MSDR��~w\@F`Ɋn�i׺�՝/���Jg��UX{〯,C��ޥp��tJ �C]��	ٌ�	 ���S$��vp��Z�#�;�.T$A0�a���Z~�Lv�7��&������H��(�D�9�=&�g��L����U�R�/�6�B����og����q\�S7����Ŋy�\-��i�W���4�Y�p����Q�)�܆H%�=hl��zN�H� �E������?�)��*HԔ����ҹ���xqE��M�Q��Vr��t�D��$������ m@�&�a eF�UTߟ�a�'
�;)�B�x�Bg��L�|�z�>��^�mJ�����������Q�Lx�0o��Z���7����@4׎��������/���+��<����,��uF�Ə�bB֡JCF�)DI� }jĨ�Z��#)'�*�F<�������#�v���RZ�yue��
�q ��Bk��f�ម�>��x���a(wxp7�˳�F�v0r�m�����14OL���{��B�ߡ���/=ۇL����-�#���p=��N餈��&ފ���٭th�[�ԍ$�hb��D�)�'��+ԕ��!���N�Љwb��z�vQ5.�o�}�����9ɿj���>�S��)"ȳ�����/��J�!⋌�بR\	��F�j�1��:)��e�p��6u�S�����ٟ�7����2�ũ+��%?j5�浼{���;3������i�L?lQ�-�"����(R!���-�f$��i�XZt���5��%$ R6�ҝ�9wp��M�y+h��զDE��X`({�B�щ�;����Ua 	���pIJ(|=��3R����t\� ݃p�����蚾�ةW-�<�X���,�D]�c�b¨�Rg1.�!lk*�8�A���V��g��ïo-�&�z��`8~�&f?�=�u=}��f�*�0�Q{m�|�=m�z�Ʃ� \\�Q���d�CB�g�]�acvT����yY���?�����J?O�^�˃)%��?��aG�8�:vWά�Ӝb�]�������Rv�*w"����S����.
� ��#Z�m!Rb)�X-m�$��#G��K�?)R[�l�B"�!�<�|P*�̏��V�GEd����g.5y��WNE�'Y�VvG��r��ŌDϒW��Z%�%^c�\�m�wm@�6�~�<&���橈�x�	��+��۱LД��]���W�������p��E������a#����P��Y�x��,��}"Z�b�9���e�i�h���8c��� h��ϻ���j��Fj�$~O�v���X�ޅ��c�Ӷ�ځ�k�,��q1R
��']I�jk�{��h�Mv.�ǰ�*�woOE���D!7i ��O��;��HӒ�pc�σ��~U��,�F��1�0�H��T�pi�']hck��ؠρ��n��?\�a� �V_$AI��4	YTM{�P�'���<X�"|�]ώ6�8�c��"�w�_Ry<�2�����ߚ�����o�R���ĩ�<r�m��a�D�y&��|�Vp6P�c���1�S���`�R��Mq�s�*q.TE֤*n��ZyIFD�c��E���zQ��:���~	��^�^6
!�t�'ጊl;h�g�:늶��C�G���u*کJ��9mP4���q(͜Q��Y�h_����=C��2�?��hp�)"�,ȍЯ19��N�5�L3���*Jy�8צ��Z����ZTN�f��&����4��}gm`�� Ȳs��i�'8E������$}ע�
]���b���G)G�4�̿C{��|K=;�:>�B��6j�\}-�+�0�}&���G�0��Y!���Q��B��{�_�Nx_Gʽ��.H�?�OU~y�~�ㅕݜn��05 Ȥv�N�gYB�T����@�o<^G��W�ȕ��ɣ���B��\𘮙6z	���_&�?
���	�}P;3���ac�(ә�<P�3j�Iy칲�T'K�E�F����S��ho�J3�eZq
�y @����c��8�xRHT�
��1�R�0�h4�$Է#�DJV�\���)7�������͠i��?9����M��<E�<�8���&]JV$�צLXӴ������E��7G���-���b>���I�tu�;tC�1�tR��5�.l�P[fƭ�a�����A_�M����9򄚴���/��Y�X{��͙Qɣ��/��վ��}���_�j%Y�������},5��``��Yy�&�ܶ(ă/���Ǣ~Q���a���gy)���'���
Wՙ��M����(�������_`��b��Y+�/ j|���*u�&qNbC>�7���N:?���j�i����q��T�N��y�tOqb͆an��G�'_��&����H}�w���`�>7��d�)��4���Q�Spv>~q�1+��S�0w���c��y�Pj�u30�`���z��O�y��xܪ�Ё�ì٠��q8N���㡉��F��{��6�O3[�Ml�F,�B�\�.�/����NCU�|�c,_��(!6��X*0K���Ǵ��k�?u|qJ�����qRm8VZ�22;l:������Fez<
��iB&�z�)��Dr4:���͔��$��9�6�=6�ܻ�?c�n��3��"�1d,��u� �!�zŇ���G��ӯm2����6���zW$B�#!*V���� ��b$x��(kn�;��%�G���
՞؍S�	���;2!<Q6B���>%�t0���:l;����<9��d��$���fJw�>�Q,�1��@�	������uȍZ���7��0�p(c�	��tE�*q����L5�_���8|���W�o�
�S��p�U[��x�/��s3�*��|5Ƞw�	��ݭ%��D���QײW�(Wà\��>�C�$%Y9*��,Y'�?.	�I,ހO�~Nv�_c�%6�s3���X����F,���	�w��4��it�{\��S�N��f�w�߭(���w��m�;�ߏ��e�X�;�-\�E%��=�~Z�M��f&g�?��P�ح�gg�/�]�����F���޼��mI�1��Tu{d򍣚SG�~���hx�i������F�{ �-ԕ�5����d�22��	�XU���H�@͙�8��$�h@�+�~��NH]�`6�A|�{&kܻ�oU�j@� U���>�n��څJ���~�\u���tL�2�N�]Uwޱ����ϋ���)-b�(;�\R�(��d,P}�H��i��u3) �a�w�b�3]��Ȃw����-�`��o�������c��.:�m�SHS*+�Y��i&��܆8yŏ�ʬ��^͝\)�oݽ�_�mZ�k
qX���J�@L�3�	�|�I�����T�7�d�����᭲b�����tU�q��Q&l��H�$aO�( =Ʌޚy�P�ԪW�c�
0�R�XS3;�m�9�/�MTP�%��4C��i��(�c��	zTn��[_��E�S�t>��י�x�|zqk!+6ɠ��@�e[�FO�Q�P�u�:3����|KE����(��6="�;ei^�	�CƘ�-
*\��!͏Sܾi�Q	��e#�?Z�����P�7�g`��)���?vZ�Nx��7'�kc����ݍÅ��f#��\���3'�"�2I����/-�qL���n8,��b�ChJ��ͬ4�&>S��s'i�)@���ڙ�v)��%Ko@{� �q9ɲ>G��F�e!�?��/���6����'�ݸ�ԟ�a�1Y�x�$&%q~� %��� ��{D��%���A؎�؈�t��l����J�(5u��.c-����>��^=��0*�:BC����,�D��-���g���D�E2!�u�ƷI��`�����{���55H �	��GR�S��+ b��1,��܏�z��>�5��:������\��L�o8��;(c�_S+���U�ͱz0�///Mަ��Zv/�d�_(V��#JA4�9wwo��%�e��%���2`N�f�u�f�Y�3S?S��֜�C:?�NN�#l`��
g>�AZy����d��G>o��	"�$��yO)Xg�!�Z���<<�Ǯ������lN}��'�6i�pŨ��K�.-#!���۹|��wZ�8��:�����e�~���/IWe2��	X0ǡP�Vb�u�DT��]��t�}�}��F�b�D��6�����e��&̍��|��6aB��2��}޵ʶp�)���[Z�p�W������k�F��^>��ib�>�٭8Nw�h��sA��,w85�T+�Ǿ�[���D9��V�R�` G&�4�ߨF��������h&q)�^Q~a�1��k�[��s�|�p�{~��ػ�9�"-������4+)-�8<��
��V�|�Q��u,��O�/ �o��TM�G�'�Il�+P�������vja�j�3��a�,�����)�9f��c���2��^���d��]~�mi�?Ël>���t�"o�����s����Q�\&h��x�T�n	�/�Pq��΁�+BÙ���~�a���б������:X�`��u�"
�b�A&H�F�7��]{�6TL�m�����t<=��l���S��Z���%C`<��o�-�A��*kN]1/g���E.P�$��!���!~�c�?e�M�k�.�`�J}F+2������T)sy�R�y�f�X�`N�
��b���Q鲫�����'�p����x�5�����L�}Ӹ��Y����~u�>E��c��"e�,�>��� �����P��
f8f������ߕϦ��Gb�ȝ����UǑ�af����b�����H�͟�A��gM�<�I�K��a��ϠT��T	������l�+���ai�����ۛr���	���K:�$F��
�Tc&��*X{g؊�������9�+����_�������#	�P��P������P��?$�5��ݚ$#=A��1,�*~�%)́o��"�!v
���t���jw멯ȸ�����7�#�]��z.���l�>�(Z��^����1��=�?��[�P�l��C�fS9��/��y5�����zє�-���	  \m	�n3f�f�t]��C��WÁ#熞�V>�"���/{�ۂ|骦��)9���Z\ϫ�ՒV�fۅ[���֔oYu!�~9"kIY��cO��O4ժן?� � A���N�J6*�p6����i��^��5�m��W����M��.!0vM{g�Ԙ}\���W�!4#R:L
�|��>�MHW��lld�G���1�+5�ۢ}^���4z]���@;?���=�X<��k������~M��w��kQᣞ�Q�;��su�SC���J�`�/�~�/-u>�O�opT7��$��QL~YKa���fy,�V����@c�A{�=����M�\�}3�O)#K:� \��Of�@���"~r�s������t�s�*N$��(�"�bl/q�i�����?)Y�ĭ�N5ه��j������h�;D����8/�:�8i�T칓�����VG4
��rGm�������JjWl���٥�����]4�h�e:��h+���;���C�"����Z�c0g,��\��t�EW�(�(�A�h:O5<�Aq�L���̀�]qxG�&X���W���mG�|E�jJRꡡ�����䅬���D��"��cX��blF�M!��)Q� �o�K�=!�������ɝe�Ζ&`�v�s,�a�>䤾Q���س��A�*�Q�;ǘ;��l�Y#]�F�����k"�«�m���9��s��Ns��yj0[��z��n�>� �� ��s����^��شM��O&@6%�}U�V��.0%��l�ZrQ��� *D�<�7������A[�8��ܻ��E�N�Vn�7ܪi�=x�LA�k7_��.���Պ?�T�m5���]�nB��r�B�y|�B��69a����z+���z��Meݖ2��D��)-��k�
��<��/���}%��4V>�	���L�gL|Eo�w?�9x�B^�ca�'Ԃ�&��t��qb�c��y��jW�h�xm]�v�Y������js�&#��C�:{`z��}�x�&7�u�	m�[L��o��ګ7�[P�|aL' �tV*�W��{�KZ�1#�ـ�8�D��V0��IO!;����6'ЂW� |pu,�Aͷ�s�}J��br��'��ܨfouӠ�#cYn������S/�'��s�/s�:��2C�e��F1�+�-�`z��'e��%Ȝn�g;H+�7?5g9�>�N���T���\�C������C�0��#B�Q=��g3,�aT݌�Q��
lO`S�/�餉����T� kHDr�S/\"��~<>1h�t�b��i����;+��~�w�5���ohǬp�J����5P��ܱ�g{/��T�b�g��*�z�*�r.]��em\��>��/4��5� �9kU�%�����	cl�z���L2E��ޥf{v���9çɎ�2�)/Z\����c[�zk��/g�W�9T;����q��Fx�zYcm@���8q.�˲R� 
���kyU�vjf��A��*n_�݈c�%�FQY����)!��}dsS��k�Dw/v �z.�"�q����kռmF_鴐�N@)(��#�+�������Ե����m�u���O���ز��]��hz�2�UNQ���=i��w��ϓ(";�Ye���<��Ey.���>d땊�7D?��i@9��(4��6�V[�:��&W�&�0r����<��JFN�(S?X;�\Pc������Rޱ�"�t~3����a�(�q�JE���'��٠�	A͸�nD����W�||��O�)�mF��9���4��A��;������0�t��`tN�DDO�{sO��(E����Њ�ϏQ�%&l�(��vM��##L���A-��I�T	N%����Pb�2[y�0����ͯ�L<���t��C�f�a}J�C�ҁ��V|�;NٶZ��Z+%�� B j�P��k��	�?L31��3��˽�d��<gs���n�,ҏEQCmݟ�_�; 3���ɨ����n��1�`I��y �����2���5W7�Q�dt�v�&6�;����Fz��ݵ�&���4_ߏ�q����������m��*�2'"�Յ��V�:�T�mOX�j-32D���'nNm��}4��a�b�4������L�~���aO`m{L@/ן�έ�7mr�T��������c�k�$��G��v���uZ�R�pN�'�A��i�N1����3�Ea+�"0�N!VwuM��/�4n�*N�NL��*�X��"�����7���JS̳$�L�J�	
	w��#_�`���a����l�\dyOeqiO�{�b�6��ȩE�P�C ��5���6q�c�y
e�E��fB���6����)�7ⷜD:x� �>�b�|�,,����nO?���As���YF9��bm��~����F�]��L,�'���j ���v���,Xk�I�d���8{Z��eT���
����S��x��>�	|�g=���z�X�:c@:����D�a��>�O8����B��;)S��Yج��]#B��t�O�(�/���r;��,�k�1����=�0�͟�A������g���J���<m�*�t' pPU����/��`��c�Z�����JR��x82��+i����������Vq�D��l�A���:F$s�REذ,�����
醡��>�N�[;�ć�&n-��kXY��R����s�Q�}D>�H�\�u�g��]N�p�����&_�b
S���#�m�fm�����>Hc��؝5���H}���ęr��H1U��K����;gX���<7��X�Cg�h3��J�*�C�}���H�͔e�#܈����?pN��I)x��=D�SmH������^�G�C`��6�D�O�ʮ������G~�r[�W��ۇ"~*��Y��1Z������
k�[��SXv�X�i��-��a��a���P�b����s�4�����6��M�1�t�x/�w=���J^��3t��X����j5T~=S@
D.����m�J�r���e���b���'���͑��<x��;��h�u���2�Kc7�1]Tj,w���.B��ћn�;"�A���0	G�\1�h�l��Y����E ��H��,���<�ŕ�d�p�V(��x.ɠ�����<|r�'� P�j�R��!gCЌl܉�H��>���$�����	�K�i~�(U�&�� -�|nB;�����m��u��!��E��KD�Dm,-�`|Y?%�2���s+I2=Uy��v��u �ͫ/
�x�e�d�dg�Zic"�I�#���S�>� �_{h���	��^�T�
n��{3����kbx2�����>�����Ձ�]�b�zX��a�<���T/0IB<-5�8�sb[":�?�OZ�i����
�W�D��i�\�f.��(䉴�F�[���Q8��4"}/�,�Gv����m!�Ox�11��ա��@C#����y1��ʝ����!f���*�?��1�"�n��"e����s�p����,�z 2�k�ж��2����t�A q���mNM�1,{
_�r�[����V��F�4���x�~��.����;��"�����ͮ�@Q���n\_ը�f�;7�D�=�c���2Z��Jr�M:?��*Z:ܢs$^�9%�M���\�������3�8L9�"w$O侸�/E{��L(������JI1�t�b�*O���V�}�<��-��*y�W��(���\0RNg�hU3��3͂�v�"��F��Z��Õ!1b�tqL��]2s�Q� ��m�����lKtd�u:�u�����V( q F��a����-�sI䔭!�0A�����i'�Qb��ܘө<�N7�m���+ɭ�,��������a5y��|��u��'�w�d��|�TaS��
Ͻ�h&�����~;�W�e���!=�,�&
Fg�f�7f"=�
ځ=��_�'S��Tg|�y8?(`�b�r^5�3�{a��YJ����U�9��(9nb��07�R�Sm�\���z�c���hpeK(H6�J9X5Ӏ��N��]9K�$fSq+H�V%���������7X�.�L3�P� ��s�om��]y%�Q��~�#j�xJ�����v��7�\�
fp�������[���to�X��DBa��Z�d��l6$KJ`1�_VҌZ��d&��kAՄU1����ufL;-�e)̛��v������H�!2��,����	d��<�u��"�$��8�B ������淞���Y{�7�7������0E��Ί�]�&WѼf�ť:��*������SF���T�g<���B�5�Tp�Sހ�-��g�9��>�yV�j�V^��^��y����4Գq�����u��\e	؊f�:T-e~�jnIO�ԛ�%��If�O��ܴ0����CI4�1�-�@������X�U���3�(h��&{����iiE�pn^C�Vs�̜�[�����֡Be:Ɨ�������xƛ0�X����Ĝk�c<�z�o-
�oC܇uEGYDz�����jړ$��aCï	� >���V���5��m(��|��z��էm��S�6���f%��ϭmS�\ŒEk2-�:ǭ�I
�0�P�.X@��j��6��u�8҄�C���9ח> ܝ��,O�+��2[%lgZ��y1k��	uD1�ȗk5�p6p�9����d`y���R�Le���c�Ɩ�ۍ�m��~�Bχ����p~�I �$X�La-\_��d�}�W����"���PR)�K�Ak}P�Y�.j���6�'5m�N��5'3e�0|ٝ�B����o�[)�>�5��5B5z� �L7nq61����:�̃-��K��h���eL|�S����P�X'��1���}V4���:�����g��<���s�aG�`J��C�X� }"ks��,�n�3����=�fu�2�>Q��2c���$�só��D���:��ٯr��:l,.R�Єʾ|�P1�5!��$��#� ���~煱�f:YЗ?�V3�p=�[�Y�V����beg�����0���.>0h�:��p�c�Vz�.�L8��U�E3��x����_K�^����
}����K���߶���: �?F��)�D 뱖y4^@>��4֬z�.7� ��p����.3']f�X���_I�j��=ݑ([����<t{2��ò�p١V�D$1�gI��H_���fW&HL�#p��zl*��X��3$�������Rf�F���I"�U��E�Iǌ��B3�����j� <�!���b^+�����xJ�����j���n���M���s�8"����Ѷ�����"�g�U��^���hӹwު�6�?m(֕�&"�p`�2�t�V)�LI�+8q)}ܧD\`w�]�c�RP\�:��[��^��1�k�V������,}P�����-�ٲ|3����<�y7�ˏ�E�b�i���B��Ԅ6�Q��o}����"���
���.J�_��6S��Z��g���d���(H���B�1�o75MI"6*�Ng���yBQ3vj�Z�.��x	>��K�-rٶo8��ќe�N�fj�b�Ň{̌�1�N2�z��`������`>�ڹ���+����gTtU��+�����/ޮzu�D߲~�W�ág�w���U�Rް����8"s1kO��XP��Q�˩[p��7�,�G��W8�6C���n�\6g��k��N�m����{w�h'G;�������wEpż��:��k��טE�v�,�+-n,�׏F�i���
�8�>��L��C�x��d���Dw$��m��ۆ/ϾG~{�e�9O%�li�0a�
2��?�س��1 _<>�=H���T�@K�B�ɴ�I#{	��5��@�ws7�y�:H�Ht��n��jBpO$�g��Ĝ��%���b¾�şϒ�����t+c	x���]89�휄p��l�=��a�S��m��f��a�si��{	g,���E�:`�a�*P��%���Y�T�X-y\3���$A�N	��ǘ�L���A�z�8�*�N���7*1�J;�S��rJ���L ��%0���|�
⪵B.�;4DP����J=<ǋT!�6��ėtK�ܘ�xA;Z1�s.I{�5f((���{��~��
癭U.{5�⺇�p�w�����u��YY܀zzP~�.��T�:S�qV� 8��Ou��\Nʍ�P��Dݣ����!�H߂&���Y4���|��S�����4��R�����<;l1�)�Cb��1{yǭ(�޽�-�:v�SĀ��G*�1��=I�:y�|Z@��y�2i���G����;'y��;�%�=q�)�`99�:�vQxOemu�GLc���sޞ�R7����¿��5�7�2�Q��_l?��_u���A������i��߭���-$�n}Z�X�Ӡ�}^�ʣ��p�C��څڶ��
[
�VuP�3&�N<^�@r.;J]l�`�l������݉��d;\8,�2z��d���S�W,LaL#P��^�᪰G�%�/�&A1O��,~n�{�6�͖$Xڈ�t@���p�Q���u��j�������pQ��E���B��������P[�ԫ���ݝ�9n�l,�����4��e�#���޾� WM���n�̓p�2�RI[[��)^�<nM�>��ɿ������NA�����ܶ^�Xd��Tg�_Yoqg�d�n���4�w�.{8S��&�Qąh�pt��d<}1�o����fDJ�oQx�!X0W�F%��jp)���>�݌7fl�i�݅Z��+��4e��E_w�~� 9���\ɣ�ԡ(�OUv�*����y����<�����l�؋D�ʛ4g5Qo��0~�)U���l�����L��_��-Wv'}}ZfD�x}���T]�Ah�����cAu�@���i%)~iAr�W�x1*�LA��Wg_9��xY���[��1<;����dI�8\�Z����O�}�|�>2�us��I�.ʗI�E����7c�zJ e�z֢b�7.�����qB����ܻr@�nE.��.il�}&��1�''�{d�R�^��Һ@�Ee
�������`�Ki�+'�JW�e +�݄��6
����(QG�0ǿf���*e��3h���^O�U����O�l U-��s��/u,m8�j���J���wGN;�OMOor�Nb��������'S�������a�5����)
jW.�Y|�샰��:��E�}�2>.�c�}�~�Obّ�?�Ư�>��c��W�]ǭ�S����`!��
�{�)%D=]0��<u(.ߪ�v�s���"��ɷ:��C�}^�����q�R�5�4`>�଒@;�κ�-X����*�`D)~��E��$X��Kᑲ��^����H�5���]�5���?�ލ��GSh��&H��b�Ѡ�Ջ����a��M=rt�xn�+A�1Ȟ���ASMʱg��	愉@ݨ0~����=c�����c1�����;rN��6 2�%��榯\�J`���#\�P�z���9��88xZd�y��9��zʴ�*\<�Y}��|#Ez����d�<0���v��J,�N��1�"�f�y����(C�:Gd� $}��E�Xh.�5;u����L%����>�R�qn��=z�������?S)�l�
l�	�P�ɇ����� �ф¡�ׅ� ���aĭk���r72i}��yN��~F�h�/yc+�YJe��Mf���NO���u��EeX�/y_@؊�#��R���@�c���7&�*|�"d��.��iN�Vɍ7v�<�T0�^1&��&H�*ZI���YMf<O�9O>Q}ɂ�J���,"����B���톴�k��oC<{�f.&Z�;��Ly|ߌ��y��g�nQ���SE��yز*�ο�-��E_�0�;RU�*����-�$ �?�K��	��\����:�B��yv�[��D��7}��w���s�{]��op�����<9}�,��i�VL����0$>��QL&O��B�\��.�=�����x����}�_��o ?deX|�_��1���>�-�O���r���k�6�[t<��mtH�/��Į|��ߞ�[�ƌ����Ja�4q�m�h�\H�1�^���'Zˇ&�Erk���Ň������1;p�P��,�6� ��d���2Ҋ��O	˄4/�z�l �J��Dխ�Q�q���8�\e����L����zhe�Dy�//)�x���y�W�����;����d�&�����&�����#�+�b����Q5��:P�H/�W��C?��A:�,��J��˳��@ѭ*f�+(���knh�H m9T(��ky�"b��eP�L��� )�����u�5YX�H�{܎�h��l��j,��{�D4#;p�����0�H���Bv<[-]1�b�J�_b���}
v���F .�N.�.�I�Ѓ�K�I|��#?\s0(����0Wnu��J��KD��Ԩ�mN��k�������B�9p��Кɦ9y�-�du%����YL�'o�sQRd^bQ|3�P��nSkM�N��T4S���FLh�ob���[��2+@��Ꝥ�л�׆[�vLm�������a�\-s[���2MO w	M���I5��D���HV�mIG�itD����D����k��%H����79�ͭ8��$MWti���#?�{�4�f@E� �tL�#���i%�z4�E�?^d�;/���V��ܹ���J|{�C.+ U�p,��,q�N)���˕�{�sq2� � X��:�OB���OP8?��W~�zG�
?�.PaА̉'�]��0���[� (�ϯ�f{�P篗���������#��͑g�4PjL'?��H���]��&o�=�kя�%e1���>7��ˋ�^��q���޴t:�1��׀`x%cT�ʝ�Xen���u�+(Pn\�TJp�������1�'��Zad�Z�z�R�̖�jDH{yM�>n1�k"eԾ���,2a��^�/oP��7�)�׏t��bt�7� ��Z_���h�f̄�bBVKg��?�� ������2������[�G���eG��pph�^OdO�b�^qB|i�:���
"��W7�^�3�Rg�<Wh��ゑ�*͇Yc��]|�K�s���
�mN�e���������ʷZl��w���U#)�T�e���&�[=<!�9��R��R���۸�Y��4��`s{\~5(��8�T%b#�n8�h+Qg�T�R��Pk��zΩ�q����Yg�){��$���}9��Aqk�KAJ_Q�)y�O��u����~�Z����G�J���9m�����%|���af����t[�C&�w�$��nD6��T����b!`����Wm����g�/��9!]�*�K;E�ֺ2^y�����s��3vUv,����&:T��؁���JN/��3�25���Ȃ��BB(>H���졪�NE���SX��r�>0�Zñ�-�aRvn7��c��8?���x ��5o���Y�YC;�@��d˷	��R����a/�w��K��P��kæ-PB��[_��_�0���5�1@��`P_�o��#�_�*��4� �4�o��<� 3�
�<���*�M�[�P\��OѐF�$� ?�aw9R�� �0]"}R��^b�v(�4�OWpcף����]��G�c+�;�� o<�#6�I��h��k.=4��de��V��Q��>����b�9(,X�hPen
�݉	\YR���ɇ�P�G� |��J��"�}��BCF�.p�SE�7���=1�PM#��Hp�t�$ ˲G�}���E���h�EȤjl4�1�ŉV�rf��'^Y1Y���{��Y�<�rn1�:�|����������#|	 
�.s�,�T�F�\�j�1)X>&��]]����W��"�����(�����x�[	7C���a�C��R+�`�61���{<�:�E�kO�)XI�j`�%_]�6�]ғ`�ɻ����8+˯62�Y�Y.����*,�_�ݑ��Y��_���@�D�L�-�Rff�fa;s�*Ө�x��[�����g�n�R��x��j�"-����X��dn$�^gbg>9B��YZD*~�W-�Z�UHDp���6�m�/�?�������V���J�$GU=��\a7OF[��3�Q'V�%Z7q(v��-��곥���2:Ӿ �A�k�1�������r3/.��c�KTQS��8��t<Zv �����q���}
6��y�g}5�fb���S���%���jj�j�L�r�4w�y��d2�]P�)('G�s�4�~�!]��'I?$[mr^R��XC�0�ȹ"�;H���Sc���t��8�.PV��A��6��vbU���.U
ѴM7��iBN�4���=�1KB�����Da�l`D6ض�������ұi��	U"�Yw�k	2ِ�2�
�ڮB=�7����񤈌ܦ�x���*����vt���E��&�%��Kf|`���PI߅I^��\��ּ�p���x������W��Sy V�3O�sY�%�QR���v�:#��[�0Q�/3Fz ��u�E�ҫ::�s�|�%6��e����#�	[<ʛ�T,� $T���-�?�������>y�ST�IAQeE蕩��b-��~�2�[?:��M at	�f\H��� 3Z�H�tǘ/u��S���M�s�9+6��0?�Z/d7�ǵ ����.nؔ")=
v�PEz�%AE_�H���o3ϲ%3n��9Ճ��� ��G�"P�� <@�s�mG�b�t�y��A�$g
 ~���d�`��&9��!�@��q�d"��\�߹-5��@b{�e�cy�U���~,أ�1��9�&jBT=����/�8�mE������L^@g�ܼ�ںD�s��$Td��DfD�'���a��h_A�iؔ/*e���}tI����]@Qxqj`��!�_u>����'|�k+@��N6v(���l��������w�]�z�	����zs!�r�
)�-�H�Mq�y����1��\��%��P�Pd�-������+ґk���u���{��L�$�r�|%U�8��u=F˒*f:[(�6�����g�d-dd��lΖ�:3JOU�|.H�~��3�I���~�V�^U��ԭ�Ӯ��.ί=!�z{P��S4X悘i�QL+��6�V����L˝���r���2>$3&���χE��W΅���raMu�����n"���2�j c�&������-y	�⑶����ޟ�D5�D[��m��N�ܦV�FMf���D�!�G8y�I��'`3R=�����*�H�w�^�ٚ�fAC__R�|LJPQ@��A
#���۔����VZb�)�T�a�$�![�"��f���3�f�ٴ��,��q������m��<��}$VH���о������!�3#��%'O��[����I>�%9Y-�J�@�O.'��|��_k<�X�D]�ځ\k�)�5�K��)��H�52na��:���cԿ����{�%�;1����,^�%BQ�X�V�;����x��R�RJ�1��| ��P/C�s��gJLe#COֵ����K�#U��|藙
$i3��E��+�yᦍ-����(]A�������K��
��s
�';�`��*Jd	gߥ�L�8n ��(ʍ�k�$@	�Z�=�646�/�tS����w7ojZR3�#���e%��ت��4Z��W���Aʱ�@�x�ۛ�d�؁6"�N�I�y���&���E'P���a��+��B�n���[7AF�ʖd@QS�aѬ}PO�y������ȧ_:}�Nx�a�lOZ8]Ĺ	�P��'�1JD�`�b��u�-#�(�������������IX0
=A#R�i�X�p2��Q �����{�5�ˀSEG��g������t��힨crT��|�E�·Ѳf"��
U��q��ә������`ƀ�KIU%�X���8-*o���>V�(N�L�I��E�fN��������B�8D��Tbf�e8!��竀��.7&�@c�3�+L�DU5	p��>ГPU}������W���2h,^�{(Q"��$F�7`�pM�	u�L����ޘ>�K"��n��|*�s	,����`�:3J%���x��@ʒ�Z��9��?���\��a��� V*��CX��K%�q���פ�����Z`��5�Σxb��k���uz5��PT)r���.�_Hu�������F S�4�Hw���b�V���+��b�Y*���Y1F�m�����Hu�T�d�]�S��� �c���?��Ldz����B���=�����~u�KC%�R�
n�e��V9��ڒo����Sj��m�k��*?��x�(���؝��7����O
xj7�����I�dck#S���7@/��y̺s��FI�y �25<.�.;,�D(H�xM�`��|>�%�8�I>~��o��(�0L��*�0u���c7~SZ2�!���D����f������=yjj���y����FB�������ĉ[F~���,=,~�*���I�����3��	��x[��n'+�'b}j�pŇ� �{8����CN�8���j-��\}53� RFi�U��P(~�S:�ˆ,�D(1����/!l�?� �{�XZ�K.�,�4dD���.
W]���������w6*���;�7�����#SP�׬N�,tSJ6�Nf�Lk#��	�)8��f��@�>)��Ԙ1j�Y�#��F�w0=+j�*�\h�+�G?�k�r�!<��N�讠3�������s�����7�ܯ�p�� �����ORk0r��ΰ9��^�O�;}�Z���?)G82�ON�iE ���L��gi�yҶ�T�\!䲅g�z��e|ڞ�2�������4/��w��������G����J�l'�W��2wE`�a_涰c��By���"��'�,ͪb����x,_����
�c���H��G	DM*�Y �����:����ʶ�����y��%��\n��6Д*��Tޥj����0���ʛ�i��2e��4���v�h�Ȝ-?@e��/�����8J����Q�_���y�u�Y��@W��+��(>��kFlfr>�x�|��2��M��Ǳ�zxrA����� � ��7�la8(��.P��_IX��Z����(�J����$�U���)��x���.�u�Q��olu�����&��Sd�o�]�7��:M�V��\�p��X��>��@�73�uh@�۶�����H�~LaFl��
�~Z:-Jc�AҔ:� ^>�]	��[����]��z�or�����3���0G�>�Z"�d�?�Gj>�,�=_{Eണ����D2�*hV�8�ә��v�4M���6��C,h������\��z\]^�~ft�'�B{*h�P!7P"q�W�gp6s3$ J�6�QS)f�[�A�(0bA�j�
j���GA�SGP]?���ǫk���""[o�����lo�6W�;��b_Ɗ��e��o�	�OJ;��(6ė��lb�q�Ø\���(��U�n#P�<����ʥڹ�DA�}�SV�1��n���?bh��F�Z��f���J�<[��ج�t�������J31ft0�3*��i���Mq�3��C:��@3N��ܣ|��Nc��k(�h`6s��j��[���W�^X�ڪ�>��!?�5�y������v�7�3Xa̟U�Lk���*.:���i�2��<���h�Ms!i���f�� �L1������\� ����|�YP>��������������E3��G�s��I����U�5߻��+�^ax�eTi�Qe��gHޥu;�����]-ʐF��luH����If�t�+�D�`���n$1�ey�
��\���}`_�����t*͖w'�_`W@_v�ٻF�(�r^���mi�i�ԟ�|뵲�K<�#��\���-��YWb��'WS��}�u?Z�N�-��℆�F��o��='���"������#�(R7���ɟ���Y��]�d�ҍ��uG��~���\���G���+��^U���_�p�[bْ�R�oc��1oa����x���q�̠�Z���ui� �"��N2��ܕ2������E��`���D�*��h[t�a�'�2����Ѹ�<��&����vU���`0�'�I�z�'�]d�g/�w��qT���	�U���m=���O�q�1ڴ��6�a�(�9MN�X�����o�ڟp۬<�8���~b�T�9��_R<^��h�vC.	l'q���Z���t��le�r7��h-S�ȯW���W����׳9[�=�'(z��[L8���kI�2ւL�%������G�����Fi��_H�{�ߗ]y���V��:.���_�����i��Tg����Dl�^��ߝ��.��@Z	�l�C5IB)�3ߓ�j��B�"�gXV��LA\&Go��?�X��l�D?1r5毦�>T���Oq��2T��_f��7�lހ1��� ����&S�}���Z ��o5U>�hD���j�^��Elp����&���B���'���q���n"5;!�Q�x#t*���2�Tu��=���Y欧��� ����%�9C��M8�|~��Xf�2��L�c��3��8�u98��k�D6��+�?P'-��<����$Mn
�* ��:�%X=v�����c�a���_����D`���ђ��P8��)t��\��t4K���|B�p��Q�!O��ў�o�>'�O��Kr.'4lP8���@�����[����[��3g4B��V���>,~�2�A��4@>ߦ3h�Q-F�-*�<r0�@t�?���vt�ܬ)��R3����/��_o� ��?=|��3r#Pz[��aV�ؿ���NV�7��Ы�ja;�n/�џ8`�#�
J\r��X<�v���2�!8kw>貞�w)/��q-�\����'	|����y��i�ǔ����c��(�Ő����E�[JU��P��>;cVOGF�ZR>R)�S
dsN��a��
|��sy����~������t�`ׇ���f�Q�'PgtRV`��KFs�i�6��7�[� t_E�K+93`IIO^^$QY�q�=��hp)��ERؒ�
�>��J_�:cL	�t��ƀ��OZ�_0ژ�/�7�L�F�N�0t1��{�{&~���d4�v���]A�@{ӟx �?s��a�l��q-�I�Ձ���#.����P����G3_�4
����4iG�i���Җ!�$x�BZ?tP�/$</䶍�� N.2R�2�:�E��T��ӲI��@3$T���8rk쩺bN�
�tI�ǋ~&Z���
�Ҕ73���G��:��qH�H�S{�n;�1'Xդ̅z�9���K)��B'4R��Niֳ�N���r�>!��|�c�0�պ\\0�gA1z�?�k��tV�%^[��x�ɦ�"��Z�>�l�N�Ѫn���Oi`�����M8�<�`.�HTǙ��M�^́8nJ�Q�z���Or:!(������_Г�A��^q���Ѿ�aad�<"��寝0�-��\7�����m��t���(O�I� �w�	��*%7�$%��'�euJ;�Tbxf��а���Ԕx�O�<8����K~��ݷ���������|��yZ���Rb�ǵ�x[gqWji斡�2��a�`}���.5"7��B��
̖�{Ik+�һ��>�'��̎� �n�bnHf
 C3)��kJ}-�ft���#���"��֫�C/ȢrU�[%���Χ]2�c�fW�r�i*f-�w�Q����*u�lS�^��ȯ�ED� �6ϸ���Y7A��րT*`C{����;�|��IQ"Z�{i������`��O:��$r�J5i_S� �@��kP��/��ǖ��+z�.�����H��� �/�`v��(x�����j�S��d�����͏�i��s�>�6��S l�����Li���.��
к�q�D}�_0��Q����9Г�;V����b����g�y�*IJC�/c�(i�ad/�?N��M���3�f�G}��+ ��k�'�A���C+�5������Ep�5?���H�L�f>�@˫�< ����ۅk�_�}U?�37t�`�Q�	a����X� �߃-�xS�t@���:Qey�.>)�t�F!u����nX���*�7�{��/ƕ6i����i�#��peB(&��,�my�y��B6/���n���l�!U�o���f!	�.��*k[��ť���gP���qC��9���	� �/h��\3����يk6��大�l�9\;̢̝�����������9{&m�
���� O�|�_e~�4�8�m����{�Wq�>�x��ׅ�:����µ����
�ل�O*�0�xɯt�Lr�[�� LM�����n����߈>V؃P�9�����nt"E�==T��1O���"���\{=���q�^��-"!G ���aҺ5u���;Rn���zi�U�;��ptcC� UR�ʴy��q�81�L|U�A1�
�gu|�������b�.7-����F�*��P�D\dn�UZ2	�ȳZQv£=J����ЙiߔFk�@�:A�9��{��g�L�_�?�6*�&ѹ¯�\h�֍�X`�_2����
5�3�A��N�����S���X�0����w�W6d�t�s���P1G�^�^��q���C���Gwm�D~�nBS.X����Q!�
��hp̝FR�gT�p�V��c��'W(W�q-���6Ed{��#t� �Y
�Ɠ�US����΄4C�+���v��������ܸh᠐��M��'�xé�M��w^�ǆ8%(�-p���-�۳� bT����\&���3s�d;q��g�kB���e9���Vjm��Mʲ7`|��z��Ln�����ewJe��0}�Č����8*	�J�������X�qy������}WM5y$��b7�� mǏ�J�^�*Аaw?�v0��s�U�İs
��(5j��Ŏ�_��UT ��%����D7�0�C�c��U"2v�ynD���(6��o��蚳��C���َ;M�����@�2	&!L
��3{�K��"�k�y�ODe����wb\% �4�A:)���v�ܰFP�k��g�C�-����'D�(����󍀣�]fS�u��R���U3�S��/A�"3�W5�<�=��"�k�?zB�l�v~���-��IN��HG�����#gq�o�+~���4C(���@��Y5���^�J*Q�[�,&!�I۴���+�����uѧ���������I�s���r#�<��D?#�+[��3��f��9$��O�L �i�?��Æ6��T�]�AtJw�%�	�;��!p���p���ܠ� @��dm�J�x�}�j��L�g��S��^�@ġ�B��n��z����]З�`U���ä���V���&�&t�Ұa�z2D�A/7����G�Cc��5��g��e�Wu�T�s@$�^v综�.��%Ւ�,�@�?"e}�����en�\�P�]I
�#��O!����G{��Z��C�X�fpNqǂ?R��9������-��O	R�����E�L�cm�$ܝtC3噜�Br�����j4Y�o&<jc�mz8�2��ڕ�5�v�!��D)>�����ADxFMaMV�/�گ�4  id]X�o@4�<��_+�JR<b�iߢ�>~B2�m $��P���OE�ot�jHn�� t>��LY�ch��o���YY��Ni{]�.Oo��ls2�̽\mj�%hx�R����࿘*m�w�?��b9�����U��pc����"�3I<���x2=�����t@.n�w�
�����L��1�1A4��r�I�|�W/p�و����&LE9
i�˜�1I�co�p� ��9K�и.n�+g�k��Su��.�^/�`?��jP�d���S�Ƶ8-Up�5P ȏ[B��L�Ϫ7��g��4�<~�5�f�
"��&Sl�	���L�9I��K��:����[���S��y��  �V���X��6����|�P�A�(OX��UM�Ìp�"ZiӻDs��S��2�ư`#n�ƒ���%���+4�wV�uz��'s;�����sf^�dal�9C����am�W֠�=��%'U��g\�5Ku!�T�D��Ճ�@�����{�8T��{��n�#J��L��{�﫲�@�g�3C}���Y�4`��W=DԹ��Y�]-NI�H
�-<�W�
��i->N�O+��VAh�؁"��!Cw\������5*��X;ʺ;0��4pݧS�T�e��0rʋ���tЃ:�UU�	���U�T|�.!��^[L]���ε�����(YW앃+W�HF<�&\�����6dL�Z��!C]zz�̈́��
��ҤE6�����g� �,���]@>�/�)�W=>���%b(�:��X����&����
�[��G m�QӬ���8�����V:3:��&q�|�"-ǃ9=��Y��x�����.TS����滘5
��Q ��J<q�d#�����26�2t�'����I;�UW�9;9�:��O�t���W&=9b6�uR�{�O}��D�j��P�JO��VF�v;��l�wU
v�c��������{�r-X�y~�n���9x��N��_51�v�)	|xK#2�צ�����L+\v+u���i��8�U��>p��ZЎY�ܷ%Wy�ef��ô���_ٺX�p�Y.����tX��D�&L�t�p��yuM;��,�H.O��2������h8=��[T�?#�7l��z�*-UC0;6?u{&?5=[.�J/�'/���ֳ��*ջ��;d���_'?����A�e��EGQ�n�5�M׹�*��������p����(WK���6�(S9"�c������[4��O��~� ����{������*dߥ�BXN�.T���5�=h��I	j�+��֛�ݷqjr��4/�_�B�pMy��q�m;�ʸ�DF�6�I�/y��1$+��6�%�7y}��T�M�av�)���ꊢGͮԐ�JIj����c�VS��p���bn���-��rӴ'1�C���3�Bˎ��Û� ��,}���0et�����^@�!����m�5L�?eF⁹��/ �%�u�ӒE�u����W [���WI��Ѭ�z}%��a�ވ���@i���y1�Lj��a�xkm�<��mɍ,E�;7F��Y�@V�8�V\�����½�]�e������7�r�ߡ.��ve�-_��3���v�#�Ś�ڴH>�#%s;����ٷ���Uz�l�v�U4�w#�G�fd��I�4*��D\��*����(v�`PЪz�N=Oy}�>�Fp�:Oj�;@�? �
�o��U�(�◅ٵc���)W=@��k%�>s��󦺎��ϢX2v�f���	L;	WR�h� ͉O�����25��T�nZ�� ��e9���)�dXA]�	i���w���q��,��jʹ�:���NJ��բ��Fp)1����wW�\&c����G�&�a��n�U>H�����EH���_��ʃ<�,���72��'i��+�#�{|���pc���w�.��|��+xLLO�ҽ��9P��e��k����)��efV����zY�mM
V�#�*�v�*
��!߇��j�6��j�#�"gͪ9���1w����n]P��Xs�Yw.թ��f5�_'��u����n ��(�S4a&�>O"�`l0�L�\�hB�! ����
��n:��!o{�ٓ� ���{U-�{�(��A�^��DĦ�?Z�d'������\r�`j�j$;�̐b��o�σ��ڭ�9}A���4�OceJZ.�����G\ӕ�'�\��k	�4N�X˕tV(�[L�čy:��
�]�SMN�of�įBE��3[ѧxh�Su�r$��YmտAY:�o��lAq=�L��m�_(�^��UF4;�� 8�J����m�>C7�կE�i���5@hD(oL�&ΐ�lC�(�Ӯ\u�5v�Q�����5v��@���ا�3�Ϯ�X���n~�i��o̅���-U];9 ��oy�5O�v�����K�X{(a�3��e�鷍L`��zD���i9-{��^�9���;�c�>?	���fs�3�J~�PL�(�S��l��ϲ.M���mj�Ƣ��-��{J�|�Z��rU����%�"�tME��3�-	F��_
��H?��B4����
��%�{�'�=1]O�	�ZM�	R�67U�4��~fʳ/+ɮ� �V�G)����8J�;9��,�p� P���26�_q3L�Ц���,���-L��9E�h��IX����{770����J����h���1�)��t�'�g[I�;���(����>-��<֧�kNe���u�ں`�����P̏�%{�=��eдL�&Q�/��j!�ť>�ͻ<���D� �BZ����zu�ISh]U�5�E��7Ll���l��J�d���]�LZ9 CZ����aȊ�I�E����t����QZ��!�H.�!vS���D�i�XX��ko�C�	d`0��`օ<��ī%�e|^�k4�N��3�>�ۉpQzao$����gŉ1�!�ТP�4�#��^G2�������rP8o�����l�R��-O�TEd��(BJV�� ����kB���U�ϥ���Tf�w �2����e�����$�&U��6+Б ���~	��/�1�ӊ#��ۻ�K�a�i��{�EX*�ǂ�v6շ�-G\K���r���\g��2��8m�j��H��0���z�!dO�����w��y�ټ��CF����p6� �M� m��b?۞0��>��n~��V��*�p���У�MQ���+~{<���;w���u*�ק��؊��(\�4��3�o�K��X�4�ؼyR�siU�Vs��3�s5�Q���m96#�h���%e;��#W�!/�9��.61_�q|9O9��N�ӓO����X}=/١�>%ʮH��dqXa=4g�OO4eqetV�D/}%��_��os���p L C	P/Ȟˠ�յ0(,Os�<���Y�sso�h�asB����6𞢴�`�.�.���?�dΌ��6���h���K+����d+;��_e�tnT���+�v"2.J��Aj�د���B<��(`;|]�'=�B^�ׁ=̇��x�Ǘ�5�#����D��Ś HO�1r�{���!`��vS�9��%��{�}��Rf�L֔m��p)|�����5�;�Y/���;���m�z�>�d�p% m�����(�wb�D�ص#Z��NaW7^%�,e�� {U�����|��Ȟ/�0�K�T`[���wI5ߍo����dy�Vb$}��}����֍�C5��&UN򥰫����y������)�'"�N���. ��@�Q��.|6�
(ˍ��[z5yuH�К@�-i��W3a� ?�2�u�ƅU�e��;�5�g!a�
��yn�2�n[XBf�ܖ`����%0��z8:Hێ;����5�ɟ:�V֩f�?-�ќi_5��6��$�+��)����jC0�{��Qr�SI����=_���8�P�>���9h�b+AaOV��?���`�������*u؞�G'�ف ��
�V_R��x���6��k~�`d�X�Y��>��Ä�	G��g��E�OH��=��G�r`O
Z`�Ɖ��"R��4{�� ��_�6���~1S��eB/���#Х������P�F�}�k���Yɥܞ��Bf�lO��YE�H�����ÊN�:��>�F�Y�(����d�ja_�}
�d�&�W|W4�C����f�L���IŴ�����Զ<AVմF����G�"S��kt�NT/���L�n>1Z�uT�Y���9���X���2��"se���}�Q}��k�t��Wa)�i���'h�F+;����x����i�5����![���Z��2������Y���e�{eD��ޅ�LΌ�~����f���}IԦ��Mh�z��a#ة5���0"+ѻ�"%�i�۲;�=�z^嵅��0��,Ǔ�~���Lk(��U[)��AL�ˉ�,A���;,���0�b�N�}B~O
}�ُ�����`n%�#�)����α.�p�K���d�h��5WJ��U�Zy�r�|�r��������5�F�k�.��Ǉ��čd�W^ 6���U�Nۨ׫<������A��y�TPF�>B����w���)>���H*>�3~&�T$r?8���tS�%��qw�WZ�9���g��v�[5v�D֜H;;��"r���'�F%k\5�32���`�/l�7�1�cᑽ���������ш�?e3���y��;P�e���[��7�C�_�2���~�&�ϩ�N(K+/B�u���@���5�R*WȮ�)�`�8]��m�ݐ?�)����fv^��ɠ��E�x��������?Df�p�t�z%����֋�`�JO�?���l�7ё��P3)IR�R�@]��2�,u��$�q"K�a����_�o��;;4N�ecP�?$�C�@��^AHI���kzOo	�%��h`�܇�õ���~`�TDB��3ZFO+F[|�=_����ky�ɚ�F��
�Z6B%�����3��,���Pk`	g��H87�Y.���3c��O��D�i��r�Qg����-�q3b�������u��7��q��z���L4��c�3����B���������?E��㴧J���x{�骩)(��o���C�%��'Ę�ӇL�+˵p�a`�E� E���nۿ�r�� ?�ƫy�Dh��f��{�����GZ�m~q�r�1�O٩��o�1�r���RPu���HQ%C�A�:H9���â>2r�e�������\�aYV�/�W��O��z��x�/�*?�!�!b��oN��$�}l���=� ��Q��Lw���E�j�W�g����.��+盝}&C�9���%�_��{�D���V2ɵ2p)�yv���o͸��~�:�O���:�+6�� ��)�Y��kE���.h��ݲ�N\���M�E��>��[ q��Y�v����;�p,�����%��Fs?Fe��8[�9�x����S��{��%4Nh�C���M`��鄀F#���ݵ���nP�ۃ-�Ñ��l�*U6��dZaD1�����T��`}v�Dc3��`!���zW��u��=N|
#p��/[� ��0�Es�=HA����}��<�>C=I	��`�gL_�Q��[M�H�x�4��)��"�-�o�+�97fbk-��7	U��D�*l�ѳT+*b�~M��z�\��^�Y�鄬V��gt�(��6�
��#�w�ؘט-��^�KeQWa��|zJ�M����
o����c��alȰD�9�"$6�����́ht�wYf��=�h�#))}Ѥ@l�_�vs�aϕ=-e�E�J	gZ,r�B��D�Rp�:0�[.��PAۅs����������b�� �ѹ
�~k#0+&y�)}��K$*�;��iq,"aٗ`�k�!(&��p�a��sˍ���r8֧�3�������KW#-v�Y��y��b6�gZ���r�0��G\@�Q/
�&Ya�I]��U�����X�T��5hC~����;��b�"@V}R�ك����!�G���ui
4���F��|�p�N����Ħ���,����u��v��Cծ���[���m�ڶ�Ƞ���ᑴ���q��,W�Ֆc�tg��S̽��5�����",;
��3�E�%�v[wuU������l � ���ß8�c'���шY�d�3�nv�~��k܇D%�}�M��=���ޢ�ߡ/��/}�:A`�.��!}�������ǵ�>��x�8aS��(�������F[��+(�h���[W���Lz�*�H�n�ʵ6g��u���w�k�9���T\S/��m=P�M�,s��,b]���}�_��vt1|iF�O�w�R���s��(�G�Q;��ϳ�#�5)��]���C��s�ӳ�gL��D;�+��%;�*�@p�?0�o��zt%��/L�i���6z%a�= �ܩ׾ye,-r ?�ɅM��0F��K��S��g�:�Z����MN�O~���A�q���-w�E�����*�Meb�ѵ�Y��t4Yg�#x�vG��՝OPn�\w��&�D|Ǻ�s5�ָ#�d�(�X�I�;ö��۫���Q��H�X='N~�@�+�e�k�vP�A�B�����E�8>�$Ғ�ך�r�} ��T~��OZ�  ��gQm���5���Y�5��]�MA������RWmG|C��c����w��~!�X�C��2�7�n��.���z�^p�YA���H���ȉ�F���s��{�g�Rޑ 4+?�>�B\����gQ���Qo/���-��KM�B���>�����1C��K�\�ӊV͚�h\t0v�W�ܘ�էJB��~i.�i��D�������f$�φ9SZ9"����Uw�F���\���'}\`�pA�ư\�Ǣd	j3��c5�ᕁ ���A�����J�Q ���F�g����ǚ0���m� f�����GC���2F��n��r?:ǚ��81�#�Qpc�h5�	�fA�7"�`�M�xф�7�M��6HkE�#��܁b�BjoT�3��E�p�ԓ��It����Ӆ�'�=O,,��A��*Ѩv�Z;4�8����*�z���;4����i��C�{�������bDŘDl�ƫH���u�D�!����D?�i���=�d��C@�ڎ�@kt����[^B��xgn�y�uCkwtd���G �#;m����0%���S�s��#�t*80-�h@��7��9���5��K�o �0cț����/�L� ��Z|�lV;���l�T$�9��:���2�w4���3t-����
���v��w󛯖�����2Rο=����x�c�`Q]X�0>�_�gT�g����*�3�-u����\cO��Q�����@,�HѵU����{Ǵѹ(H6[>eR��ȓT"��aN��ga�e%W�d
���z'Rz��:m�>�V�qR����1Qu��D:��JÀuۯ��d*�y����{���xx$��ŏ�akt��FD������a�<��|�c��C<B��i��}���)&3t�_(.��������#ܳ�� �� �<;��Pgp���x��/�[��-�9��}$n��3��|5����y�@�"U�a��LJ˵�Y��~�ls+�ysἦ�.���S�!������-c���r���t�yΉ����p�����3�e�B�Ku<�_��j4`�h�ݳ*�%���h�Z�d�͚�b�Л�[	%�0.�!}���/F����S��s(��ח�eCo�m��|��fj*8~8Tt��r;ϪSE��R�]V-��@?1/�6�����y�]	���_ �<\p��6�c��.�7xPe�hz�j���ԃ�2�Bo{���N��\���)��t�p'~7�_�$d�ɭP����ܐ�������O�{v< M��7yF��Ģ�T\���'\G@�}������tN� j-��Gk~,��@L�Q� �� ��!�	��;ܦ�f�lT��/)�� ,!5ر0~��
�o�Y�H�͑brE@�"�Mm>'�i���Y��p�} j���92t���w#Ї�/�8�n��l8ƴŌ�Kj5VaQ���H����B����D��Q�&v}9/�F����<��/�Z��p��{�x��`a6߉�2���3j�۰�+7Dϧo�}`��G~�|;8�(�p�?�z��\�X/5�ݦ�J�G��P�ˡ���� �D�p��+���r%oqR�{���h`f��1^��Qj�Șu�m�tf�|�"e��)V
Dܠ;�)�&G�iq�kY�){� � G'�;?B�<S0�h�e��]��*������̶Dp%ܩs�G�'`�n�^Z�޺@�x7E��,C�����G��ȫ���D8� (1����V�+�11}���΃�e�E�۪X��S��qIh��!�>�I7X*����Zc�A�lET���!��?/9��K���#��t�^m��eH�jZ�c�[�/ŗ��r����Y�_,�x��F�ZbH!�\���l��(U����:$�L��[���nsp�� �MS���8q_B�9�Hl?O��W�����$�G���6|IͻJq=����w=��b6�mJE"��\��M�� ���,i>F88!��ɹ�ß`� �tpj�k{�ȃD/�t���SAm����6l>T;	˂��Z�3v�h�oj��ܟ: ��z���4�8�)�f���C�5��G�H;���PQ� ��4G�����m4��Q�����t���3�K��!�=]�#5��}i[K��;���'�!�Թk^�-Q�m��m1��e����G{�/)l��ʨ5���4;X�P�F�^�
5-ܭ�bGe i���=j��1�( ����/�}�~%O�[ئ��@��a��ԤK�N�	�I�/9��Hє8[L�����m݂&��6&��0D�4H��<���l+�e�&o�$�|rw�L��+aQ�����h����K��xE:�~�NU�H�l!ߠ!�����(5<������h���A�y+�α&�M�G�
f���'S��c��a�Dƣs�����J��q�4�����n�S��u���S:L鞬[MԌ@��&L؊Z��,l�80 ?�H9J����������ĮZ���r�g^ε���p� ��������ٌ-����4Y�Z�B����C��K��%wT����h�^L�:cx:���I�_�]�a#��������Q�t��8�-˩JV�}h����3|6s�jp�cv}�-ɿ)��JP (���YlC�>���m215C.��&����̜�k}�5��Cd/1����!��!��c���}����A�o��� ���)@�z�]��=��Bc�o�*b��ꅛP���=�4W��(׀�W{/�A��;d���� ���^
���t�r^U?�p������qf^,W�Jp�Q�i����0H��#	`��V�f��΢J�E�����TD�c�B^��D/aӋ�0M?���Q�L�[�(˽��6��'�{j�~�B$�A=K��9���o�B��� }A���0������	��,M���F�f6�6�O�u�x�����ޭ�#e�7��+8>Aํ�1#���G7B�=�_S���]�Đ1��zĖ�%��� �O�s�ޓ�3���oi�#���2鏎FX�V93'�ʢЛ��+t�@�}�x�_P;dt��E�3�ңq;�T�|�CcVJ�^�K�Ծ�'e�%r�����5�]_ٴ[���邆����Y�'�)h�&%��i����J��j
��〪T�^�x�'g?���쓹]��i)���.����#s�m�߷���9���R�'�w	vMHU��2R���W��6���(���FN�ēeQTd��D`0Ȍ�C�*����q�p� "��PM06,u�ɚӱ ��2��JQ,K�pFj!�%B����άlP~�Z;�r���XaF�Z�AR�궉ϛv� �{��v���C�7�~;�w^���{H��	9�\����?5�ɪ�e.�)�u>�����g�9T�'�o�K������U�@��fN5b�v�94�t���At���s����qx0.����I�4�gIH���fj�=Ἵ�N��t����Ɛ"K�6PC�ҧ߸$0���G��혆��
�`�����A|wtN�mbC�UYƳ��
}O�z萖d��O��K%--t�"��j>�
��1Qb�y��p���/`9R����&�e�u������,�\���
�~4�	��x
�[حM:i� B.�0m��-u
q:D��ew�l��8/�9`J�|g#�7���*bm���)=~���>�����M;�꠿�:���Ձ��첤5��> Dڄ�bv\���h�ta�ku�`�ڃ�O�i&���E���#0�K�@@�'߱���NfH�7&�iMT~����1���P� Ϝ/4��Ƀ�I��_�QϑVgƪ���M�_T�DQ���L%~�a[L���۰�
g�iNg)r�'#�_�5vT�okp ݑЮ}��9|��4�#Lݩu]���J�q��O�?ޟ\�/uR�@/�sx�f0���3ݝ���b��e�״n�[r�<�O�GOc0�R��;�)���~4$�"��&�!��3m�Mz�@@oP!}b���	~_.�uE����3�`Bnh���{�ų(k��R	S:����л���\z�>���ۖzܢ��U����ݫ����5a`%SW�a�g���^& ԣ�\���;�wn�܁}ݟQ�Yó1���&�q�>|V�
6Q�|[? H,3�*㛙�ah�����V�*�JBDRr����/�!Z�Y�2m���u���%��{(*�pdE	\��Ty�0�^�+��� �w�6駃�Ǜ��m��BQm��z��[���),[�[8n
)7e-F�� �+8Ã��2BgVQ�z'VLdV�V�fd��FL�ʫI��|LJnL���Ÿ̓bI��+Vo��$?|����+����6���m����('c�:5]�;�u3��j���#�WN��'�eA`���L��'�R��S��.<q�2լ�������𿡕��I;���T����J��=W�.�d���r�EAD	�RK� 5ڌ��Z?�N�'��6Y�1�qgG�r��e���%��{qw���j'�[hi�;Ö�m��y�Dn�H��<*�%.��b��8�7�P����_F7cx`?ꅵ����uL�}5��P�?��>9~$�N�����z[����J��U�cZ���s�xQ�8҆��(��R�Ꞟs�4���w�s(�>��@���M�C�+���ɜ=*���S�\�J,ph��XC�۪'V!>Mi^T+}����̔.u�wuY���L�ܫ+M�E�ʷ�cmʛb�ve蘸|�&�H@^\O#��.�@CL�� �D��\��4�A�q�S�u�m[2�
����1ZM�.�m�^	�ۧ΂��C'Y� g�L�wm �l�ǰ���ZJ���	�K�C�/Wz ���aD��U�$�ZIa�8Z��`�O�b1b�ζx!L��1�����8���g���_�eG�='BmL��\o$�&{�@����|�یATa5j��,��n.�Fuo���˹S(�
覠#���<-8UvQ����b�̀/���F�H���>._���鬩��.V0(��f�N��]eX��٬����t�ά�`��� �|��Y����H���]��j`����vN�,j|���Q[� ��:W]�2E��Yb��	+��@ouq�'<�����-RG�\�<jzy���z�F��$��i���"ݜ�E��~�'�� ��rfŜT������,������	�O�,*��A8~Js~�֣N�*�\me�w>��0�7�8���yW:I~Ǥ^Te���#oE7R�9q�^$��v���(+	���A[�����!Q���t��O=+��޳��V��^��zm4u�o���ξ��s�u�֡md�-��+�JaU�p��2��/O��+驆-+��L�=bu��D<ѦQ�b X�pws`�R���s��U�&	�a8ۍ�4C\TJ�S.��Ӑ��
�!��� 
�.�D�o�MX_��o��A�)��6�e:�T�~�;��i\O7;��)ѿD�&6�a�8�у�zq������Wl������ʤ�-�' Oa
6��Ǯ4:?���kW�rdj���)�v�8�h< ֊bݐ����.�Q]~˽8=C�f��9�_BmKq_Ei*�7��8o�?l�&ؐ�s�
�ER����{MŚ�}��.�a�pS}��^koU�?�ǔ��ց!Jq��@�V�x�K�'08;(��i}a��`�9� "B�Un���uШ��٠=y�uH�2LǺ©n:O�J�(&�����c,(O��R�;����j�VY"�P�Vid�Q��ٔG�b��Ъ�gsj��;��×��E�a� ���:򍨶����Z�OHU�m⩭h"[��J�Ttd���ߩvr�I����@L�~ui��z}��$p䒝�i_��u�0m�ǳO��~���5X%��^K+i�>rȺ~P/�����A�yo>[b�O"��4�u��q�䪚���w�wk���n��~�ġ���R�ėZx�+��ZY�e�ę���ҒyW/�AX��$�Ӧ��e���Y�g�tȲ��]���~�SEg�;Vw'6���O_��bi�4.T���k��j`
�^�gw���_"A�>��Cp����Ɩ��ͬQIW��=�7}����Yw�@����ԩr!>�y�wg�T���\�Uk��2`3 �s�h��� 2-��$u�Ǵ��I��]W�̰=��F��[B"���;�� ���-�/S��.OL��D(Y��x���׻>1�-���d!�#��\���/�3yώY��b-_[ �9e�Y9�ן������)m^�:�Т�}m؀�����dl�`3-d	��z�ǉ��Y�#X�v�\�����Jb�k/4d�Z6�oز;\BuːZP��^x���V$��`�rC�"����^���'+`��^��
q�� *3a�1�9���� ��`f�ݹh�ᲀ���|��c�(�P�������#մԫ�j�+��=�W�6g]Y�6�����+�����ӱ;{D�gŹs���;����k��u��WyF�x�4��0?/kl f*�U��`��g�i,[�z'�(��b �t#G�~H˻*N�`�� ���l?]��RΡ�ɱ�F@AX�S��a�c�eF�ϫ��V�o_Z �s�����7"�@T��h�³Dl�7����d�p�.�c��&�`�gՅa�3j��X&�M`�'��X�#E&���M�1�c�^��⼥a�������l�u��F˭0���l�@���&�n�����!�c�-L��=�˷طLQ@��R�hW�-����/��%c$��Q�r�6
+���^QC�GY�1�ټ��@��1��N�^Y�`���UfVA�F��|VJ�*�?_��%C�U;:�������A��J���
�q�tOu�Q�1�M̤����c���g���^�.q~ez�yW�b������>Y(*É�J?�?:7��[N��V��9� �_���]�If��ez:� I�7��z�n�+�s[�4��o���"�?]I�[z[җ����\;=_�d
�('���U�9F�@U$�W$�~��˧-�34����Qnn��(V����;�a/]�4���Eϧ����\<��Ce���]+��j!@8^   ��j�a����&�Lؓ�� ��dJ�͈ŕ�*�Cim:���]+/C0leS�c��a�]fȠwY�Me�Y�sĜ�o�4O�G�t:O�b>>@��d������`�@��Q�����GG�D�l��#���c�^�Ыj�H+ }`�}̨�Fd��4�n ���r���LG�_�#Q�Й[��O���j$ �
��M�R�"����ĸ1���'>�d��=��,���/ -헳d��o@�(8��"���G�aA=�H�黟4T�h& I�6�	�x��P��i��N��{P�y�������D��������?���R�#\p���C��4zX�xd��!OP���x�%�8�V�w�%����G4T���re ���}�J�**�@��� ���	�(�~������P�+Q�� 0v~�3�+� ��挕>���B�"�]s�}3��W�4��J��Σ"B챸��ܚm��q���M��{nQtG�Z��$� -R��O����r�8��8D3s�(��B��ȶ�q�����~�G�źI��h����nu�����[5J<��!��:�c��	�YR���Ď��e�}IR���7|@�LJة���ޖy��m�r$�+�:o�icnM�̀J�s��-�ۼ���B��R�yĒg���X��Y�$��T��K�y@��O���If�p�� �S�2��z��zq�&����=q����=�!�C �DtkF膺�0q&!0V�w�ׅ�̘�V6a1��?�����������ZRoe�JnN�z.G�S`��Ͼ�G�'���y�>����h�u@��C���\`o����l����u��l�}aެp�S~x����9��@trX��Up[������~M���n\ ) �B �f�S[���2#����ﷴp{�����!h�cԙ���O��IXI�&N"�E�_��c��=�#�J-i+Ix�j�G�z���x�d������)BP�8�`�+S8�����N_p�-��C�l�㮌U�s ��T�,�7�"�;X���ƳI�F�}������b��j�O���(ZR��
=�1����Yh�&a���,;h���GR�W��ϐ��Q��Rk�3Nm+ O Kϔ��k׮R��k.���O�s�,a�@m*1PK*���lc(J`鹿��aU{��c��;�A��Me}�W6��?�iXKQ����?QS�M�A��K��m�|��]�ݥ�̐I���'���6����~�}����)�	P��5 !�.3�R1XF�����4�(3+��Ќ�e*,wW.0:U^�2'Lu�JVw��P"��鉋R߇�`kr(jZN$�{�� ڂ1��+�n�k4~��%�ae8ג�a��,����_9�z[y�&�!����zQ��my��~:��Pj)�tl|��Z��G&�n��U��^T�rǱ;�H1���CЭ����T'��L;ݳ³n ���G>!�Vaӈ]�d����k���~�d��<	NB�iO�$���Z���}����^Ҽ�]���xvf}閵���4�i���«�A~
�O�*	��?�`����3uM�bc�Ao�8�̑}���n�K��k鹧���]��|���+���	�:���X,�M���~E���9��4&K�GqÚ��:������ʑ�U�?���5.I�rY���9·dƚcg뇱L�|���!%nO�/�gV��W��㖨vik�Y���kң��]��˛QO�N+@eI���1fC�.��G��عzh5�����Y�����9�w>�c���5N.���{�^o����䖲�e��+�dr�J��� {�Q�o����K���+��fo����D�O�r����]529�i�G�|�#V}A�|��i#�q�j�"ֻ��v~�E?V|��ϳ����\Y���"���{Y!J�^EH�d�����a1��s}�� &Sݽ���]vV`�vڗ�(	6��"r��7�\�FX���Jr�|/��[�wF��]p�W,6��IRs9F^��W]�^��ٟe��ǽ6r���m9ODyIOҝ�)F��ps�ε ,�=w�������U�Q�����C���〮re�N�YZB���J�v��OT�C<A�뱉�
 |��~J�#�rIi��xK&Y�8��л7�i�χ��sn�5_�;	r�Kw,оl(;w�2ig��YW�U�Ĕ�$2�6*�(�@I��X��0	�����,��"��(�C�Z=�2��G`o��Q]=�PMm&�C���9�2��Z(���T�C�p�ȧ������rN=���(+f�4��!�^�+m� �7��u�l���Vd�"eg��zF�m�v���q��xk7u܀� �y)��᝿�HO��m��̤~QB�r��G���p>4!:�r&����J��	����T�L����$ձy��\1��b�{w��
Av�#�<W�R�jz��
��u� ��?��̋���5;�Ru���!Ϗ*�o@-����k�C�L���8z
г�$x5ɀ.r��K³M�n�;$��'��`�2ltV$���4Vө���8�����:S��p�µ>~�/T��i��9�6)�
M��ZH�]J�q�5�}?q������$�喯�ٛ�J�e���ם?&Y})�Vϭ!�v%�{]�B�h
B�����"]��83j��td���0k�t=f�6�s��|�ҟ�k�D�p��r�P)�xyΊ5�YL�b��㗗O����EtѬ�VH+m��kj�J���9�LfCԌ���U��R�~�5�qʭs�&�[PGo�/nࢿ"(��4*�W��V4�\+:�α'��Z�CP��D�Lr�k�ｹ�;�q�6��j�g�~��ۏҫ�W�쌁�I��d��2�5`{�qꛊBȠ�ru��&t�jWR������ܮК"q��'/|�[6�$s��o���6����mh�F��OY҆5��9j"��w��y%�#�e��F�I>�p+�(]�������`%�� p�pq��װG���y�p����t��\��kY �}:w�����S@���&�*s<�Nx��(�7�s&:�9�@|��/%�`�t�n���A�«
S� Ib^�W���P2�I;_�����-;V�s+R0*Ҝ5b��i�SY~C�Q/��Y��j`��P��Y�"c<���ؔ"B��7���~�!���&Q�������c��d߈�,�b�1�FnǽoT4��_�")`u�2g�6wX��1d%������G�]��)�nТw
��,*������p@����V��_��VM��2��À��i�7�N^�A=��4�o!M���bN�8jHhI.Y(]>�z}x�D�x���x͟oc ƨ)�tx����ԩ�̆�&�W�"�FM�n?�Hzs�w��58 �vz7Ir��.�{Zm��1����{7�D�3��t�h�Iⓤ����tQ1r������hWO��Sn�(�ع�&�
�jʳhn~�_�{D�s�γ�Z��I��mT� D�rp�ż��eMQ��~��dU���ҏ���6�_�����^F2�V�nx9QBX�n�#�� ׿�B
^hܧX�ZaA�t��x2�dŇ`�&�W>�H����Ӽ��0V쉝� W�eK&}*me<Ű`M�j���ǩ+�1�"Sxğ4M�O��z	8����K��M�`p����F�"}���9����.�������@0�1�V�VJ��n'{f[q�5Ё�<km�A�� �`��|]7��y�%��HR��$A�<�iq������Rnq	&�����/͑��Wv�0l�qqs�A�x��j���9�=����==�{�k�ƀ�m~��s
I���T��N���>��{��hJ�Y�q�`E�r��u)Z]�-��Jw8��p39 ~	�=�{��hy&i~rԯ�����"K�)p�9��Jp7�ׅ�*G��67,Q!�R[u��*��O�6<�������-5/|��44��1}\�6#��	S�;��C�?��^M�o��::蠟�������{"E�]�l��e_#,zʂ�aXpp��F�\1��Z>s�����嬞:Q� ?��>��/����7Vsۓ�л���(��/�	;�?O�%�<�A̚��dv��pUʅ������WÉ_��y���Ӈ+b�(|(���a	1X�R��;%��4���7$̊���Sκ��0��7�ξb0��z���3�db��)}r��р�[��e/�<k�䇢Q��~�S~�Ђ+�[�# &�8�u��x�O)!/�0�
d6:a��umxĎ4sC����pRu)��Q�6���@Y����=�g�u��o'-F�j"N'l����g���T���)T��X�\���T�!�7f{7c�d<)�!D�<1��d�d�]�om�'�鍉֨� 9ۺ#�MaH{DV�ƽ�k���/����uPi�����&BC��ȊN�Y�2���~Y����A/��� �X��<v�����1�TI�{f�A�j��9^��GG�o㼫�s������'�]�T_~���6e[+��I喽�S/�b���)X"��㮏���%3�+�Z�e���8��
o_GX�`��j��Qv��*�j�����w_���p��f�O$���~�/^�V���#�mv�|��*�]�}��Hp���^1�r	M�DB��Er�"�޳7�`#�v2-rA*��`�K��S�1��w��_�����
Jz5��Մ��DV˴�k�ɫ���d�O��j�W��%	�
U��A�&3T��1����`?p���~�"@�A�˫u.'=�d>�' ��ب�����c�=0���0������W��@؈�'RF�ᰁ�ui�)/�R��F3	-x4x�݅I�TK�Kbʋ�	tv���W�+��7{�ƒ�t��":tX�d,��%���e�b�rV*蔺)t�Q�ON#��lf��UPY���*��B�$�nZ�����
,�zO➖y,��A\�������lR��n"�!7e$^���\l�8ܒ�C��gK�ʦ��:~iVC�F{�#L|t�l
���j;?k���]�H����#.�&��h3���+f)3��k�����WI�#j���#>�<�BŐ��a��m�������/��	f�a?.a�||3}/�D�i�u�Ok�^����nC�(� 1r �f~��Q�U|��]5��K�fsj�#f�`[���0>ULd�����n�u���M~�hJ���܀��}3'E@LQ��ev'��6{�����v�a�.������N�q��
(I��p�S� }/+�%�|A�4>�xS_}���5 �l���]2�V�����-�6S�5\�+&�O^Ɨ
�.a�ĝ��,��PO�!'�r����4t��4P6�y` ���i�{�3�"M�G�^��F��dڟ���nll�`5O��jp�~T˽�m��;~طĮ���;h~�َ��mC�i���A,��Q����;�m�;PU�?�K�s�'R:"6��7߫iv���c J۴�|&�FhU`WE���1-�`�Sd���0��o�Ͷ"-J��2��2#��� f�F�c<���!��$9Q�% ���aIy@f*���묏��	�=�3輵���&yfS��H�^%�����d;�';���j@���a�L<�K$����e��s��\ۋ;�\k���`�u��wz��!��`����m����7F����u�,x�^�PC7��P)��x�tp�Qd�pg�oF�`�-��_m�y�?�pӉ>o�"�A	y�|�8_��,>� �_��ɀ�R�����ɶ����k����(��P[#[�7�[9�#��o��<E�Ĵ��J��
O<����i���s�x���>�¡$��X��p�k��˃��ZEb�m�w�r�Fb����s-�pa1��v"HAp�`��B�I��+��v��!<x�<d�a�$*�ք��#�=�x�M�����j>fV�6;��Ξ�҄�%q]lwƙn��ި��鮔�����ugc�f$�-�.?&E�Cdnbo��PX�֮��wHb�b�0����l�M���	7a]�]56<�^�%.]T�<��UtWC7K���y%� 8�nLN�(�� �.�m��y��H��d"�yXf�5���5��I1&a2��מ{�����	�����W����fbǝ2h&���r1욬��|>��	������=x�v_�0�gT{�g�	b������5�C6�OB̖Ʀ|�ɸ/a%[�EK�W�T��X�@ưh[��Ӫ�8#��b���[h)��n���EN�_y�Rx���[h���U`I�;���푧@ꁨ����-Z3� ��?,�]���-#�K�<;�[/T)��y�%�0�� ��������!4q�������c��5�o%�)Ӎ�nQ�e~��s�]�o�j��4`@��$S��gR��,���6�o8#�ӑ��r�G���J��f}�D��s#��BE��2#G(�L)� !8�dD���x��f^���g�tU�l��v:ᱹ�I�<�e��t#�:���9¿=��N�e������y�<��_�V;@�QDi�9�7�"Y��h��pʫnQ<D��,!����6���ں�/�G޴��6���5������%�� � ��ﵥ��A����o�m�)չ&�^�Y��Lݎ�����|e�1;q?�x_�mN�^�
�Ȼhq�zN�c|�E[�jBO��,l��B�P�[����X�t��yɺL�-�/��T�{�Ѽ�D�\ �{."$�nm�o�ĉ��2/�,@�b��N�Í�A���|��5澙0`���תs�wGSm���1'i�x���	7�����Z��M�7N��V�CWt���a�$��[�D�����E��Dx�Iˢ����PE��Շb�_�;"�o5��n�����W�2�N���9�-M���>��ڊzǷFo�X}F���y=M���_<���g�Aq��Z]`�Q�"��qV��+E�^l.Q�".�-���	\Q�١��|eYy�(6�<�~��q��hUK�O�b*�^=9���l���5�ܣBy�D)�~y���@Pb�=ٖn��J�%7�-љ_!.{��$�Y�T��X-/�?Y�6�6�
�������k	�F�9`䆁aF�ȑ�6'���<�(E�R�-�%�<�Up���540��[��p�ȑޮ �;.�)-���U�N^/${�L)�Fdy�}���ם;G�ߖ��*�E.+�Rҍ�şn�g���w��&��%r�$O͚	F�2�o�]zY��V�����NB���?���Y"��?��}�%<\єe:��g��v���)�f�d[������|�����ai A�[��FL����d�5c��if g�.!�!i��'�?$�+G�O�=y?U���sB���%̫&dPڿ�&��H���
��h0_�fH�J������}���=�"]-;�5��"�1�:���ڱ(�_��ͩ���ٽ�p
q}�G�k�wK��BO�c�����+ݯq�'�鿲t��%eAG����R�0#�݄��7y��"���٢���r����Ap���O+��cv�'�piE�6���ʭUu��Ʊ�hY�6O��h|+ז��g�� d��|\2}�~n�"N��q��ڂ<)��������A/�+�u��ae���d��sc��Hl��4���dɤ��~�G2i/.�w�}�N�ՇǕ��!G�����h�Q�w��w�\��oE(H[t"^�M��l��LWY���9`�V)%�{V��FN9'��585�]� u�vv��@;����ЂxAD�csr*�t4FX�Z���- ���sm��^�>ø!e�L�{|��e�8����J��U¨��o�7�ۑ�a�e���S5��'�'#`*�č9f�t����ɍ����۴㕱 񱣀Vn���J�g��Պ��P����Ϸ 8V��y�$�G���5��;8k<Y�cN���G8�X	ى�d���ܗ��M���@�٤���<�@Sk�}�j��$���qU�&�B�$.�E+.��*�8��1�_��y�1ã�&�P�I �*\�-�=�Zp�����G�с� ^�mEG�&��I�-����N���E�z��^�5fѮ���G����7m�͑�T��>��UĤ֡@���)�)�~l~�4�d�(�>5��^�0�!�J�RN���D&.��F&�n�4�Ĭ���!����Z�.a>Z�&�˱0��9���4�%�B�,0����ؤCISK<�Zޗ_����JX�V����z�O�̸2��D�� �#hc�y����a�#�Fuc�0�0 7b�6��������h�!T��T�������-&a�$��������=r2��v�0K�{eQØN&	��%+ Q�,,�@<�)� ���v�����T��V۔��n���������e����(��n�zU��z������ɫ��Ö��!�mw�+� S��=�R�Nv�E2�a�%�14m�J���S�di������ЗC/���hK�n����� ��'K-f�}g�<Ow�H�/t�)�;���~��.Kzp�RWnuxӳ�y���1oP�/���>_�g*��u�뮘i��Q�g��P��5-���mw��3���p�]卜�_-$��5�\Ö��$�1�p=jb3ڌ��$��r
|�����k��y���7�����?��$f"a�
�C�'��9/f�k|ҫ����fF�_v��1�ݹ�=��wߓ��|c�[NkXߊ��O �[x��!�U'�#��\φ޽8]V.��e����&�WK5io�<U>p2��I�	��dX��-�V �����tc�
Û݁�����nT��[���H�utԘ<�1@��5!�0i�q�q�~��@�sHT�hh���#�x�)�^�����D��><�dpw�l����V�s3��K3=�m��\�Q�Y#$#�$mj��8�B/��i�P��ѼV�Ӻ�`�^��-��MMkm�5 փM��lR�Q����P��+/�Y�#�x�
s�$�6��ʝ�"M�m����x�-�x*�du7ȵz�~g� ��́�����9�
{\^$!"h�|���B�:N�4�w�x�e��� g���{r�T<��ǧ(f�g⿝u�'�߿���E�J4�9��� �w�D�Q߮>R�}?	狿Y|9������%HGsC�T�Jǂ������t-"2�6�j�ޓ�U�|mU�F;˕�݃oJ�LfC7���Q_��ej��T.g�(�;�13��9&�B��Hq�S!SL �@�3���ڮ���b�<nہ,P����N뀒�U�5x�07͂Ϯ�ޱ��
t�H��x>A5�b�{�!h��+��<�T�$ș�dr0})t���$5��`XM_g��k�̄N��|�O�P{���K�޲�ܢxн��$E�sN{nE��&`�/�eD��*���������@�����ۍ�}��ڟ���,�|C�[]�F��C�	�Y@���^���d4�9�;Kk^�Y�#�(q�"A=9".�r��֘���=�^�b��G�u�4��+)'�b��g�y�����m߂�j�����Ρ߽c?T
�I}m?���QkN��t�8� �!ބ'>V���+��ۭ	N�GV�	���W��*�:�xA�mJ{�l�)�%2�Ku-ۀV�ĚƵ�>y��a҅���R�Y��:n��������ߓ�Ref0�[���{{nX,b����Шd8\�7�g�jIQ�/��:�r��;��,�Ҿ
��`�H��!���2S�B6�iC�ĕ=��g�j�����CX�{�T�� ��l���s�Hў]y���ز��,���a^a�N4�-	#~gZLAe!2+�C�v�T=�iᑒ�� V��z�n1�'����H���A��X)vm��I=c�����]qB��ߢr�_�'�G�3Ҷ�ǖ\�sY����Q_�NJ�Z�f����x��i��E}d�E���0��+����U�r��I�g����*mIi�����}� hв�hs�����(�Ȧ�LZ�af���U��<j�xG�w�;�+��(����5H���{��h'ၹ��{���H��i&~�I�7���~�3�����DՄ�ϛ:�*�T	�o��Y���H�Ǯ\�O�L��!b�����}�Hkl����6���#��m�x�AIs���]�S��M���{���,�(N��]t����p0%����]�����T��ͫ�^���-��_�$Wh�Y�n�b�V(�J�zrɆp[2�@�=cCt6[�-Wp��2�
SF�
,�+�����B8ח@B�<�"#�����:���Q����� �;yK����B2��o�(���+�>��0��CW�v	e��|F(�x��������g?����i�dh.��>ʱ�}�1�{
�ݓ�9�L�l�����/��}4Y��1Ԭٖ<�>�铦�eF*����z�b8�"�]����=	$�-y�Q%�?�����IeA<�>�5�!�a���J��4�#ѥo�$O>�󤞿�5�N��F����K�K@�u+e{�V'��S�#u�[ X_��|�M3"gkVՇ�4��P�����7�?�]�`/��Y:�o�&����^*���Òs~V��(O=-Y�h��l�����f�&]���TB��r	s��X�Ѐ��.]の�Oh�3�BP<8zi	�\q�|X?j4�����s�`�	O����c�h��,;Lz S��*mQ$f�0m�B�+�Xi�T{�#�zFQ^�g�iE2�\��e��J`P�;�c������`+}=���rv5'gTj�<M�=G��550�Ͼ�u[�3w_}�txC4��ח	5+#7W  V;��x�.m�2t�Z����Iͩ�e�M?I���"W�q�Ms`Y�JB��NRJ��=�#-c��9�>'NѪP_y2��dӴ�ծ߹ ��C[R�2�G}Ug�+3���F�N� � P�C8O�=j6|c�뵺��p���l��{E%���Qm��I����b��:w�A!6���8�1�w��s��+S��n�Py���������9�c�	õ]H�z.&���ЄD�Lh��v�D�f��V� �󶱓CMO{��8�RuŮ �����T�ԫ�8bYt�
�ڝ�H3��'����o�� Nb��bT�qz>��t��O����B�=R�Ɖ�:�A�rfb9���8-e)W�|(��7x1y�M���,�"ܕB	�,o*~W(��O� �'u���@l���'v�	5T�y�#��Ew�VdXO�p�¯�#հ}�-K,��ɳ)�]}-.,���j��bW�W_f���*�m�����h�2d-٥S�-�H�qb,(DM��b�ʇ#���<�Ru���X�2c �vm9��#�������u�Ol�  ��k��G>^;+έ������������c6,�;A�,��[���'E�5�p��>._�9kaI]�Zb1K��c$��&'�hg6�2Us[�n���hl6�vI������a��qt~��P���Kk�q�.V�����ơ�۬@$�	�3ZY�}�����O����c��#ˀi9�jv�إif��lB��t�4ę���y�2D�+��ck���Efh��f��r:�B}�`���o.����g�0�Rib��(�?�7�h������S��NA(1���ih�u%X�lC�"H�--�R�؈��#�C�4v��b�@�b��)����S�"C��ѯ��4=����WUt���}P
RP8�����B��e�=��I���f��x��>`Vb�r�A�!?}�RC���?�d)��,HȦ7��j(dY�+�bd���DZ��CH)���l�'g�>H�9
�z�Nv|� :F�v��i����ӭ�c\*#Ȗ�ɶ`�*�P��Փ����[�o��Q��cj���=�ã�_���^����5�d�f-vڥ���(�"����
Q��zgD�e�R��Q~|(����xa;^ޏ�*؉�N���/v̦+�Y�
IA(5f����ǯ���J��M��G�\�><Q2\�(W���RyBTXƍC�jx��^�����Ee��RG_q�ֺa��w1�rG��$ԌSd[���p�`rr=�͆����ri�k�}�n�t��峭���+E���4�&�7�jtn���=��u�X�_�U<ӓ3�O�7M+w���3�VVf^&���B*�(���e/�)�I|7̻DZ�Y�<��f 6{����j����"=�V)$7�Pk���$X��Q��W`��S�CyD+K�<��d�M�}�q��G��[������z _H�d�?�6V1%E�����h���^��X̢=d��q5j�*��e8�ww}.b��8'Ը4D��@f��*9�{�q���NJ��e�n��?g����X�`Mww���0�B�4��#�M3���Ģp@�~�,y�'Hxّ�n��{/��ѭ���,�
&��)�^̅MO���nq��
���#]9�xk�Uҙ�����^2vahg|.�4��z�vN'�W!��F�t�	�Q�$��-9�?g�V����K���ʑ�DFf��Z�y��\���L8P��R�i]��o�?�
rݬ��A��
Ff�?��P��O��g9�O�@��U��P�	����C�h����/��ջ�[��jK���h��A�u0���t��l|��,g��9�A�caK1t6�h��7<*��+i���:��>ivh�Ƙ�����H1��β��ۗ�#+�9.�:�}�#��O�+M��oIT�+ىĞ0$�zm�
��S X�rA00f�|���Rn�iR8;s<|��3�KE��>a���^I�7o^L�j_��F�G	3I#b�&�.S>?G�azԄa
��)ukF��ǹ'M����ƫ� �i(�D��(�I�'Uv��:K>Φn�5tx��U��G����Oܙ�򔗧��Dd�6�U��g,.F6]�h�	\2�xJT9Ny%�X��xt?��w�m����I"Gڡ��Vg��-y��e��Z�1��W�˦����8��������e�C���J��Q�s&~#����G$�����%��c-}mrn��A�WXy��<��Ʒ�QY��00V������5�m�Z9������`�Q��H���P��08�k�x��bf>&EG�/�Y�'��S�8�(�C�e�w���5h.���bM�U"���X���R��}8&H����u�9@-D�K�#��	"��O�tR��<�	�?$}Nơ���+[+^s��<\w6�]�6+�f2|ɧe���S+�b��X:2x�����n��>��툅@ 8A�������o�zo`0r` ��E�G)g�3~&�͕�\�RaD��3��VN���Pyp��G��<�"f�;�n32��V�.�A����^�:ܷ��6XrNy�W�j� ���)6$��u��#�p@�8���T�1%���#!�o���������O�N��R�~��K����.�m�R��M�O�Δ:O�����Ts��T����x�o�p��h����i8`*���ӥ3:K��d�PSK����PjY��J�k�M(�܀�Eo�ML��/���R+�Z+@�YRd�;��/)װ��ؐ�����p���ѵ�ױ����ia�̄����� g2���a�P�����/�NX�
t4 ����ʱ�o�d�"�"
���9�|84b�Ag�e��w��l'�1�|~�g�~�mRuӈm��lio;_��V�g��������1ҁw����G�d�y���-�Q`%��N^��%�)8^v��6��/*`�[.���3��t��}����0*�ע|d�А<�.�6�J�=���`�b�B�]Y����?ރiն�,a ���iUB������}���a�1�)�qq�wh�Ӑ���-��(���Nu�L�D��T�]�SE���+��<9�a��Y�r���d�I���M�3H%�J)��g*��1�8�������� ٌF}?��&��t%�Oc��2���J�z9��X��
�r�;�E�?w �����鵅��2;�A�Ѧk���Kr�(������ ������&?PH��{jB�i�խ��y�p�L2R�����╊�M��8����k���E@��+�ɳ����N`Fz^o�9T�mJ���1X�1n%D+�diS�kE�E���oN����8��ŏ�,B.����UGst��\]�����c��	+z#uA��F�O��;<�X�f���y�ϼ��V#�(47��b�2w6' I���~;���ߤMhB�']q_��1~�Q�QT2DkN�P{_w8L��d�t�ފ���68p%���e�B��p��QR�i��{��p��3�d��'��0�`�� �=эNT����I2�OB�j�
�������w��c��6?� S=/��kY�$�&[-I��J�AO�v�Ts��I�S���(a��W��'�|!�D�/���]��F��R�Å��xG�=����(�	W8+Mbdy-���%j� u���� �#�o;lN$�b�.F����ų�ϛ�Qyv#��¬���(�ʏ��V3�ű(D�5�e'��nZ�.�ļ7ʖCH����@8:4uM� sK!��ƥ�0WC�#�E�g�.���6�6��su`��g���&���r_�^�0��y~\!$v��;6�����z[R���c-�ҹ���'�"�Jn�v�d��i���E ř���!���Rf}sW�/�>�w�C{�_4a��f-���I�D+>Ȑ��xo~6���MBA�-"�t���s>̙��`�`���\�:�LD�(#Ӈ*L`��nk����2���]��8ծ�yHt�dku��?g����J�(%a�� oC���U���Z$���J�>�p�d	�wn��[����'��s_�&B5Q�1�������ˣ��9À�X�D����[�x�h�
����<�w_p��tk��tŀ[�ݳxj>dC����W��	W-j�5���r���ǁ�B�_x�0vcd<�<��ō�l�ɝb+���#�˰�>"�� ͛��74e�X��[�lT�p�g��2��bq"c%��ٹ�n�A����'E�'kQ�0Y��qj/+EFH�K�J��$���p3zH�%q�m!�X��6��>܇��w`�h�I%�%�p�u+Pd*{�^[�/���0[�zB;�qT���O��^$�ƚ�:ݲ�/�(T*!,��9�+Kd�?������ԐL��8T!�$]*��Izμ�^r�؊Nc�c�AF��Y�[g��gꛓ�(eҌ�e6�w���0��Ƀ�F��<k��E4�\/��r�R��z��;�^�.l�v�:��A��?B�8�^������WM�O�ǠQ>�=��֛M��\(K5T�f�ur6ǀ��2�#ȿ�$C@�I��z��|&���I��@܎����RcQ5���=r��R�b���K�i5��E����r��#�{�'`�x�+uأ&�}"��q��
?@}�H/Y1�b�����A�����jO
ֻ��
�q&k+�x�ӓا��_�]�s�*eҬţ��o@Zu�n���An)xN4���ab��8L�\��v�~`��'��;�.3>�SS��L:2��'�g'j񩥫��@F����B"�.�q�]"��+�8���:�Z�T�g�����V�Q��[��`a����uj��s�qb�ob�������*�?��-�w��n�d��.���T�l0�����������~�bY�l�ҙ;�G����$�;	3=Cx�U�gLh�c/�Wt�f��&�a���	F�>I��t�&����P$oO�L��������鰼�྅����
�G��?Dd���f�����kY�X�B� sFK���h�K%x�)*�K�a<H�Ǐ��=��AĞ W����[&��yƮV2�oz|b	�W���z^#I9�NY+y�@��}�l��҈��t�t|��X�K��z��ٟ����ƴ�5���ϴ/�CQU`��$f-��Wq�Ud�j��<""�B:�e����c͠2��el��q�܄�-�GsA���E?ۛ��v6��T Gh�����+\�Lߍ���5�U�
k�H4��9O�K����A({�>�x+����A���4���
Ⱦ��_'n�8�xG�;��`�c�,�(L�ФjՆ��Ƒ���8Hmg~�4�t�pɷ5�V��Oڟ�%b���M�C�Q��0k0�G�gQR��������A�ýS����^Xm�C��&M�E�ǅ��$}�C�b�#(�A��q\T8�>��)��^}#�]l��bՎ��q�.e�@|�_x�,���wH�;��I�C8�¥s�6�$���I8r����0�<��xPǚ�CJ�۸��2�+a'��[�vQ�9�G��Z�{�.����j�8�h[�V��C�|P���%kQҡ���
�!SnnG�[�J�l����e�ݱ����^ =m��!s'y��7��rq�f�W��rs۟dS��i�rk�]B����T!��E�I?�����HrH#�Ӷ@4�)ɇ���qD�QT�<d�I���p������$�G�r�*��z<����U�V��VN�����{}	h�sg� Y��&=���ae����zw��?3<���>��9�����������3�j%]�m�2��ھuN%����@r�]f��a����Ôp~'<{�%ˈr����t7=�$�檥#�b��-�9��`Z7�j��I3�|��<p�';R�CKgI^J�9{�X�7w�Tq��my�J')��w�N�-)�:�JL��#Z�|C�p�d��V�BI�i9:NY��.g$B���3��F���@�f��(X\Q|��8�@�%v\Iꅳ�Tdu�~r�2*�X��u�����&E�}6N���h�ZQ�?7��=��;���`��P1��~����<�s���棅7�f�O��]���!;�qV��I�PG;eʬO�Z�Z8U�����&���>J3��v�E����i�~��؃J����0Lq�E�Y�ъ���;���yA�FZ�vz*7s�o�1X���2��^�C���iσʔ�;�? >c����Q}阰�P��H��+��)��U����k�7#��#���(Z��	s�0�AD�2��R��F������ȯ���r�����W ������c�lu .��O&U+�V̰�n��ʧZ�� ���s�����*�4~�������cef���y>ʽ])���eb�K���Ɠ��ap~a�Ԛ����qv0� v�]�T��j׶�ݮ��85H����?��g�>�?�F�j�P��p�~�?9��+X��Z��@s�	(P���N= ��0�m'k�+���|۽�t4��H����'+�E�bN���!�zLj8�O���1+�8�5ƓYN�}��@�e�=������Vz���.~f�e�)�R�*�� �7�����Z�SIW���&/��w�[
]|{�6v����Xgq��_��n>QQ�Ě�������7�����o�G���2On?�H��7��.��KAծ�2+w�����f��ޑٟ-:FB�
�ڼ-�\_>��}I5�|aW �������1`�����Q8y��F`�le�o��!��|�����<m�UG���D+��~��/��@�.���~w�Wn���� �b
/P���*�3s�Ȑ���kү��vHA�����N^F�D�ՒzRfE�[SlO�1�6�E��l�Z�`��S���I4Ά���H�U���@�R��+�S��c4dpY@�t�X-E>��������|h�/q�p�a2���>�AV���/�;�����v��"�_hnmܵ��懢pdt��`K�a�c�nf],<gc�jÍ��]NnF� [���#�s㘒Z; bcC��A�a����Ee.��X��s�DP�:�:w&?�!�b�r�;��i*u Жc���d�
އe��o���kVL�?E�����i�=�/�W�|����)Tg��W)&�X0��"S��[����~�h���Te"�AH �4ȿ�k}Gh��s����(h���A����+�Ȭx�^lρ�[�ϡ��a��� �?�� �a�5)��mƼ�V̡ �˲�p��h�W�p���P'��j+��W4k�&����XgG���U�z{���=,��]\�?˽^�3�u�3J�+��[�{��T�5������m�Ձ��P1fR`-)!�
ѥ��Dˬ�g��f�������
���1}��Kh�R��` O��a"|A�ې���9�
X4��鯑���%iZ�"F(��ȳ��%�f�33Ncql{���M�����CeQ)�OfJ�J�By)1��,��xL���%uyH�\���r*���9\ҙ�ڋ��he0�
Akes�uf<pe&��(F��oQ��B��s�-j���+���g5-��ʖ��윥�Z6�0�$!�{�ȴ�i$9]��y���=Y�[C�Km����
�}���e7��#�%+J_hH�}t��]E=O�Rzb��o׎9O�G~���#xVW@� AQ��̔D�~��(Z��ئ�=ֹ�c�w鈏�m�s��o�u_5��Wա6��Ig2y�3��0���7�y]/�$Yҋ�H[�B����A�����(���J��N��X�<s����gŌVuWl��ȑ�|\-��sI�!U|b;��\�>x:X�E$���f`s����"��	���|�#4^��6�Vs�W�~����HЋ�8�E-kG.��b"u��5�T�����E։�d��~�.�?F�Tl�;ܥr��=���V�_Sma��YٴcJm��Z�3Y'�t������"�a�Oi�7,���|�RQAR�e���3���8��d��D�yȠop3Z �H�֮X'�BgBy8�.c�E0��K�9ƪ�EE�?��5��WyJ ��z�zj�z˭�>�.�*	D��;�Ξ2߲� AQ�[��b���@�Q��=�$���alQ�,`S*fW3�]ă�A��Xo=�R�����A��!=��$; ~�N�I�1���{t�?�T6��̈́J6�;��<S��н�L7U�-Ϭ�8xK�K;9��|M�_d�;�ֳ{]�̻W�X5+1����}�&$��]�5�*w�����U\��.���U���'d��nӒ�Ґ��b������ߎ��Q��[�F�^ew��;x<���-�])F�M� �U2�A%�j���R; ]\]�=�f�l@�v>����F~�%��+���L��t����ßݠ�zT��djM�3]��)��Z�.�%��DK=sOBٟB[�Pm_�0+���Fzw�ϝ�`��S9K;��2����\�nZO��I¤bP:�d �E��9�cl7�����H���:���4y��(����ñ�o�7���Kx��~]�h��Z�y�� �!<
`�?�@��e��K`��d���@F��>3J�Gp玃���G-.�c��G�(e!�$����k���&_;g�=W�Jϒ���QK  Qё��^�
��5���arIu��!�j���PW�?�⹳�nޗ�:��l'�-$-�+A�*ڱB�j-H�>e�@ه�&A�	��]��2V�$U��F�E���d���X�rw�sa�?�K��R��L'���3���Q�Ԙ�-�P����A�`��~1e�%�~ď��xp|�Q��j���Q��	�ބ����5h�p�@��JB�k����qTc�0��.���`�� ���#Zn�U���-��?��"�*�ӝM��(�@�{�'V����IM�iI��l؈nw�ե�U��z��@���I�^��P���!�P)�Q�(���EF�@� 1�����Q(\<������í}QKv�2�v��&�Y� ���2�w��{���a�	���f��l)��� �񃽌�6�6$��˝NĽ=�i�$	���a�E�g��W�:<�r��Kd5`����X��w-X��9�]��υ�Ή}u���j�2�(���cT���h���rC�c4p����Iի�抁k��53��H���_���șQiꌒ�m}�%���m>��E�n����2�1������0�����5����sQz�}�j���@�:De���w^�!�H����)M7+!p�?�u��B���*��g�&��㇁�S�6}�2�7�-�	K��O@!(�N��BO6�"?s]Hr���&�~I$Ѝ�+�Y,��ȍ�7r +��:��y���-fw�莭�^��m�&y;�P��rO"[H�� �t��{��u�w�a��$7��j����|r��u.��+82�NA�īOW��Xœ���5�{CyKr'�{�傅#�/�]�p]�7i.n[�DǾ��]��]8�>[�pSw�htk��z��~w�%3��z���!o����i�Q���I,7���!����b1.Q�����x�.$�j���Q�\��*�KXb�����6��:z��HZ�	�lFdl0U�'�$R�D=U� 4>��А'��Ci�Z�\&�	�lE��Ϧ�mm�+�؋�^≼�f��+[��29�[o�(��]�9dZzK���b1a�FCf +P���I�hκ3��&��B�A�%.�,3i'�R���
����8���D���Yٶ�*��, ��I���_�f���yI���x��P}��'��Ğ��V.��⶜�?��ܫ������� ���7��h���vn����>����Y���{��Kx(ߓ� K�tÜBi)^�}�Jm+K������{͋�� �0�Y� \d!�[Q���<�c������`��f�3�]�5>7ОvLcȐم덶E4��J�������U��~9~Iu��dVB�_���.�/W���?���U����=���ĵgfT�1�?�;|��_��A��y��)���snK*0�z�՘��z��)~�Oc�'��IC�jD��!�))�^�u����g���b����v]� `$ �q�w���'	x���)���J���L��)�Tu~3�n����Q�,!���s퀞�5���Rn�]s�9fi���FV�3�d�k5�Ӣ%�����کbh��z̹N��qk����Ds�(���@��_���0e�Y�CN��
���}y4�)���{9�s���\�m<���k���@x����$�W�P�Z���b�%D~���,�X�oƧ�u߇������Sz�w޼.��Ի��W�]ق��x���u�?��CբV��뗚|�<樓O���B���c�`l:F��/O�:�H=�� @63	��ע�9����!m4�wv�	��s1�"�ŋ�t���\_��Vt"���.������#�i���kx��K�͏�c���7�Q��zj�|*�pPJ��!�-���{� ��� +L;�o�����G���hp�[�}�k�[����!��Lч�.��I%�ٲ������	�ӄ����i^�/d}*ՙ'V@�[�j���^�$��Y�d�ɫt��2/1{����8IG�pl�����F�)a��K�6�ǦB
P���z��@;�8��R� y��ӪU��R����?L�e�.˗q��~H�P.�"��u�ꡱ v$܉�7# Gm')�$ni�R�@	.몲͎�������d��g�B���Dp�"�����[m�
ʹg���H��U6�]�o�<�Ҙȟ�aMI䲪JI�������L*�Q
��)ڮ��*�G?a<f�5j�@w���!���[=K-li�FՊ���Ь�Age͡p�\���ZhE,㜟����ay�-у�TW���
䤥�ǓX���W�ԣ(���^��Rgћ�a�	�*�2������	�~�n��)�zݚ��OӀr1K`8+C�ެa�Ǜ#��ǽW�r�N�ǩ�Z�|�#$���$�C<�(v";?��\	�BEOҞU��(Ō�&����L��H,Z�{s�BiU��ar�:�M�%撂�o^	��p4^+���0N]�W^I&uB"��Ђ� o�_mj�`�;u�]{���[�����\U��~���]Q��P��"�t^��.0~�'��sQ^��u�!������C~��Տ�Eu-V�7��7p�+B��@.�Q�"�:�RU���+<DƳ� G���&��xU�kgP�$͏ǚ9F'����U�R�9�
��ՔhH��M�ސ0�q+* ����G
��~9f�u3l�a�a�w�r��7j�	�1F�/U��h����W�1�%lͿݷ�~0�'	~=Α��4�k ҄���4��d�Ƈ��#Ծ��+�{�Շ7<�7q�Q�:�<J�h��Lɐg�E�9��%2j���@���*A��������{�5���(���Z��p���=��6a
���<��[a��J��i�Vp��׈��p�^/ t����ye�]�+�yd� ��qAW޾��B�[�[k�XKK�w){���v�t������~��,��'&��ᬛ����[�g">)M�1r�O���cQ���E>3�D���UĂ��U������<E���:�K� �	���M��R �n�=;��I�[7Àc��LU�j����Rfߵ��)i���\��s`�Jn�IHqG�]�A~R�k�\],�6�p�  ��TF�,]���ժI6����U� ��Q/s,`����J9�_���\����L��nQ4E����T�⃬}����N3��|Vl��:��Heg���WP8����g���ېe�=:ɲr������lc*�A�%���R�P-|vv��������XV_��r�ڛwE6f�e���BM��kL��b���s/�����~"Ek� �R3[����It�6�_�߂Nhw�xZX�{�^'(Sa�U�'�s�����F	F�]�M��ǰ��3��,�5��;�K�s�H��b��r��-����j8�FउK�hp�Z9��F<� �n��
#�N�
�քJ
&�ﵽz��y<J�mf�"9�+d6�>4���w.�7-��穭FT�u�Y	�}�\���}��"#������BP	�x5,A��p�L㓕��ޭc��\Q�dA&WsDk��	Q:�.��+���<�������vM/���dq�q̼j�?�k����q�g/�$�Q��y�uΖ}A��6u!�U���G�5��b)K�=�l/n�̒�[��i/���&�p2B�j� wy���NE��	���8�Yf��Q'B٪-��B:ನ�*�`����]��8��m������v�|�����^i�X悫�$g�z��^hX�㰬>fa�!�YpO ���l�?F�?�*���UI8�r���o]Y#�������3<�N'"u kQ�[+-�vX'xj�}B��I�(�l�%
GtmH�l�l6&�w�R[dq��  ?��a%�n%i��>����̇/�
'-��L-]�%n�]��E���Er��)*52�Q�N�+];87�
��/"��Ѝ*��I7���U 0�J4���^{>Ea���O��4�N�V�����^��*�������Y�Wi�Wx�Lޞ���M||B}}VZ��fB��2,>LN��{(L'Pg��w�)X�x���	��jR5	əg
p���į��UAO����*e|�߯�paq1ټ��uL�%�����@T
KP�'��п`~�����5���q|���>zp�.��  �� Jj4�x���ز�5�Qe��a��xG�$C�u[u_����7}��[I9Ե�7J�T=��Ϯ���ֻ;��u�y"�]�P_��7H�����BX/�Cs�W��q�)��Zر}�/>���"�KA5?O���iv�� h�[n�#�V5����˵���m �N��LR�W�W�Orkv�H�������8�^�)Ò~�syR_�����켏L�w�Cs���%���k]�s��az1��=d�������k94R��a[��5ٮ�ó�1L);9A��Z)u�7P7����ϋ�,��(�a"�R<v�O?�h��� ��5k� ��5��'�GG��T�=q��U��Z_u��jSym����y�>�h����d��7�M���%T�=9��s�E\�M����X���r���<�&�'�֔�7�6,����p�rj�[�>qЙ��}^̤-�����'>?,���L7~$y�TR@�g"��ꂢ������^[U��G?|F�6Og?Ș�Tj>/g�Ӱ����?�m�n���Dؾҭ�<
ȠD���p��J���R�9��I/h{�nI�K�.9��h�3iW��n��Ϥ$JS���_ÅZf\�$!T�e_M�^�
�[��|B/:�4�������$����Ӈ���I�Á����d�$=��������A��`�1Jdl��5T��4�q��&b	�ԗ��2!M[�]ϐ�  ;�N���r,���� )�a�B"�g�+���E00rR(t��j�q)W�W�F�VZFk�4��0f�h����MϚĕ� �^Yc�7淶e�Ky�!���1�0���^�Q��M�u0�!�Ы~A�G�:*����^:|���[�h�䈔wV��[^%C-��w¿�±:F�7|����}DE�ЯNo��ը;�*�")b��	���}�����a���ϩ;���_Ez�Ԏ>g��$}}��A=�=a�W�p��@4��0�IkŏĤg����G�) �4>̼��
��r�X�+��]��丌���~Bf]�ۊS]���i� �Q�z=W��(
d�S��>J�.�&�td��stո���N2��`uO^"�
MMPpT�rC �9�6��	��~�pD�eu�>��-|��AyW���)��{=W��r�G�U�(_*�ԠDn�B,�&M��[���r�Mg����ʌ�.=0u���O���\�pA��
���&���a�p�Iؙ���5��+��1G`
��*�0|�?
/S�z˾���Qd�YD�CV�d|~��c�M�"�X���s,"_ p���A���G�\z�a ѝ���"I��im2�
c�<�RX�ԝ#�6d�*4Dlv�`.��2g�a��������+�y�}f%�˝lPu�����e����r�QAt���.BC�P���e))r��"�w�HM�����P`���pi	���LP�Yx��-���P�N��F��F��sk|F�9_K�2Ղ{D���S\����[{��ߑd�k�@iJhN���q�;�T��y��7��K��q�]rŽEB�'�ϐ�'��D�
ޗ8�\!����_FY֪�:��!�h�Vh-h�k��]v�o;v[��f�Q<a�`�h�U@g��~��i}�Dv���2�#c�����'��Bc�j,����%�1}��R�:n������h����w/��tu��՚���j�GJǞטn��=s�)��}{t�<�>sh�iT뉭�2�T�����|���a�t����։����w��#�o8BWt�>��~�K�;0Q��b6['(G�BB��1� Ä�^u [�W��IB�K(��G����J����ھ�S���Yh�N^��ܸ��ݠ�AR�j�H\�7͑��9����c���l(���� M�:��޸�f��z�e�,Ig1�3���s�_�3!+�O�K��n=č�c�����ۯ�n��L�ޖ�G3���76P	$3�.��&�`��G:��f�+�k�8�]P�{o��-'��zk�a�K���͠����
���*���~g �=T��nV!�	/��i��[*>�Ze��S�|�y܎�+�1�]f�=���^~ٖ��5=V'I�W�{��wk�����,"~�u^Wy��f��[#�,��/l����$3��#pD���
��j6M�b޲�k��,���N�`��S��L0��i"��J�\�� �:>Iu����i��K�����zs�������a�%�/�i�P�k�M�1��(��j~�!�u�G�Ĺ���Gv�gr�l_� �4�C�t�cu.�4��D焵�-3\������%�\��z*�y������o�E���8(�n�>n�c��.^�d�~��r��\+�KE���u��=�8�9̉�09�5� ��6�ND�;�cһ^Ž|��8���`��y��͑<����!S�!�Jt����X�����0�JG�K¦�@����#1�Q'u���|���2���*�������o�)Fi[�
�R�:��+{���]��h�^%ƈ4�a� �;",��o%4��k
,�$O��6�ۀ/ॽ���xȽ���I.��Hv�߾�|�dj���t�����i�u^AZ�`x�F�~��]�Q�+�	�WFՑ��n��^z��w�� 8x�,ߞ˩��ih�W�eKMq������Wǽ�ҽU��N*��j8��&6Y�i>jv�}���F�c�����k���[�k�!��(�3b�i@F�]�,h_�
Ί:;�b(f1�{�)9�.
�Mq��X+�����y�1�i<ԟ��	Sd���AA�v#�1F��Z5s� Ӿ
!�d����$<���8�Y@��H�'���{�?�ѡ|pv����K\E�4u�A/y�5tw�L�����CB_?�����m�,����qo�<�V�2���+0�#D�8!y���>x��}gy��y�F�ꚩ���~�^l!���0g�,�@�fД�~þD��3��f�a�	#�(;�[�������m�2D���c��ϥ�Y�a[������S���6� �K��2��kW�3u��U��-�n�י�9��V��c��%�q��ѵo���i���Xl�ZHӓ�]�A�Db2U�\�.����ŖTֳ�DĂi?�_ uL\�+��6w=����1���j��E��X7qn�h&�n�%�$���uܝ����!	�!�TV�}Z�'���:-���y�� ���V��"-��%|h!���5O�H�\U���ߣ��fD�`���	�s���w����7�â��d�� �%�pf��{v���tb���j��X+
 +R	c��%#w��aNOTs�����nf�c���Od�F8�G8h�EW�K���;�S�%�!���m�`e�nA@r�r�+��̈́�a�7������~Y���B��=��K��UAJ�.�q!�P�ϡh=���Ķ��cD�G��&K���ĉ��!��:!t���h}qϫ"��rcb:_.��1Y=���67���L_	*ٟ�И_p
W��t������������Hú,C��Q[�)C�M��T���i��/��wg�m�`�Q���S�}i�:C�\�l/ka��{/~t��b?#u�0U�WCZӌӻ���:�
�Ojb׌��%�] hTN�%�x���mG/�5�!f�TC�ذ|�6�.[�I���`A��C&�����Hv�~��ʒJK{61}6��!+���+͈v�oO��s�;��o��jN1��Zr`�lO�А�ۼT]���פ>���ِT�3A�~U��������`b(��($�)��ڽz�F?̭���4'��٘�����1���0�`t�5���0�vZ��OM͏��G\�M��w�jie��1�|Yv!z�A;Rp_{��(�L'(k����uldKOdː�U[ц���K6.D;�f|
jsxE>wVJ���ܣ��!�-F�h^4Fs��m@���{�C[���e1	P{� 1Ɣn�T��ts���{.��0I�6k�2��rYlr	6}ΛFx*aT]�0��uҁv<x���"����	�����ob��T��G,X�����Y�΄��ܛ�(�~AL���#Ǭ�[�`�����܏YR�����{���g{� ��;��-��`������^7H���	�g�
)��>��XZ	��:�.�[:5�[�������ϼo�ki�Ě���Ow/`2�1�^-լ��USV�:��G�	��{G���Tk2���<�}�����y��]�࿸��6���#?؊+==>w����0l��y0�0��R��� S�oq!TM���*©�
�@w��r?B�^1���2�u�6����.Q/g��OH3�iEB�̒x��G**��do�Πr=gEJnз'��³�	#�(��xs��P��J��Pb�w&r���>� �5��\!���b,���K����ي%D��X>���ϧ+��7��D����־�{���X�T��0 3�R
�/xU�*�W����+���l�ۦ�$9��&J}J�*'�bj�eȟp�'5����箧r�'�O��ŵ.�
߭��Y�0����1�V��M��m��Ƒh����W0bl��ZO�fq .�$�8GZ��Y��!Q:s��Rh�
�@�0{&�J�\T<�c�ެ�)=���K!w�����#痤����ǳ]��j������˂�\g�4���@�EK�E�W���(�}�R����#�C=4̤¯�P�8z�AXu�<�A�$�g=�*0Ǣ�xTvR�.x?�[����hB�J_�{_nn�N��E�%nK[�n��?�X�f�qh�Ҩ�-^��U��}�9�����}6K�T$��w't�-�����z7��������m��e�jS��*�����sU?��]�D�a�	�|/7r$P O�w��>8j����m�f�N{!��	�T�ק�����=���)��f�:t�k趒lƭz��z$?�R�+QN���%Vv�z1����lXB��?�z|�D���	Fd:/eB[����������R��y�m�
q�;3��R�Í��A� �Q���oوT�-�"r�TuK��|ynZ�w-��*�A�-.��������7>I���S��q�oxR����}E�?�ի�V_��*n�C�a�¼rC����;g�閣���	���8Ӑ���`�R�/x{K�gk��^������c����ɵ9H���S�.�Q�
q���QQg%�fs� ��� dX�%�L��~�7)�;g�P�1�@4�Q�C����1��ϋq�<!`�b3b'�8�>NP��(�D�Z�
�Fj)��P�e�҂����jd��<o��n�q�'BL�7�=�gh��=����Td�)O}:8��1u^�ieP?�l6?�����/DQk�ܠ_]�)�3a�C,2zgT�YK�n�C:I�g�Q}��H��-��%i��c}�蟦UV W�s���Z4U
O��1�L	�: �t1����&h����X�|1���pt�]p}_��:Xh�w^.H���Ә�w�)^�d鈏5*yP�0�ip!X��~c�k	AD�� � ���nS�͠��y��1_p��j��iM.	>|J.>�߲e.�utf�F�瘐BIb�{�P�
� Jh����e�0���ן�f`&k Ɯ7�^e���1<�I	.l�h6��t�����J֜��Ш�8H��ٲ�� ѶU�C{���S϶�1���\���K��/���8�Sm5ɖ��|���8`����9��a����B��K#����^w6�Y]-h��~x�[�B��(RX�d�A�C&+�9'D�Pu��^rk���2 ����4{�%7�fz%]���Zz/����%�o�
�����7Dqv��6!9�-�������@���YT���8t#d�Q��k�F����H�(���5P�y5�*�mbڥ�Z�KP�*r�lU��[�g���z[�@n�}ǐ�9 ���U)u#˓���y�CEdV��`�W�~p����/�
�D#�D�`��t��9�^t�vP�7E)5.4�����+�� 9���{C>��g���]�t�p!�ѐu�\֟����2��D�z��Rv�6��/�Lc���h�ɿR�`F�Bhk�jԨa�-�~��{տ]/)�,�5�9�5;2,�-�'�£��ߺ�xH��<����%���GwB?_ -Z�r�h`S�up�3�>����ZPc((�XD����� ���GafGq������-�l��XVa"��)>�{���a����4-i��2��.<�]�ph���7��~�� l]�8�n���`!̦v9S��x+X��\�׿.N
�p.�TC�Io~c1R���l�Ƌ���a�)8*<8x�'�Tj�Wy�%���!!�{K:DrbT'Q>w٥&%[ �x���\�.[��9%߃��;CE$��#
l��N��܊�$�h���
O�B�{ iۉ���+q(���͡����H�:��?�K}]�Pl;���i�p�� J���ܞ����������S�����Y�v�������YZ�#e�\eV���*�X��G�
��Ȋ�,F1�憪�:���}�p������`�����Ec�E�6�Z�>F�ڴ>v!�9�$�j���>��n`q����R�+�2����QS�ƝX�r�DA�/g�3�Z+$��u^0<,
T�R���B�L����� �Gx�KHU�}�㮻@]$8i$��@X�iF o�������UF
�:0��a�Xi��?Z�3��_ j1�ٰ[�xvE�T�:���x+5M��y�+#w�{�;$xe�}����d�QN�=<Dj�;�#��@�b��vK����������$�si���j�Ң
f��5�z�f�W�$�۰l<9�y.�:|��`i_�����BP� �ͷE_�[*�lm�w�1��FL߾�SȬ�&��Z_I��XO�[ޣ�Z�g�������,3�������Ud��j�e�!�~v����xg��.��iT@�����:�i�}W�3Q���`27��yٳ.��� K_���8!�K����`)i&6rO��cn�ʘ��̘��|	=�iX��X�@���r���q��<g%�]ԭ�{�(S�P4�bC�h��{^
��M��WD�%���s*W=/i��j�̝L��>sJ���%�f%K�H!ZPl�l����ѵ�?&���h��0�����=P�\$���2�n	�t�4w��򂪯����"�s�wvprK�3E}H���l�dV;�].P����F�>�أfPq2!�̹��41B\}sq�7<>�u�怲��:��p+rG�e��6��5<��F6�Fǉ��+d��lc��MkCt�Jr����}+�R(Oe�k�Z��_���;	-{�c'������k	9�3gvO���Y+-�w��yn�r�F�K���m�#<h�U'�fc�.�M&bb��(��"�B��p�����GS햺�`�;i�gaҾ��h�[��m����J�dM��T,y��YBm}1�ޖ2o-G��#ӽ��K����
vA���泺��M�8��T�{������2�')*�<o��]_:�p��5��ۣ���C'}��\��"��&�d�x؂M�[X*#NK%{�b���;��� \�������Zy��6�?)�z��#�w̸ga�q� G5�8�;'����z8�����Y���Q��н��� �3q��e`,�q맿'�Ծ�w��p(sQ���}�C���F���B�G�_��U�?U�60��C��hy-x��㔟����=�Kf%{I�zETM�b|f��`�OV���H>Al5hc��V�$��d�eX6X$H��i�w���Sjy Z���z���jq#)1lJ�B�7�i� ��[b��ǚ��D�!&=�l�W��=|E*�/ؓV�>��P��燏��4$��M��"}�Β�#��� �ф���A
��O��A��L���N.�t��u�c�Qoa���L�H4SE�NV1�v8nQ�,fR���^+}'�c�T
�'[�����%i��sX�f%�L�k�K�Y���BG�=�3+��~��gE�|(!�!H�+�����q)st��࿕��}1���0�t�Ն���謖��0S�M��������;J�&$A�[+ E�zO��j�1U��a�s��S����-@��Z>���~/j'�B%*�����~�Gm\B0X��.��]��)i�*�T,�p�����V�Q�K�:ۜ>�M�NT4'��ji�gԉ����8�k'"�hnXI�k�e��a�z$0��
$޲���.��Hu�<�]�b{�+Z��*���'�B���P^�=C�����sj�ABA��{,5~t/��|�F��.����x\�c��ygU�׭�/bAz6'@)���-���jf �/!QG��^*3��ˈ%�����]A �AvJV�P�@��cb�%��淀t�2�k����i�b�y�5< mH�vS5���ǑΤa��J���	9�j;�S����{J�Z���}3M�������]����(dg�=T�q��1���	�J@��g�⦷#���%�q�,�P���-7=W��p�UQ��^E�4[��w1 �~�3�E��B[����+3C�������#��B:��L-��-N
�QRAB��h��ZC��=G�qG�����'�Fh�{�m�R�ܖ�GN�?�$x��H�"�tLm؟���><I��ՇSش�[�s���¥Z�J_��-q�bE��i-iUA�|��ȝ)�6����v�1b���(�W�	��ہｻ�'�=�i���O����$ڨ@�Q�椒zs������hTL�2\LcF�4�������'}����j�1S3K�p��sU�����A76�Q��5:g�Vhnֺ3�s4c�R�dS���y�#�nl;Kk�B��Q|��"��T���j$ �M�)YV��L��_�Fɶ~�)��z�-��`b����Ͷb����Y.�l�P��A�F����]���/ƩQ�\��R����0zw΋p:�v+���#�@�xBt�����0=6�dR��oY�n��Ϲ$y?ւJ�ݟo�Ge�eu����x�"���ذ25}9Ch�ӄ�N<b
$VBo�t#nč�H��*�}`���/z#�xZa��_j� R�,�MF^CT���(�/��)3��p��@�♡�u1hg�7��l��C�m�d���䑦����ӆ�d͆L���qJFΖ�ׅ,�ƙ�^�y��1�_�{�NSt�\��?y#��kf9��m��"�j|��+�-�@���^��^P�LK��g+�`R�eM��c�Ñm��ۣR�� 3`��K��Y�u/{�w�N���M�qT*����m���^/�~��>���M�.\�)��Ŝ���5�^��r$O�>oWN�5����R2���1�>I���a����ߔ�ɨH�K��Q���������H6QwB��n��͛�tax�\��	�d�\��$��=��[F&�0!-��R��(E΍��<!y�ͮKW,�Bż��n�̢�'zC݉�&E�S��z
�3��`�٦�:���Yd��<��3@Ì@�x��Ggl��0�J��
��2��ňf��EH}�0YgA`���r���:[n ��X-�V;l��G����0(��,ֱ:ά��<�x��Ю|d��cu�V�"韕tVEl��=-��h���XJӏ�}
�+���B9����#L����$;�Ȝ�C��C�5�q�~� ��-x�RM���=�{����0��� ���6�Lh��W�ϓ��_f��t�� ���������9�[!����O?᯵)aE�������ڵݡ�4�.d�߬B��j��f4��+�ΐ�!df��"�2e�� X�$xސTWaU�Ԉ��m�m��w/M���e�!�z�O��w�Y$(�&Z�v�0�X��<�s���sm,V�y�q�F�/���f��v��ho�]X�꣕��x`·��(�Pa�zX�ï�7F����Ib�Yz,+���+T'�T�x�r�}�/�;W�G��#������Q��]�6����,�ض�����v�+,�tS���$�Յ�P�z� +�)���S�����ƛ��f+�Aag����������yfj�ĵ͕����W�/�I�@�ƟU�ce�UH#Rpl�Bi]�BA��Ⴚ_xv����s@���=��t��2��.�t��t	�kq���7�A�Mgv���U8dq�(9�����H�=�D���,=����ыDO02�,!�ϤX�.?dA ~���i�$A��4՝f�A��v��I��FU2Wj�x��!%�7�6V�9Lz���F�n� �P��4�k�|r#�;g<���@Ma=�4��F4^+��Q��խ����8����}����[�`�D�gX��G��*nkI�S��g�&�+��tDm�Oq���ٴ"LD�K�캮u��.�"����������X�;��]&C���A�L�m	HT���ք�� U�ГR�g�e�F�r^��"s\ֹ]V]���@B9�V�u���F�v��7�C�K]r#ぞN�I>�b�!Ǉ�ܼ�z�B?�|��PKM�Z8� �u�t��!#���7cj�H�Yu}9}��V������Q�
2�Wf�
����J�s�rx���v��Z�ͭ���{a_����k�gRy��x�^��k��ĕŜMaB	���%n��x��g���^o�_;Bm�ix.;!�ν>E��U�>������i�"Պ��@*J�`��\��Du���/�� �Zɯ��Kc�ؾ�f��9<�YS���c�&s�S��`$�fI���k�:Pe�.
M.�@�xZ�x婑�aT����͎6�7%t�s���!k�T�z�v/��m�ɸZ���%��q��N*걤3&;�H��%/�K��&K͟�����{�en�SD�f�����ͪ%O(��91��(�@WA�e#:���N�_0�NhS�sx��5�6l�$��$S���ۦ&I#IhY�%�%~���V��ũј{�:����u����K^K�j  ��w`0�����h'�k��J��3��Rێ>������,����j� ﭑ `���
����7n���&����heg��:u���{m�Z�O����'����7�^��و��M�s�O+���_�/{2/DBt:C�83���LF�hQ��Rè���E@���A��$�h�Q���Dv㨪;%�<�u-OE�lXtr��0p;ܫB����%�x�Ie�N��x�N��ͩ}���k�D�P��.a6mf���+������[2����7��uK��?8 ��@�{O��(a��<-����2Wm|b���Q�	f�}4�f��m� Q� V��
{�b��x-�<��o�k�bM���K"�	��I����|�!N�h�;1[��M6;t?$]���"G�5�]q z�Cp���@��z��;TTD�1C$��z%�`�e?��%* �G�3?(�q(��jݨt�K[�h`�Ђ�'������|[aћX�Z�osj�Wc���<P�v:d�N(M8�>[#��(C���]���lV��ú6a�u�y����ߓLdĄ"Ī����'�ZHj:�ky�����b[n�@����h����ݻx}�R쀲T�������Li��۷1���M�:
P*{�_S�:��w̎�U��gY m�&I�IaDj�N�Ī�j����@!����<|ȣ/��Z)O�N��y��My�E,(+�-���O+�|���/v�(+,lR��k1�[&�{b�N�[{��Y�E:������EjVԵ�+��+ʜ��i>e�f��q��S�FY��0֖B�q�y�Z!�CA��"�, ��ull��'f���|�U�])\)_��_+���S5�·B�a�̢�9d�mS=�}����^C�i�m�	K�s�x����W�3�bm8EX���9'��v���\_eI�����R�}�w�A�{U��Ad�o(wǐ�fu�0�TVL�YK�&(�4�17�U��Hv/NXF�VDQ0i��ؠj���X��]�jk��'��^�'��3v@	��AK�xz@DVKY+37)�g���/��L�W_k�r�H <�S���7�L���L�%ί�l�����^��5�td|���t�j�'�n�����:J��J�����0����!��!Zٞ���ʝ�~��R��'��-��+��F˿�lA�2I�}��Ӌ�P8O�"]N��X6j���	](�@���D��0��5#�4�	�җ~��@�Q���+�m��!t(��G1�9Ţ��s�!����'� ν��@@�݉8�Ţ����s���tL�fR���*x���w?%_�r)w����7,��A&8���q�b_huF��B�7�.�jy.o�n�R�����H����j.�Y��f�y�>D|*��(���� ���L� �V�U1 �d���&�%����b�i������W4����d��N�G��8�����+{_ghhj�t��j>����'�ov7PANt�Ӟ��_ �7wP$Ԅ�a��`cvˮ~���J��8�K��e�<o�vm�Ku�&>̟�+��E.��BF�f�=
�[��Q����B���2QR�7gnl⋣��K�!Ǭ��_�m��zD�<��fp��Ԛ��{*l#��q~�{�S
�"��X�գ��HQG�A��B7Ӳ�ɱ��4���$öR �s�2��[-9:S��M����I'6��r��Z�8�K��P���<�'�u O@���,LT��GQ����Uz#|�8ʙ��6ހ0/��Vh�>0���B\`�i|���fb�0i�֓���x>/m�	�,OS�L%y�y�M8-�r��Q!�� <^A_6eM��:�_�lx T�c4��8���V	�%����ЍIE^�ݖg1����L��|�<�=�h8_��u�)&|�vG>�$�w�z�4��hҟ��~m>�]8'%���.e&�Zy=�ݔ5���0���A�l��a����H���=F �T�&QP� �["Ul c�x@�S
[dI�	�$8!�h�+s�d>���#W-7����6(g�,F� ޮG�]o�yΤ�<�&���l��Q���|D#`WGSI?�r�fr��� ���E$:���.�jwLÅ�&�<�7i�@-�����H8�1�?����d;������Ԑ�3g��t� ��zh�<5��D����%>g" �� �֌w;�i���ji�΍8��Q?m��׉�$_���U`{TO���/�~\A��}�ak��џ�}P�_X�b������VJ�y��Ip��;����3��/�����+Γ��S��{�:Gk��w�X��"��?H�Rpo�;{	ҍcf���:����ym��%�T"+q_���<�\��,�� �g�`�Bşp�>�d#E�4B�stwГ�+��YÎ1y	���Lwy�z+�X�.�Q�B∏2&;���+-�*�u��p�(�IGO��wo����IT�"e/��d��o*3]�1X���'�뒬e~�Ӄ܄�q�/ښ���k\�m}}��P���[����T�өDְ�#�?��],��ǭ���D��4��Tu��a|K��6���Mw��'�U�\u�z�U�ޫ��.�9�С_x�<Δ�3�?��냽V�#?O,����a-y�� h���ߤqZF�PI����^��k�m�P"RP;���ݥ�ܼԮϓ����3R�#�S��i��F���s��o�:u��D�� M�2o���Km��P��!�'マ���;�d(}̡���;���3�2�����w��	,![%r;�f~.-5V{�u_:��%ucX�U`d%iY�"�d�>ÑҧіSf��8�����tف�&c�8�Bgs�j��!�xU�ڨ�aan�k[�̦�O����nڵ~wk��iII�#׃����#B>%i���s3�Ɋ��/���K|qw�0c��Q�b�3"%�c��}�d AH�X�K��>�ݟ�.�0N�7��bFzn�>���4Թ���ߵ�LLb5�N��F��>ӏA�JI�f*bp��~s������c�aonQro8��J�`���	����r��Ѱ����//��2+�q��D~���%�Ĉ����GCD.IL�ᕣu=\�7����Ϝ=u��m�X?��c�0^�@ͨ���rK$w'���M�����6R�`փ�̂� �U�&�I�H}D�)�j��${+�z-
E�9��A�@��G]����S�:�SZ����a�=�����!y��2˳qs3I@���b`Z��#��w�o����fR��CY��: S����Ar���l�jc��x�i`
�6�	"8��qtŃ��k˻�s����އ��Ljy���g|��q�2FQ�J��	qpw/v�Dg���S|�'|
�N��I�:��ݘS.�z�0	fȾn�Aиo�� 
�$���?�m���1��27�����fT+�Ԇ�Aۡ�M�vP\������T� �A(���MR������}����(;��281u��L�!W �>���.��s��6�۳�%�Z�R�=���)�c9F�~���O,~C8��%?�՜��)"D!��iȶM����i�l� 8l��^���*l��H�/�b�CpDː��-6��E��@�����E�& �2�5�t��m�ɣ*鞬�6��(��<^	&\��
���}32Hb3�]1�E����F��A�׾\����N�o$��	`��� �T��B�ly+�q��ZJ!���	��r�Д D"��݊[m9�v� ���QMw���HQ��礫���@���������\��;�ɒk~�{�!��*Xw���c�E/LzN��DlϘ�:�.J��p/7�>��H�����6�q?����`P�$L��bS�o*�eU�����>y�;Fbs)�]����w#���(n�?�(o�/�x/x���R_y|T�Q�#;ឿl��b����8>E�|rd26����K���h�E�.�@���SG
���'M�>y��S�#�vhɝ� �E��<�L�HI�ށ�|�`��ħĀ�L�
dݻ`	������p�x-8r��c�e�����LF��k�؛�f�ie���?P�sӚ�ƿv�7�Qz˶W/�����P�=�=K`��_��]����J+�$����8(��T���%�gp��SÔ��U���=���j �KH�9B��~���獗����)TT�L׮�?��m;���ؔ�`�vĚ�22/�� x�������F��$,�x@��)A13��"Ɇ���J���&y�<�36U��z�q5g�6���3�����鬝��n�_��F+�4�C�b���g-{��	�];����iKI�՟�*�[���x�&��Q�:����f���3C�-o��rI���B�_�5�@L�b�l7C�NN����IMq�������C/:??3z�<�Q���WuP`�
��0�p��9 E�i�YGÒ���LÀ�>�s�F�)V_3�c��?�O�ZI��.�3�c�[�Ԝ��FbN-#�jNX�	H�k黨�G��E=����D8C��J�t��Ϡ���bE��ȕ�k]�n���"����A��D��0� L��a�����nRo�)�$f�`4e��h@6
��k$Ո}y�"�� r�Ü}�P�Ěq�S�M)F�<�]��Cp������<0�vB;��i�UQ�ī�۰Ќ�Tm�� �iP
�M���;9�*�X9��H�$���0 �:T�����o/otBv���M3͹e�<ծh%�ȉ��gHZ1J~p��ڲ!��h���i-��ڙ����z��ƭ۰E͈�׽�+'��}�O��X0�p��ު�M�d��|�{(�� �I���S'
�^{t. ��O�	��Y"����x쯈,;�k�F�*�=���*�k����IE�b�ŝ]�d�.��Ju`�܁j
���Zk��P�yg��Sb�i��C�1J�1�n$�&~��ȥBM�:��)�ǾWd�q��=$�su��{��4��Q�� /0O�-��K��8izI�6�˟P���G���O�Y����K�lɞ�����b:��n�{>��s��N�"O;���
^@�>Ƒ�(ﹱ(�r�$���E���iݱ�+2B\�����Xӫ��+��֞�-L�x�����g_K?L������i|&��D'}��A�-�OF�sz��Z�U�?�Sq݀\x˰���wA�(9� ���D��烡�C�,Q�)�4Y+%�_�7����N$�����H�L���$����b����R��@�e6$�n;�3�]������I��-mr92.�a�(G�����C�o�M|�*3�[���-�Y��G�ˏm�k��/׀���~�ʐ��=�F�-��ɼ�J���i�z;���ӗ��C��D�sc�!I������P��uhj�;�>[j����9o�n:���Y��G�;�&	�l��<Pw�P�=�A?	0ވ����d�w�X9H1��ǖ;4�f��ޭ ���e ��t3z�j�k����ON�??;K�!�e�1�"��ZB�!@@}=Ic��̽J �GU�ĻX�*g���!�Jݠ�g���c�j/��q.{�U^NP@*3�mz�j�"��l����F� }�S��)��^�!4�Q����+ʼ���%��RSW��>�齣@�t7>�ņ3z�O�e�
�# �5ԭq�]ˇ:�7L_��V�7�<|#J[I^J�x�@�:7�"{1�E��U⭏c�O!�����?�w89T�e]���8��ٚ���ų�q���%S�U���ή}$_@��@�=�Zg�y*3����A��>�eHX�띺@�Z��K+V�D�w�#3s��u��1���9)���a��?��-f��sJ�6n.����{H[S�U�����m��y���̰#D�
8�F�$`�_RQ����>�80Y6�״���I�;E'��WFo�`H6W9M"a�N�������8'�s,�*�H���,3�]c��3�A�/�LD;Ϫ\��2�I�����(�:}�����3��;.�a����$o���`JY���X�6/�t�C/ϡ-i���*e��"E3�#خW)K��v�C���>�Ag��*�c�9Xc�W�W^�tM�m��{Z����&(�{����"y�H�� ��K�$򄑕ܣمA��!��BCcz�1����x����>c���ѱ�"9���%R~���Sˇ2�<���亟,VŹ~Өft�s��w���e�l	������Eu��Bko�[�oV�]�FE�#2u��w9�Z�g��뾄�4�&�e������Q�~�S��*R�M����-eX}�o��B �*9�9M�{��<ד��E*>����~n%���g���(��SH�ˉ��2�mu
i6�.ɶ�T�����L�� (s��g<�)f�B�J�V*�s���Ϸf��ug�s����0�4�=����J�)-ɞnFB�O�����z""�
���6h��<�]�3�ѣ2�t��K�Jeѵ��8��R�Z�t[�3����:��s�ط*���o���knm�p�KLT:`��l�>�A�s ��%��ت �Lr�D�F)���@A�t�pv�T��{�$K�.�xI�;�}>� _eI�Q��6�)l4�5���Gՙ��LҽE�@�\-�nR�I���{d���֭�4���b��$�;���j�6��Boӓ��8��< �,��*߸QCjŌ�h�U�d���ː��Z�^���l'��B]��h�)�;.��/Z����dXZ��G
X��$
D.E�,�r�`D^���ܽ_���+-aa���;�U�B{!wA6����&?��(<��Q����C�n��.���{aEHY�g�'v��ǳԪ���;�o���x#���[E�ǽV�$*0�?���� "u��A�h�򟵰>J�B���e�=���1�#�E��V��o{N�f�Qf}q2��A��k��|T�zMt��߬���n��-��ܭk˽n�.y���G��Y�ƚ���}�>����IZ5��1�~�w9�*	 ��ˎ	 �[�"Ck�F%�C~�x�����sZ �m��o5��Z�2a�r`F�)��]qJ��w�F6���;�d�w�t�����My���P��"�
��Y�
'���3y���q��1��M����u-�p*����A�b�k"1??0h@X�����v'Wk�O��	��`)X��(�ͤZ���(e�y����`{OfLd��!-�U���b{@��k�j��;�J&3B���0#z\��3��M�����GV�{��|+ޔ>��R.yNDd���g4�K3�wcώ@����/�#+JHMQz��{8�17�3T!ZR�ߑ�J�%*�e��~I��ˢjmp�W�QB�ANj�0cGo��2�(|�e�nѩ�Ü�F�e�tC��Xh��jt��+!/��]Y�6�/����A�Ge?~`:������OE���F�o�X�4_4��;�D;�%�H�D}l��|�jnm��v����_b��g{~�i�T�ɿ�[����,/������g��D3e'4�dpj׭�����dWV� ��m��B��!g�_X�}~��h���N����{nC]����E*
�eL�M5fm_��,ձ��B|*!-Z���Gݮ��!m�We� L�2Ŋ����<�=-����8�Hܝ���i��4�_���+
�>t�4�I�e]v{{$aT�C�Uvx���	3á�s��dP��V}���?�Y�%�����Ź��������n�94P�p�ٔ����c���,"��O��>�"�;_�E+s��QO��R�~��.���<.٫K��[�X�c��L�->MG�_.?uBX�b�@/{E�����2 ?u6�5\*�
φm�B8{��N9�t���GŨ�_�E���Y��u��m3���rfs@�m熺ԕ�3����'&� ��Hi�-z���GN��7�֝�?�X}�q9h�&|��� �5�^��T�p�-J{h������p��A�
	�̦���@:��S�Oe��rf��D��:�9ON2vY'�<�n�9��Xܧl�&����C�ˢ��r��4@Hn��|��z3*6�݄md�<%L�'��q�>�P�����4�P�%�������|��6`�[���'�CH��ե���߇�[@��NL�����<.'�ՙ,\��S�-g��v�.����6��﮶�q��͞E���w��� �h#(PY����a��J��^���R��Н��6hI&��w��.(w旤zKc�h� �E��p�D���E^)`ϲ�f43� ��2���zB$mj�B��L���;R�'�գ�'��x�j����Qr������/m���2�J.v�������r:Y1�p�
����TpF�Bb�&���B�!���:Y�$��4�o�N��Մ��׈��\�����m�W�[T�&c���)џ"}L��f�p͂��D�2Bf�@���K��4E��~�W�4�z7�olU�F�������S�Jc}�#�R�f�b�Y��p��t�c�|�S��ʽ�J�L�;��_~fb�u� �go��Í��%E5�#E-xR[$��:�9����L3��A���E��$�x^B2���h��?��'\�&�2)�e�&� Ŧ����Ȥ ��-�f�	�s[��Ã�<��Ph9�d��3Ů�&��*�8��)g�J�<���*����	��G���:���OW�%�QS���ш� �)��c�3<xv�$�xSnm%! ��D�$���%�+��?0����:�?�a���� �>{
�>���Ԩ,�e/{�m(��#9�<S��z�x<�CM��d�-���bN�I���(���&�~d�$�Ƕ�{{�-E�m���֨�?��Z���"K�W����۰R]��)sh>o��������j���"�.�MS�Nnf�_��F
���3.D��lt)ʷ��lN���f�8FY�AE<�Qzē�n;�rh*�� ��w��5�d�(h��6B��޺@�x���*�R�y�_��m� ���m#�,!�9L���g�9��#�v�3L�^�Qm<b�y���u�嬅�;�L7��]���4�ΒM%hK�B��G��A�}|�����ڍ�68�nHT�:S�J�̳Ēy%���`�ȎTF�ٔ�3o��YHӚ�/?����N%�AI)Xy*���1<k�<��_��k�i'[xi&L��"���I4,�Jg�;]�����&M�Ba$��ؐ(V2��dᕥb�'i�hw��+����y�Xg���4�˸X����T�\��I������'<Otֺ�lf��l��lr�z�ś��� ���@���RE:�|`͂X�f������m�4�cb��>ZC�h����e�RV�t; ��#�Gٓ�si�\�g|����"��)tN�^z.����JW�4s���^-}�p���έ��=f�dԦ%�Gnx��W��=�S�:�R��|��J�ƞ8֡���p�sP��5w�?B�E����B%R�gD)H�����#8lQ2,u�G����5�\�S^F�"�!J^�r�^��m�OL|}�ݔXzK �H�[�����S���������-ՖJ�'��d���uV���7#Ko����2g'�.�H�]���(�7�;���c�\��$�"� �9��;b��D�S%�$~Na ��	Hu�T��Q)pֲA)y�����i	���_��K�5ȟ�	>(�(�m���BG�*%���8�����~��C�Mu'��h��.���Feh��������<[�����w_ �OͰ].�w���N�C�G��Dn�`E�k���S���	-���zs�xY��h*�O�V/�Zb]�qo�^���\p����ą����;J{��g�6E'|@����U���q��U�!+��4�y�=Z
��Z�����ʩȢ<��y!��c��v孓Λ����]�'�|"���xrn��8��G�C?��ŵ�Ewg�0��Q���qD+�uJ��+��(Q�D����+O�MELs5(й��-�I�;����ԜKڻ�,�7�wo��7_{I�=H~�>E=�)������yn�d����1E�m��|B0xN�@%�nk{\��3:|W�$OM:�__�Q��4����ƣҼ�.)�qI;r�9�f���mT/J��WW�rdۍg�Ä 	O"��H \��6�_����GD��(� K_�����4���g-���wpHՐe+�����s�A��6���?'����������O"�� �}*����2�k2/���U��Ǵ��l%���2	9&+z0�7B)����r;�蹷w
��f����DE�Q ��\�~���J����D�#TI��$h �c�0�INjWX�Zt��ѯ@��,rR���D��'-�pk|��F-�^��(Ø��5k�ӣ�K����k9m�g�}ȋYҶ0�
{��xr��Y+��@g�Ď_���#�~K�M����ٹ�@n*�������m�0�Sg9��XYQ��3R���o��"wԇ��UD�,�u?bW �&����Y����5��ܬC/��`ϻ;*#�6�OH�Ռ�G��(�%�=0��3�e3{�e�!�1G�[�Un���瓘S��
��d�-��D#�ϝ'���r{�4AX��fr&9s)�:7�M�ں-������1�;.���¹��QB�y����i"� ���7���Vx`���[F�7~�?m��m;%�Fr/�U��� ��=`�~	��b&'�yM��0ڪ��^�s��U�� "i4K��A7x�#�2F�o�Yҽ
טg��dC��Y��I��}n/}ɰ\���k<�.�!$K���{4���AP�s����1-'^B�5ao���f����ȝ�a���i+�ꭩ�!}O@L���		5]�m�4=Ԙ�iqBy���X4���G�(�A�����.�� **q�G�N�V4箩f{bL� '���3=����Z0!�'���*A�R/SEU��W��\2��r9\\H���X�������a��t�kBN���5��4���o���l�HlCn������|�d���f��:�g)D4]A�a�T��,(�&>V�$����(
���Yc���`��~$;��A3�]������C5�����|�5������Y��D�~��jKt�v��,V�),��hp��gvB��5ϒm�f����(W�Z
"�-��OQ5�'�b<EM-��8�-�M1V%�?�e�7�Wi�;"2� :E �/x�M��=�p,Ti�D4Y�d��/t�4\6'E��p���� 	籣F�D��"'�nw-���LA6��%���3�����xw$�A� ����_�_Z��;h�?�+�C���b�2��]Ap�`]�H���me�ؑ/��m���s5�*9�'hhG�����F,vY9"�.�a׶xn���M8�" ���y;��~��O�8Ax֭�:vtA�i�ll�D�z\�c� ��h<[�D`�_<�G�H�&� a�/?i�@۱.�x)�M��솢��Z+�^�eԽ���|]xc\3�N��� {[Z)o�:�DJ6y����b�7�w�I����
��,)-zɷ
���D��$Nĝ��`�A
���3�Z,{�%�l��r���؜e l��ن���Lvzi�z#r�3v	��\3����o�Cr�K\ã��d�b�	�b�7:v������I\�%����0����:N9b�>H�7Y.L��%��ӡP�(5�ڴdyϕ?o��O�mT��}3�����/��k�ЧIIg�eXc6|I[씸H���=�BC	���h�X�Z)�a�Hۏtە���r;ۺ�5�"���ߧ&C�ِQ�f�k���q䦱�Y��{WZՁ:�w���/��V�hտ	]4� 9��#���U�1D"Xe�X{Q���;Mx4��Δ��k4���{���\ڂӭ�W"�bޥ�RB/�o���Rn�ڸ\:�=4���$�h��`�VQ�F�v�3|�1I6"Lӂ}D���&v�*ĕ��S�tzvНP��Uߞ�qI��%ȍi$�� ����YkJ~�goױ�T��Qx1�o7>f�M�,o��S��Y6��&}3u褧��h��T�<�GHx��5�j7��T݇�f.�x��?���#UE��%9��^]�1�C��{��8�-���+��,���P���<@6��j>���gfH�A�$(H8x§ȥ#�7q�T��n�!%�R��U�V�5�8ݪ3���Ϣ�z��;�xCu.}�k��q�7�e���[�E����i�r\�9C2[@�D��%�Cf&�W��r�G8�A���|�v���Ct�SCQ]���Q[/ש
�1������t��"�fa`�Z�nK�,�6�����9V�b�d�!�3���̴���\�6ཊ}>MyO̤f{�GXou.��;��7jP�60l,�_l�ՖM~�`Ly�b]@��ѡ�a�gQ3/�~�;��MmsԒ QQ!]��	kZ��g~(Q�'e³]���@Q�R=� B��;��4������3~F�m.������V/Pa�BD.c�{l�����P<_b�:�5��w ;�=DB�6fJTW���YNm�[�� �p��<�VL�p�1��f>k�@���Qa���!�"�����9_=dO��_y�{^��Ù9��E�V���Wr)Ȍ#�[ע� ��bj��LX�����l`[2��?��1���V��	�7o	VR�Ԋ���.��d� B�sβB;��r5)��0�*,&D�&�q�H�R�_�ɜTt$G(��O`#"/�}�i�p(�t,�z��9Oݭ�����Q�}��Fʭ}z\��V2���0N���}>���ŧZD
(��GN�pJ��-����|)o��}�/%��{���W=j�=˒�LX��n`cO�h���]X_H��6� *���{)�Z����+�)u�_3�5Έ%o&u�+��9�Qc�7�Ixڌ�3@5{w�u4�zF&�hrЇ0��%���� xd�\s,ICy�^h���x�nq�Ҳ�Z�C5����J��	A�(r8�2/��z���V@�*5�����G�y�&��d�
��1����,OR�v.%���P�;i�'"⺎i��ɤ��m?,4ޕVݜW*ѥ��?j����T�u�-���t�k��:'F��g�����h����W�Q{l��6���_�O���8=�D�RC�jz��E�s�8#���y��)����\����jk(]�!�@���	��jgL���,nzB�l+� �m�r��{���:7�;7�5�� Z���uP��)_B�P��ri���_P� H�OdX+���s>��I�ɜ�����vg�.H��p�g=�����@Ew�y�'����g����NE�aI3���}�����%k�U�Yϓ&`�+B�P�fߏ<Q��MQ��T0��K�|��9�/����񏆨����~&�g�`�[#'Z=� -�q}'c�SS�hP6�������U_tOHx�g��@'+Iy�l�����S�x��-x�Q%�H	�$<�P���v��U1�m��-`22X���"M#uB�%ijm:�}�����(p�͖��YIhR��ؾۏ�ݑe�>{���ߦ:~�e�δD�[K tx-��(�� i���1�5*<W�}�	��p��/���C㮞+4�=(O/u���ѷ�\��� �-�����%��Hdj8�}�@��|�K��%?,�h!���w��8�h�Đ
#�y"e�w��Jj�ܔ�V��#U�P#d!�zP�|l��g,�!���L|8���˽�L�����敌qysĜ��M��	f{u��T�M?(��(ĢU�v���JF��HMee��
��{P�9"��Z�&�c
,���F[�.j��f�=*���'�}j^fزm��Y�遱��U��{j2r?�=?G=6�e�I�H/d{*��6Kú���u��?:�̝�������ն�5�'�\��#�[�f���ҍ�[�6ɫ=��HYI��ۈ��� ��ǫ���������P��V�SF:����z��ի:�Ή��?g���~z�Y�	M네�˳�:g��gԉ	`J?�]t	�A�RSi�w\����V����Z+�'oJ�����X�Є�C�$�ʚ^-����(�	��t��-��͸0�j�����~c`�[-Mc�_SBDh�'�F���
c���p�zI]#�
�-l~��k�3��6�ǐ�ڳ��z�MgL�f!�b`ˎ{s�d`�=W�/���������i�9?
��-Ks o2����s�`�yR6��X��M�������ၡY`��&K��C2#��h3�M�X8���(}���Q���o���I�-��M^XP�
�J;�	L���@��S�����˝��e߲�X�)/]�?d�P� �.}e{f;��ȱ��GO��nXu�+X��Y��P8���L%/wd˘l�Y47*a���l���h����O3��&�D#��Jn�\t+�\�ٔ�Iz��Q�#����M��w��I�{��s������ϫ��d��3���&��rh� �Ycj�t�6����������	87�)7;8(5��#ܲ�g��p�p�?�A!pP��Y����1>��k]q��U��O@���W����,7�5
��]�<h���lgz��7v[�W'��-ŋ��ʐ��}��
��(��%���0*�Gd�8��=*\�p�d��	��q�7��Fxg:`��d�NpF�M�B}�5�-�]���l�c���c��F�@�O�Ҟ/Kt�MJ�%�X*��W�@�)o>ޜ������wG�ٰ���
�OP�\%�����_����� ��������A-�問�����^��A�^c�Q%�`S4�ɧQFċ�H��ú�|�xUbA艩��u+��A͏J�B.Q��g6�y��@YY��/�]#X�
�X����;z� �X���KF%fS�oJ��Z�>��w�53)q6(��v1[�c����Q��+5Ps�k��m�zA�tC<c�|�q	�h�jH�xfV<Ƨ5OzV{�3zO�@��J�~]�I�V�� �VTR@��$���#���8̈��X,��j8$z@h����,+�m�93��"����e����`(�.���CsRP#��3h����?��U�zk�
�ʰ��OnI�W���]R�դϥ*U�{�3�fu�S���_D��������,_a�;�3�
Н{2E���5 *��5A�'��ȹ�o!�a��H�#��FhT�֬]1L�pN����[i��������Q�p'�_��M4AT��M��!����N��s�vD��l�&QK����mՒ�ғJ"������(nZ�VEǗ����]���x*���l��<t5<<Ū���&\�/���n��h۬�|M��l�� W�#{�:TQGsbK2J�1
v�7R���ڄ���n��TS� 1�3|�I xɌ�|ݸm�H��fG0ȏțV�j���'���0?��M)����cK�"a�"D��a����{-���J_U���4��mXO���V�;��)z����JM�Tr�1�y�J���	��Pq��e���_�Meń&�4�L���9���Ȣ��VdrA��
�¶	��0Ze��KT}�{��W�������,�y��e6[S$�I��V�|֯��U��/��D[�&8R�ӸQʕ���}����'<K��O�����l;!�MsP)���f�ٵTj��Tq-b,��,[U23�P㓆��94�(�)��Ig��*�p�J�u����#���	�c�T�9�a90N�η�	�j���%\}xp��!�_;�ko
�x���G�Y�x�V��؟�Z���1�~t�BiQ��ׅ/!�L,Q�Z�_���=i�p��Fםmx��[�� �#�[��xP���Ҋ���M*�@��x*�}���9,�>b���?�c�ptf�,r��ռb���Ap��â(`El��Q�m�����-�ͽo���j��+1%tI����Tt�l����{���7��p�C9��1���7�}?�
�N}��(��~8��y _u�+�V�{�aO<�v�m�H�,0[�`DJ�g�H��MKpYX�\��nb�<�d��`W��`j�&�&+� �R;��f1�gf!�ٔ�ן`RkQ�(B�ws߫�t�"qT��x�vɚ�K����k�L�Jr+kh��y���q��h�HC��P��S�v�����Q���{�� �"���U��7���o��Y��U�b��]��s�@@�q�'᎒�VH]���|]�\*R&���Mv|��F3s�:��z�m���ͱ�g>� #69�!�l����NN��Ik=�O�9ֵD�
����������A �Q�ZP�`�#H{��U#}����U�-MLS�����F4�#�N�[�mop0���}����� ���+�<�]j�R��g�q�����ċ�7������U�nU[Y�낟Y�劣o;����g��Zb}WUC���t��g��%E�o&.�jN���7�ϥ�w�!	z����=nɬ#t<�Oa�0fS��H�G��G�"���&9k>h�w5f};'q�*�!���͊,8��DT��ݫs�G���y�K
��i���m� ��
b�N
�P4�p�To�Ɖ-�mO2Pުh�L鎋��nP�.>�U
i�iQ��[�^G��Z_�/\��[�|E����a�G�و�U�=-�3_is�ӝ��kGeL��y|��]3 !�dG�;�G���J�uBڥT7 ՙ��쾬��b���u{�����c�Bg�`�M�D����IoP8Y�U��"���M���P;�,~�*{�r]���#�++�"�9���X�(���n�, �O�0�6�!9�,	I�*H�9?��XF۫�G-r�X�Hy����A��SV+c9c�F`q��Ulu{���泛y�N�εJ���-O��,���&��؀l[�Ͻ4#�B/)0nK!qqLz� '���s�H0�F��ܟ��76�Ȟ�1�&�)��k��[�Ģ�����~��J���uJr��z��M
*��o*Ts"V�,�U�2��r%�d���|�ߥ��m��./:&�ej���q=���������A���	�/�����?B^�Ð�,e .����Vs �1�N`�	Q V;�8'�q���i r��d0���]�z��3�t�bv���<�G��0�,��;M9<TԴ�7+���D Dd=<u�}�_���&�{ŕ<CC电@M�h-J��kOY��E3&1�x`�3u�x���Z����.|�Wh�[����j�Y�
 ��=���W_F����!����Ͳ_"Bou��S�@�_o���U�=�����.��bJZ2h�4;���c2��`c�?>=���쓯2\��Aqq+�Y�����Vz�ΈD5U&�y�.?�Y�]t��3�����ͫ�SNc*��\S�)ʼ�N6�n,k�||��I�Hyp��]�n��u�{�,��2�-.��'E~���L����3����g�-ιC}�8K���h���!���:��%�_|���v��$'�yj�Q��Ifv������v�0�
�Jt��?8��xW�1��ʴ"�,��l��E��k�.?ZyB���BCa=�ڒ)��ʄ�Svv���q8�,�����y&�����5bAJ_
����bq�>I�rk�_c�Pb����m�P.�� 1q �]��t��Xq��k#F���9�~Ġ��y��<���Um�N��73��l?~?r�����6N���o�a�~xwɖT�kBb.u�0�2Ę���W"�Ս9�-����!����m����� ^M�H ��$�z��mR"ԔD�'���	_Yl�.�C;�+��I$�п�؃��m�p7��b��׍e�N��F����'��Zx�jN�+�И�� ㋟B���J��?h(��BJ��`B�̻�> �+ϢΩ�&�����~	�z���#�v�����"���$=���g�Q�!a�l�ܱ�*���>�d��~n_�w�V�bչ�qg�q�%
�ф���y�@w��2b�i������</����?�$68l�8܁�w�
��A���b�X��c?P��8�`AHq�z�֪x$�ș����$�i}��j��s�O�����r��@�f�T�.�N�O�����V�h���>�� F�T��/��K����^"a��*�\s4��1�J��=<-e�S�}���V7攡�Ӄ֥�C�m��`�ql@P�BR��D�c*�-�Ro������n���ě�z�<#� +���޶8��y�Ʃh�W愣�1�B%�.@������ fs!�T�$9�ӆ�^�-�!d�w#�\���/V�b	~��a yS�o�=p�x�2>x$��|�pC�jV�?�BOMN�q6�f7J3HD`O�[����ft��$�
�~��Ħn]�e�E�k�h�q������+��&��@��P��_b5�����{Ж�tV-�#��|=D�Q�g�"�ps��E=��hK4�i�;y��aD�����M���W*����^��m����TmgQX�l���!+���<�i�|�.�Ԓ��2��[��m;�l�s���A�CYby-T����Z1�K+�B?z�ޓ�����o�%7�U\K����>�p�|w��`L�����@F��ʞ!�`�Ӑ�恴�b���p:�?t_� B��K��Lԟ� ��}nl��p�26$
T�OYb)��Ww�&�^H_����EԚ�[:�(���P������͠�W�mt�P%�����ۀ[�>�0��~3Ԡ�w��E|S�9�7ºE��_��ji�����hep�O9?,m�������l��
��8�@>��N�ڃ�b�~�k�����矈E���R��r(�|�/�)1V!��"�����2BsJ�3�K�w����xؑ��?�"Gj:��Ɗ��?K$,V�a�+��Fb����汝�����:��L�Q�?��`�Cy��"�Aly��R^o��B̒;mw]��EH{�	Ԫ!<�J��aeF4o�D������o�B�߀<G�i)�ӿ'��4��t�買�$��e �a���u��m��L���+,G�WϮ}����-�/v��Ϙ4�V4�#	mN��l�$�bQ�Jy������v9����&+�~��J�1�3���/�q�F/n�֌��6^.2��],{�8��?y����rtk-��D-��,V����2wRs[k��"�>&"�`��p�ǈY�>h��TrE�il��u�&7� +���0s��Vq���˴�2�f�3�\2"<v��hS�61��eME�+h#mǸG��!�P{T��K�,�b��4��+w$����%��d��p<�R����k�ړ�c6A���X�!@��sV���cIzм��k"���z�\J�న��7q��q�N��Jх�6��zJk�j�h�6=R&����ք��ȮRj�r���qC�)�E�b{�δqk��(9���w��]��c�{W�v�1��&�����Q$]�C�x�v <�w� ��{#L���}���O��@���N�W|y��P���t���ޣ�ihʟu%�z�]��ʀ��������[J�XK���y�+,���z�WF��$黓�ڱϰ<���
�	ߖ
Tׯ{=����DH2�|�%�]�������%ډq>��d"0����+����T�&�.�"����9p�y��G��|f f��	g��9������9I�����q���5��irU\g̩pK���o�6�svD�����������#O3��Zk�z�*o�6�7⯇�	��"��)�(g���R��x��۩&�?#��DǾ�\U��?[*��#@ޖ�,$�wv]�7���6"����?�e�d/QNy����[�i��l�v�b�޿�fK�0p������l�1�*H���|_�z��u��+�`	I_�LQN�*�k<yt4��r]��Eq��x�:�>K��o����^$w�X�S\�M�\��h�����FE����vp疲g���j�T��/��g�ļ���Y?��Έ��(,����L�eY0�9N,�U�w�6��m�s����H1%��>��.PC3$=8�t1��ZR�FVy�y��S�V�{��j�z	"��/��W����X��8�Va�I�aP�\��ѯ%�R�V�9�8ؤ�q�$@�i��� n���W���[xU �+����f�a���}i�';ה�#N��}��|o��3�� p��R�s�uvy�xN0�y���7�|����Y8'�	Ր�Mg��9u���������nh�O�^�����$���T�W'I"�o�̵�jl���+�� �Һ��>.t$.����7O��uQq틇���h-YQb�L���z�9<�~��3`OTM�$l�M�������F'�Y�l�b�brn֪R�_�!�6��V�����	 ��y�:u����`,CU\~<��yo]��@"�7��w��蝘T<=L��4eV{9v����ul��%F�C�HmE��.�0[��b��x��[�i�Q2z�=��t���"��j�(�Z��ݺͥ�h���g���t� 7@v�td�W�;��~��}����R�Mힾ��ܛE�3�I�r&� .��{�=��S{	�!G������Ա�<����ZB���ú�o���0�a��d���5���D�2�1�Ɂ�d�Q`|}}�&]��|��Qј��i�Y�<���H�@u�l�Rm-�eɡ�oZ�
'P|`�\f���yO�M4��9�q���o����ApI�����e�*�p���M+�6���X��aYXl���庾-Aؽ<���~� ��Β��"��ѳ3�����%A����������yǙ�dp�Ҳ�0�� C�����j�8Qd� �P�q"a��_���}�6��J#�e�����,�}������O����!��0���kl�h�Uw�{�Y�	抔a丽�����x��&���L'`��$�*)�w��w�ǮS�=]1���:�t��|����J��W2ÝD���Ehq�螇��u��M�*k�e~�e[�Pșmc/�eFF��
�n��MD$K�A��Ft>̅ U�QLuIY���3Z )���'�Ĵ���O4Ȇ���BS�R���
cz�>�������������E|���`�V�ӡnc��Ȼ�n��Z��O���J��8G��̎�g�?Y��B��=���=�_7��bܼ�'y�fN6�}/&Yo	��s���MP�piGS�Z����YC��AZ��5e�m���Yz�Y����+^$A��_ޮ����
�3L��"�k��A��!k�q�؃���b���}&D��i�$�����4��GE[�����kF� U���ue�+�W4���۸�mO"�2��o�㪞���x�6Y�0���Rc�A�
ɧ"±�g�@���\�$��x��h������.,�k⪐ z���6�S�jf�,G��1��ga�V�6d9o�.�xC����y�:�A�zd�D~��.�V�_���-�u=i|��	�]�8|���)�unD:��߇�����?U�>M��>(�Cy���=�̿������0�>�D�VN�����N��ܷ��ÀaΖ�ڍ��75�,��a��#x>j�ZEO���s)"��	1��D�� ̻3{m�} 9�}`�+U\,���(Ò�e�~�q���+ޜ;4��B;T9xä�1'V��^i<�F��*J>!5�w��bS���T���1~�B�D�"JXj٧��8JSg�g�n���Jt|j��p��--�6�W�w�Iu�P%4*���2{��6=L+�z<�v��G���Z�G�R���yA�3Ez����!;�*�>�] �h��椪���D���k?�ho�Ar�Cy�;�ߟ&���:��1G�QSRb���J7b-�?�Ff��F���GY ���Ek�Ga�hR���H�ߍmr��EZ+�[T��yF�����P�lPt�k�I J2����?����%D�H�P8D 5��HDyc��*����R�ً}!�X��ZbB����i��N�����q��<�=�S�^N���~r	��6��}=�t�;�B�fm�9q�}�	F����1b
�[�g'�`J1�Or]�L��L��DE�5y��d��ܸ��7�xyki��7:RνAg��]8��ZL���9eE!R���]Wѡ-w_z	\�Y��n�WP�Z��R�����s����=�?�27~���R�'� 3��W� �@bFw�6e/�����i����
��&C����^~��G�Y��6��j	�,=A;B��Cw�4���%y��K��uu6���E��g0�����AKEr� þ�C~����P�m&�a���k��48x/k������t�����C�7���T��:�vKܡ���톒�Ȳ[m�]�ml�L�d��f{���3.Q>O����}�)��8����s��7A3�n��G,��^D�%_n��p���z����9��w�B
��w7U����(�l��OF	��AWC7-~B�6Awe�:s@k�M�s߫/d�%�$ 9��Ma*�y�⚘vm7آ��������F1S@��m��](&*���#u�΄�z��~�9�<�7=0^��ʖV�W12N f��^X���, ���#�@�xN������,�!��I1���^@ ��qߩz�4��Dw�����F0긼iD�&��A)��g5�\��u)�:�%����1�	�.r%CMI>���Iμ��q%����=����uR=�/H�H��V�hN�T�q������dd��h��8*:��[�����M]%���k�v������k��l����;ں3�?N�(�!J�G�p����V��GA%��b]�v*�TJ�T��kh���R�����\��|p�IP�1}E:�l���&:�U<J��&O#P�xD~�H��oɂ�R`y���9?��u�̲�������d��7�l[u�?M�-2)x5�wD��a�Y��+�Ü�y"ڀ
���:�푘�eF��8�.s^,����G���L�2f�׳�Dq�N[�1���jAĂ"��(�� %�Y,�%1��u��j#&˺";Q��*|�
���7��d�M��&����^�k���/�u�NSi1��X�g��0c7�5�0"�#�;�ńG+}|D�Q����p٩)UG��E�
�$"�!����d�X�B!9$��iDd%�1��hu}:U���f��+7��d�_OՌ\z���>!p�}����Ώ����3)A��`���{i/���oͲ��B����Ir|,� �UX}ZNs�X������(�q��)mSd �h�:��;>���MS�m�r�V�bq���_(`ZE�167�5y����F�a�b���`F��xO���O�ȥ�jWk8/Dn~dy�2�g�!�F��6D}�A���%�<�z:����Y%�Q�WS�%Tv;q���W���ֻ�Z�������.|��|�֦��\�" ��\_f��y��;\��d�)A,�;�Z�`˅�X����Y��3��N�М��2sR��(��K�<Tw�8��YgBI9[�x��M��q�z�/��w���u��W�J�A������wF� �eF�($�<bpp��=�U���iM�]mvU����)a��E '�����f𻜼d˘r�m���@�-W�$�Y�ƻE�)����l��D���*�����K ;G%7E��7qO��@�%��B��*9��m���i��z��:��\;�`^{[�I=S#D��{S��^
v<���Jk@h�4X���m�>�>2��ߴ��r�n"3E٬ΦK�'G4}�o�Tvܯ�g�JJ!
7��<ʓO���@�[:�I:5��2�<�i��k0��&RBz+}l �Fg
x���!D_������KD�y#�I����``a��]�;s_~@���S6��l
�`��aX������F
؞�D��eF�lX�-(C�������������@)GMn~�-�}`R��0>[�|c����Q���cJ�UcR���Q�@}̇=�2+�f��@��7�䮕�]�nnƔκ��y	Dk��
�xZ@>H����j,�D�h$���>wk!�p�X���<5	֋����smI�0V�jט��X�>�@�$|�#�EΩ�)��y��),�E�d���-
�0L�� �>�x"����A�c���'��6��$��S����Jt-�_�T��⪛`���40 m!��m~R9H���ծ��i	8e�s�h3k�΄�H�s e�e~�ġ�$k N��Ѻ�}kM��x���H����"*k�gݦ�:���R�o�U��6��F�������-� ����E�	�4�rB��Q�47��-b.�Wu^�%n�d�f��䏅�aaϔ��$���HD��2��m�)t����f"�������O�.��q	xP"y��c�>�oKL!�#"Cq���ޠ�w['P3��ʘY'	Of(��.�9�k�W�P�7ȴU7�}�-
�� �+T��M��hM��g�[�u@�^a�)�F%�5)����f̆���j�:ު��Y��KC
W(D��x�)ת*C�,*i�n�)R�=PVؕ@�Ȟ���	�M\�����=N�R��A�Ņ�V��#��T���6@,O�>�bb�5r��r�@W��x�?@C�����E��	8��ޏ�D�B ��N�db:.9��a$ X�\Cw/���_� ͿJf�O�{o�?���C��ҮM�C�8!����Oc����=��sT!���8p�9��Q�aHz���Aw�3~����S�\ܫv��\3�p�\�GD��2�ȢK��A�6�m<��x.��(��K��}� b�u ?�h�]>Nd�J��P�z�X%- �-�+�D4�&�B)&�b>K�h���J�u�����j?����7a��U�ʙ9���V��h�$%S_�#��U�Y�+�y��� (�δL����c���������l��2h���CʪÏ�R��2Y�����S3������SSiH�3bʶ��X�<@����Qi�q`(Wy��X��F�!|i7��&&�B'?1}!�/�����XE�Ѕ�U�r�L	�nS��0���UГ�MSK��^i�u/
���_���n.3ߎsu�D��e�B���.����A��Q.��9��E���&�+���ŃYSZ\ZNݠ%���f�����A)���&���K�m.��"�"�}wI�[�]��\��w�����'�u>;�8����];=#��6�	Pp�h���(��l
6�[Eb��3ߝ�ན<1�dnt�l��k�XU�����_ҔV#���U.n�Z+�П��]AG}��ʘ �0>bk{LLo*�����G�Fs�ɩ��%	>l������`��rG�{�ͣ���¤+cƋ�%�%�Є�QBBL��T����gUSAR��鋌�^���"uLe:q@c�_h~�/��y+��NAa�C"c���xC�N��8�����x����J��',��pz��d5�.���_����^�.�VX֌��t�7� Z�Z3׺D��#��=ސW�#1�\���G�A���)/�4�pva|���������H�� ��ؿ�|�������҈�!8���G����K�%��3�<�@�i'�0ϸ�z,�G4��c���l��\O��:�~d��)�( F(8�C+ �avJ/"�L��۠KY(��N�oP��E�k�
�Ցb0����5�k(��<��3R48�%�ԝ�D2<+���+��z �;����P���ӎ�̢Xs�x�fP��ޭO���3oY������Q2����p-"e�O�8�'���L#�L>��1�AE��q�Y���\��M����D:o&7�{��م��ڱ��@�^���O'\�k�+�/ae8�}ì�n�|�����S9% �v�2���g�2�Sc��r+{��J��~\H�_����[A��|h|���T�1:㓠�Q�A+Ȼ�;[?1��s$��Y���l�!�Y?����3<|{�ަ��b������iv���.'HAk��P�������$��i8����×E�j7�o6)Yͥ?F�<0C-=L�K��%�ڤ���`���v!��Ø��d*����ׇ�
^���a�_�9B ����x8�}�c�mS*����5\Q�4?!�O�R���A��
�|W��串��R���N(Šl�D?\%�ͮ`t����s����/����yr��G���?I��Z�,���(Y��*^�de|zi��o�{'�2d�L+��� f��v���df����gn	�Ƒ����>��M�3v�����q���fwմ�V�L���H���ߝ4!��3�3��w.M���_�#���f�̪���NV٭���:���+x���Y��s~S?o��ǎ�W��tW�n8���튦��L.N|<W�/J��1�&�Ag��bv��4�+��M�^T��C�@��.�8T�s{['�#�{$�����Og�@�� 3Db\ �1 \t�/�L��Ϲ���R�0�GҸ>b�n̫k���A��}~
g6AX��̚��)$�Q��R{�R�e���L��T������z���[u4��4�2Y�|�ސ���_�ߴq!F��߷�1P����{�e�!o������G!nRr.1���c�H��i<W��F��V�tJ�V�.ϖ+��Z�%�j���B�r�=�:��u����S�<�;�9��m;�l���
�oN�z#p����t����\�-͸1Kr��a�v�6�'���3>��yh�ΕI����l���6f3�5I� �ߙ�kW���:�\M�qE�,���Nu��_���K���юYk�<0��-ə�^������aoN<�:1�U��1�44�he����T&-�'S��E�s�aI���\�����Ө����=c9uv;�Co�I#��(V'������u����{G�j��M��f<���1r��E��YgʸpӲ���� i1��,�+<����I�
��7?����"�}�|���D�e����.A�Ri�`ۭ�Z����K-!U��,�w��-��Rw�d��>
��5y�C�e�@N���� ̋���X�eZc.�8N�U Z,�R��EΧ�J��Z��[<�t�7����F]�e6�BLXy<fu#��A��5y֙���t��z9M��7
�Kmg����:w_>�Z�P��̹ݔ�O=t�l��wI%�'g^y}�K��q���x��pF��ay	�lː�rPĞ��'9����w>�ǠOmVڣ71���zz�ҎJQ8�Њ����v�֒�u���@k8:�<k�(�q�d�b�)�����Jj��Ğ����&j���2�E����NalN�yNUV~_��c���>���&���ݎ%���ʍ j[F�P5�C�㝆���ZÖQV�ɣܥ5m�4���ۯ �O6?����}7��3�7��57�?�)�4�{��fj�03�u6Fmy^
��N�7��(;^�*��X��4�
�n�(GY$z��r�a)�Z�g��.�M��\�O0CfAWB_���x�Z����U?��Q�I�4�������}K2S���X ��@l<�����'��TM�G�ߓz
��~�4r@#.Nk���9��*���s�ʱ���5���9�M������x*<[�p�����ć�~�c��x��a�&�e���=�&�̅`JǥQ&�w��)��"�YC�%��qM�����+:��}>���,�����[n.@nҖ��o�n!z�G������&K�b�*t��� ku���?&5:^��G�x�n�9��*^�MZ_�R��z'ѯZ˳��L>O��	m9�o^�
w�Zd�)�Hb,��R۩oeFF���M}�T�$4��>) f)���#���6wb��7� 
Ⱦ���CP1'�\�w�-k�d�oXX��B�XM@�����A��<���ŗׯM��/1gr��i�A�(���Sj�Ly����+�!��  ͓h�K߃y�������G0�7����\��f8������7"c�`Y$�������i��y�

�g�!�W|��-T�оb默3�-K��<y8� f�u� r�g��lOM(L�R��A��� �������۰��H�@��P�q��v�g��܉��t�K�e��ޓ֢�&�E��yS;{�4�I��P#B�����/����`�4�U�_��<9��bK#��J%��%ː�z*' N�[oM�^���n9��~�&�:tsfݣ�����C�X�?5�H$)� ��q~Z �z%����r7"iQt���@}�-^H�e��%��NV��;5>��S��t
ǟ�g�Ѣ*Fq��z'�n�x  W琽�瀠�������=dҏ��, ��Nf��J�nB�P��s���![���_�[1�[CKtl;:6�?#��3��SQ��P�US�A(W$����> �DS�AQ����x�gU��-��Z�4�zغ,\s@Xy�_�̝�[��o�a{���SGFO����c`s9n'�<.p�>����JZ��X)t�X:�/�t~įPa+2�'bү�c��`vݾQ6�3��"]zA��?c��2/Od�_c9w�iD��c���|n"�34�B��B.w��/�_��wĞa�3�j��w�T�E}΄�};�w��Lۡ����2��_�h�5E�U�2@}9�����"�~�;Fnx����7)/��k�9P���D����c��ݵ�oG:��[A�
�L'Am	�rx<�_g����o���/�a��;!m�
Jy2E�V'̪����������T�X� ��'�� '�Q+�6���'��-5\�f��1��e�k�&��}�,g��5�I�'�pհ3�����J��Y?���C����{U�FL"��ZF�pt���Jf�C}���Ӻ��_cv�Y�[�ԛ?ߠ4��[n:��/O�L�R�Ѳ�V�"�	Uy��4�kD\,�Y�x��z����.�������N����C�� �U�ԟ.��9g�+:O���^s軏�L֕!ȂB�� �4{[����ͣpq��uR�@�$�a����flB�k2.�����I�����̵����J�G/�)f����X���^'�g��^x�[z�֩�GZ倥�NR�5W,�R��Q��eL�Y.L��P�6Њ�H��8�A1��Iǋ��e';	!w��è��0	�_�1!C-�$���>��З�գ�
n>C���������ȁ9$�������u�%�z���Ź�ٌL�y�x��z��~�gf�Hxbv���ȏ¯;�=9��B���s\!@�ś	!���(qE?pz|��K.������s�Z����.���@�)�s=Fq?���?���3b6�:�ɬ�gm �_`[@�*pK�c�@P�G�F���=�k�-��~�%瞷6�>0Ĵ�$�bE�1�S=�Fx���vC���k?�xz�ӴL����S��`$��dZ(�n�Iv�RR�v\�K�7 DK)va��it�;��z��M� '��2�XHw_�)�⳩�]�៘��xlc�-�|��oXw��N�ԅ3I��'X��u$����o�S��'=��1�^���(Y0�:b�V��H��Z���x����|��M6��}��^j(oC���f���� �DO. ��Ob��ۀ�a�GIzGdco�$я�-�2QӖ�(��a�Y�e�M`Ļ�7����ЀZ���A����M0���h8�f�����&BRǭTM:
�LFɯ$$����3R�2}Y���|����o��+!��Jܠ���۽���(�5�B1��h��XTSi႗�>�y`��!W�n e�n4*��T�t[3/A��6<~�T.<R��E��QH.g�oN3A\U�J�C؊M��޼�&��Պp���c�1a)
�SE���{�
�B��G��"�J��]|��9�Rj��4xd�1/c�MROF��aN���{xӿ�#T��d"�q�V�n��F�5�D�z��C���{�d�&ZV��v��E`��Өh�r��e���=�]��x7T�bu� �	��%��醶���k�ԍ�0�0p�@�w�nW��X?Ǥ�AG\��E��:aQ�v�}@�c|�k{(��?a��O�&��yT�E�%q�I5!uW$zaOE0�B3C%M�W���#�ZTW>j�o�Lh�nf�N�hW2K;�+wC˽ s{���Y�[f���J���$���/����g��*�6Y�����.����D,B?'��N�ʧ��jB��2Xy�m��p�Y[�q�l�q"�/�z���3��A��mF��ɪ����� �����䕪�)v-;���ʶ(����6S�y��T�3 �}�:,oA�P���h(X����K���9���e.��Բ�� '��8�Q9p�i��/<"�ϬQow6�����P*�}o�7��z�E>�&�Ɠ����!P��|�)O��ϣ��Q�`��e�ZА�5:�����ro�Ey�jb��L�� .��3\Е�X�QW�$O߰Y��0�%3̼<�GẬhu8���S�bp�@�~��v�]L��v8�|��V��f�A���_�� �q�$���];�H=)w�H���Ko���P7��/��Ԛ����~�k��;g$_�7$hռҷ�I
�]}���Mc���,+����0�^�� ,j�pBD#��W�f�,�d�L���F�,� Iǌ����
pX�-�3K�uM�p��ތs�%B��6`�!�'�5)����dM��SG���D~��?37}e�a��dP5��l��{��ĺ[x!T�{��u��t���E��b�,}��ә,ݘ� 
#�S�o}+��Y�y�X#%�r�O�#�+`8��[m;��談{|���@o��1/'��_܌Y>�}����ȵ�)���>��� �^!��M��3�6�c�Re=��e�1�|V�S�J�G�|aK����n� ���z��\Ć�Z��}d�,��{�9�G�~oG�f�*����>�}���ㅳ(�Nz�L1=�{z�{��DJ��=��u�w}��{�	�vzL2Qs���&}�;�]e��g�����Ti�#���+A�<�(2��B�N��S�ϥ$T�U�?�F�l��uT��!>��ߎ	�Ӝ�={Iv��U�}�����q;���$���)T�(�^Cpf#p�sc-Ct�C=A�w�w��4vY|�e�>���L����`���$��y�ʴ��{P��,<j�՘��ԗvz\L�����s�>��Fפ҇��
��)�Խs�4M���ީH֙�A2�伣}6c�cs�9��I���r֐Q16��淵C̬W8M�C`��C�b}����eT"�ݫG�z0�j�"B�q9�������z�ˑ�G� �z�Mz<!N���+O/|�_3Cx���0���7.���4:�����j��k�$�yz��x�*d����  :ꆼ|�p�3�g�y�����<C��d���l>~��i���w��?/��$=5�<t�ˇml�M-s�[!k����̝·f�l؎FYOz|o�l����f�lz�  ���y���e~��"�P�|�{����+�1�H*�݂�����q{��AV��<�oB���<��������RV"�m"y���8���[�C��$��M� rR�hVMa���q
��}��|]%�H� r]N�}-�UVm�O�f���@�T�fJ�ayx4]�#����r��[vھؒOj��ȡu�M�)�,%�}���{�@.����x�!�����f�[ا���yA3��� ��-�'�T�:����{F
J�F��
��}!��*���-�8m���|
Ɍ�/���F�F7���E?�c_XZ��Vgf�p=���.T��c������?Y���\	j��loE����&�3��z���V��I6����u-r5���Kq��!�A[�S�'gza���U@]N��p�Bh�L������)95���L�3���a�(�P�)YQ�"������B3)����j��`�	)`H�H�G� ��@�9�"�)2H��|�lv��&3 ��7�ٓ*4���A\��]�\0�`_1�A}�#���������U��쀈Z$[ēZ��[s�߂R�K�&e��'�C�J��PY�ӈ��c���4���������%py^���8EY��0ܷΙ(��NC,�g"���JԳ�?��H��x�X~���;h��{ԋ�̒�]$8�+=�����+�����.|��rOBhJ~����{#<�+�DȐ���)��� u�G���U%3 ���$Ȝ�DwW��EƄ�/�p�ҥ49�2�܁C]Ac�8���ȟ?3+�n��v�(�e�o���&ǯ6f�����5{}�9H�=�?	����g�y�2���#Niï�M�2Y���� ���=����O�K� ]Lᷲ&��qt$�铊�~v�>��uT����w�I����N��>*!��hL|�f��L"�z$(��0V�C����K�翓a L	<i���%�D�+��䫉����T������er� D]S�J�ŧtHW���<+GI������5|��iP���v�Hy��i�q�nxُ^]�)	�F>�c�����a�2�@<����.k����A,���V��xaDr&�O�(�E6��z/�%a=�15 5.7���Ǳ�!Ds�[A���#r��A���X�iW"1�K3Lk����kG ��ɗ�2� kvs�H�r� ����s�������F���B�2_��&�����w��)��jϟŝ�?;���YA�������G����iS����BX�9\�InՋ�y�!R���	
Ӈ3�ȷ����]0�̼^c�(���Y9H���3������u���h��=�:*ð��.�Cأ	],��'�*=4"�4Jl��� �.�5^���}o���G��<�����KfX�Zdp�Ou���.*�m�����Z
�e
�hiTN(#\��+��a�[N0
nksl�����=�;��>��|U3�&��h9�w��\�����Լ�i"n�T��Y�L?W���Z�8L� �S�r�j����
}{?$�^�/�r 6	�~����0$��\*lPԁ>�.��XpN`�"�L	1�R1)��F�vG��tpϚV�9.@��cxʹ��ҹ$��Ѥ��J�}u��v���v���yW�C��{��{��'��9�Ȟ�H=P\�⬯F�>��k7I�ɶ�b1�[����œ:��F	Q�3a�eF��ģ���X�3	����7ѳ����3��3/:0B��;3_�0�����c��d����5J"�G^��dj�i.��ʸʍ�!�^����yc���5�Fy
Sxs>��֢+V��H�BgG�l��S�M�S���^�XėK�l���J��ߓ������Н��j
�}�b���[�����������D=�
��Z�=^����G�b@��g�cu\��`=���h�[-�P�ϑrE������D�B�X��J>�9H��"O�� �|��W'n��8c�r"�dS��U~��ޑ�Qz+��M����k@��5���U];ӱ�qg��8Ï48h[���H��2|jb��L�g�P f��XZ��6+�q������0P�ۄj���i*�}GU��ٟ��~f�O���yČ��}�N��/�CI�<2]cLpv�,��D·�P{����K$Ll�oE��sY�4�l?��^A%��r��x}�[}��Ptǫl]YuQ�Ń��i3p��:��)'ѳRS��Ns4�͏_��>�x>mKr�h����1ʙ���^>����7Ğ���tm��o��w�֛Q|�s�	qr:,3�?�3wq�=0�3;�� +2B�:�;���q�PK{"��M��/V��$ra#hBn8��oަ��� �	�>P"��#t�˂�h���]�m�<{�d �o���Em����m�e�G��CZv|µu����Ca����=��q�s`nE5���v��\���3�=��7}d��b�O���
����#8�j������ܞsf���K��z�&k�Ɍ��R�(���mL8t���]U�J$~@�'��o�k}������{�Wx1W���S'�n����߀ŃF�B\�]!o-��^�-��OcÙ��?c�L���L�}�1�)�c=��%�Z��ͤj)+�	V�X�5z��,W�*�ω~�����G|x�b���8ݞ��ֽ�C"� Dx[؁ԭ��i�����A��U����W �MFo�K��W$쫔�Y�);��YO�.�Kb��a�B���nh�S���렸���Vf���I� {C*j:�u!x�����|P;�Fp����C#��%M��l������a%dL���4�D�y�d�:�ͻiuh���s�<|ƃb5�����+�FD�>;u����������Sdu`r��[��FH�@�9�b75�g݇׃���&\��!$�r��^Z�o	B^�-���vR�F�7e�����H'^�:ة��h�w�L-W�a7%F	j�?�ݗMm;	?,Ѓ+�:e��t����z4�z	�i�;��b�2�4n�-�������"����):�ung���]s=q��]yB�"R�������z���q�x�	ۯ�E~���L"2�$+~ޞ�_oJe���MT�����gMf������S��Prf~��!�;,أ>�%�RQ�i&[6�-]r��X`H�$Ȃ��[]�wx�&�9Y��_�Ӌ�rv�+я�9�s�ȏՏ�W�|��ӟ5YA��'=G&��P�B�A�F;#z��~$�y4|]��e���Hc���{N7�]֪g�ԥa=c�\P�}[����pV���t�~MD�!o_k��|�{:��L��<ӊ)ͦ?�:3 pȣ&� B��Bp=g�_Ѳ�|�,�C��f�l�<"'��E�RA��^�mb#Y|�|و�~���@p��x\`
��ʉ%"5�?4��v��ض%m����wE��Z
~��W��*}���ɛ�־��o���hZ�y=�3�ۂgbN&��!����6tA7-�N���a^�K��ꗟp0��� ����|����@r�:s��}��yr�J����e|t.���i4*�"�K��I)�y�gzJ�|`(�-QTVأ��Ψ:6�6F'tRH74��m��#N��F '!��Ն�Dʄ�L�1_�Ѵ4�D*��ӊ����� n���x�hz��8�X�"A�L��7�| D��^�Fy������`�L*|n�.n�{�+��� �� �"D��3�!7�j��FJ}�{!�O�ka.��<8
W�����3o|��E'���PZ���*�N��x�������b�f���P��$0�4[��ƀ�� �C�'Z�*Zͮn�h���.������!��D�ϼ�=�p}fbK��Sץ���F�k����=P�(�\d��C�ɱ%�L@�%y��>�(����H`������"h�T�k�q��\.�1�)�kn1F譆���-�Wv��������
�B~��EE��A�$L�B�e��z��͡��k]g�ya�����>	�0��DVi���u���T㮠"���d�,�.�#�3��t�T��2��v�t��JVmc[����� ���d��Y�j���I���<�
褧B�_�Dl���"-޶��jQ���T��蕎���%�"ƈ}e��\�f;���K�:�;R�	T�b<-���K��V�=����M*�t܊U����O-�����/n�y����9؛�Oj�!hM�E���������Ro��J��kn���"��7}��6m���\����J
	t�\ŔYcKm����rל�8�r���˰2���y8U�݀�9���sA$,\��s����*)��]���d��b �ۆ��-h	�h���ky0Nq}lύ#q�45��:���Y�2��j�S!G6��ƒk!g"�ln^I��)��?ˮ�a7���~f���U7ĬFQ�G��-�g�%/�XL�������Y�3��E��t?G�A�~� %��*ę#��椛45	L��񄐊�Ғ���QH'�Q��2�G�ܸ��c�g�!�=����ޕ�B�ZE����]Y+l6l�'ɰu��n����C +����)R9	.q�H��^�c�X*�I(���U!MRK4��`�輭��>�Q8&��yqi�޿��ũ�%��#Ygx�S	�=�N�|�޸�D=T@�����b�Gݒ�맻z�g��rj�����|C3���(>�7���Ьߗ����ՉQ��X|Ѣ,���{����c���*�jvsvm!ŀ!�b�P�>��4[�2����,Y2e�uyG`�
hܥ֬\Kl[�Ĩ��j�%}E8�s,e�$~j�E��S����\>�����60�]���)��OF�o7'���8�c���P�P�@�q� �C:�e�P�u Ql)7×��<�Va�+�����m�����������4#�ס�r�`�LUA�6c[ڈ���b���*`#;4y�֭W�r�*�
�����3f�q�Gɋ�'_hm,��z\�I���υ�c�gQs��߳���p$��u�:&J ��cS��d%O /�tK��ȝ�Tg��H�H�V�~1�E'�UB�@�)9Y(�����R��z9C��(Ev�>˸���Eَg��tl\sǙ�W��JX��v�Q�"N蠻�ʛܝnwd����KS���Lp[����FT�N)�.n&�����&l��q~� ���#տ�0��>)3ki�����A�E,%�XP)���~L�3�O�r��;Ud.�u����E -��T��;y�8�v��T�9�HP�.��S:͵�3�54��޺�e��$ڽ���,����4}Iް����at~����)�#�n*P¤]�8T@\�hͦrʆZ(��)��Ѐiːq<9��o�@w4�U�p%1-��8;5<�L�#5��9u�+�uoy��p4�{�?w��U���>�s���᧝���S��zAo�K ��c��3��={���SS9��|��4��S��Z�
���o�ro�=h�}
����E8�Wϡ�����V8�'���d�Y����r[w=�&� y� �V
����\��okB�:�gJ˟�Da(T�>jU~���M�?X��G����Dё�?u��ta��4e��ZA
 m@���߰��X���x����&�R76�����۟���&�F�g"�K����U'��h���@)�^�{�2T��TD9�4�����@�x�+�m��TP'��Ǽ\��!���g��&1�֨?���%@D]��B���u��pT�vLY:�������u��	��M�׺��g�� �ǺTn��r5�c�-�.���|�����Mg(������.�ՃB#P���v5�����'��1�N*Jx�����ƍ� ���{���� �䁇�W'�r$����a�y��a�mF�����$[����GC׌�yE뛣�>c��)�-+Ř����s�����R<vcq���g�5���/�Ҡ��ھn�w���K�t����0�Ga1 �2�ߒ�F�Y�g�f�A�6�����z7�ɽI77�{�
/˅ܟC�Ͼ�`�>�^Ze˳���2T0�7�9K(0b1��Ly���{�f:��]�V�	�{OI	��|m>�J�44dyh�1��]�ܰ=a_���H�O_�0��2�X�AzN:��4`nD�ihV6���#����F�x�O�^[�.��Č��Ǧ���2�$�
�&��t<�(݅3sq�O��~,	▗On3���H��jPk���H�b�dN!4`�agH�w�<�~ .v��1|�q�$͉^��EX�7�JUgbZ�J��Dv���U����e��|�
��%��Tڴ��wƁ5���<W��)�l���2��?~@��ŀ%��ɳ�J�]���륍;+�&u}i���p?�,��)��X��Kd��a���Ḋ�d9m�m4���'ڒ@�_�����l4�_t_FwA�"`�{9Uy��<�Vp�1N
r�B~&��M;X<�L��}iScP�d�V�G��B8և�Օ�,P��o�u9�_��/W�v����)0�
��.� S�k6|��3� �SoMH�.��1ą$y���fW1��C7���4���.I��<s�儖�FY50Fl$XKԐK&X���"� ls`�!O�h>��`�h�i�6	,ǰ�i>(4��eXZ/�)mQ{{���G�|�ɰs���g��r�A�t�>��FLwZ���݊�b&��{�z�n�ɮ$/�M
d�K��f�I�;Y%��B�:�Ɇ���64 uC��f� �i�^���	%������jS,���3w�ބjt�o����q��i�bmJ�6>�U[�����=~][uQu{��@��j�fҋܱC�`띿�E�UG&��n�.�D+���͸�i�����F�F�~�i�xQ�(�ͣ:-�����,Kk/=�œ�����J�mZ�QP&�a���xEy8#DmVzAu�x�#�XRܻÍ�[�C�)g��?LW��)�u�W�V��L�i�}�'\�'��>B����U��<�_}s��	�{B��tp���)Z[�ۘ����� ����k�J�|4oc3��kKnږ���<(�TD|�o�9��a������L�#rv�ye″�Z'��O�4�.��&��ĆH	Ol���1��2�
*�T=�[�W6O3�\C7�����.�Q�E�����̾a��6"[aO��4M��1�������`���k��y#\�-���Y�g:�A����-�ӘW����Z�ɢn�O��%̣�)�u�5(��Oz�����a��
4F���KM�0�8�S[�M&���uB(G�������X��7��8�g(\"���Ք(�B-+0j�u�vzۉ�rC��+fs��k��Q����/�O'?d�Gl��s��ꘀ����-�+���+�ؙ���m�Ck�N43t�In���>T��[��*���X�u2pC7A��0	C���B������DV�L�y|�98��f��NꃣbY��ob��5rR�"M<:����V�<�!������ o�?��s^��8���_���XY�38-� 55��'��!Ҟ{e�H� vj\O�]ZwvI�Z�Iz�D��WSh[�٪sg���.t��n�uC�ǗG �T�ty��~Ɍ�{�o�%A����(g����ѓ��Q4��Ԗ�c�w��n�5�4.EH'�:~���g�!�E��0�Q 
���b����~�0�W�� T�P�]d�����;Rx��M��S��8Ũ�6*�ʽ)waX�<�Q���u�V��\~.��X��F��|I�[G˿�ͮis����WWmd�4L�J.�r]�v�,��y>��h�I鮔A��M��く���)�Sg�0�A�䕌�	_�8���"C��l:��VO�����x<6f�1���w�jP\��@P�Un�\߂O�㏳���l��7,�����ڼ.b�"&�2����XH���qt(�������:g��_���ù�j�����ɕܝ
]�����+�eT�D��1�>���31���kh�/!y�	���x:����3Hgs3г���d��r��k�ޛ�+�o���.�]�,0V����z�*�|#UuC��z�ݫYL-?ҧ�}M��⪓ȟ-����`�,!d����eQ����̠��B	yI�1��;sؘ��dO�7��S����*O��랽Q/���d��϶�}j�p�ۡ��8a�g���$��L��铟g+g7������~s����T����k��#�L�gPJ���� �=.�p�UT#0�6n�%�!��w��e�E�W��K\-��O�\� V�@۟��G�=~�e�*�"��/����!��K'x{�����aI=�:�i��TZڐ�V�h'?ި���@Iѻ��g���Ƽ�ԬXS3i�P3k����ɑ����K$.�����@{�� �b�}�(z=M�������԰��g���y�����g��cPYk�b���mfg4/r��;��LM�X)�d�룘����w���l3o�H�g����#�܆~<�������=
�W���(�<b�ȶk��$�ھ�i#e�ң����!��-�PA���� �y����8e Et&Kx:�U����g���1���@ &�����/32���JQ8��څ�9!$��R��NA7�޹b�����l����0��������L���S����
+Y�$w�<B~ �܅wm�h��jٲ,l'ݟ�N!�����jq���pjQ��V!�͘�;����y�����ݪ��,�����c�
�����*��"���D� ��QnE�1�yXb}��3�B���%aл~^�L�]�z3�U?�P@�?�Y���Նi�&�h�V��0�N?��T��P�l�)��>��k�y������k��B��͡	�9KFE�v}��L"�q�f���1�X�G�.E��?�p������}�T���\z�F:�P�X�f�p�n��C���'�P�=��?z4b.�uW�l��PsƺW�Yc�5ܝ�e���i��ǎ��#����M;��Ahz!��%@����Gf_�Rگ~Ij��d�E��WC�S��٢<7Z�l�#��M�UF(�d�J;�;���4�� �=ڶ8�_~�c���j�Xѯ�0�>�W;���W����g��YE���do�����ޮ� 1{6�~�����zň|ݙ�i�Z��`onJ�']�*;U.qe
V�樂~�{�3�K��ͯ��=QBӯ�Pp1�_�V��f�#��O�O�¨xjV	U�0L!*b$���I�%���xB%���$�܋�<b�u+]8׬f+�/E�G��L����.V��=l�@�;uL��J��=�gl�����Կ�ȱe�ܹ�
�^�9�~Ҏ�A'" �`�������I�2zz��YY->n}CV��Y�+W����mX4~�p����h��¼o������y�%a��*�H�7a8җF�#����7e�d�|i8���*,?G/wZ�R�8B��0g��`�л��~v�5���R��e���M�rl�x�O$�'�ˌM���>9f���=����i��'�pdl�7N���U�?���Y�S��7�C�O�XT��`���:e�����^n��'%����q��K_�GJɊ�/O�v倞�ujƧqO���V|�amn K��l�i�[?C�+<�g
����5�x���Js�� Ab�K��0}=�f�EE��IU=�oͬ7�Y��in#A���z,�k�w��'G�/����*���?�C���=A+!85?z��~RW�l�㳖Af���-�>mC����k�J:�ȁ����	����l����(}��r<�xَ����6
�l ��` _PE�ěaXn.��Z�����Oy�������E�q�O�Xt��[TqQ8���y6ԹST��z��)$��kCˑհ�O�Gɺ���Jڃ��t{H�\J�����.�Ρ����n�u�O�2���y_6Z�?_�� ^�(hB�2TPsۄ�e�"x4��(�*O��9Ȭ�`Z�	�{�8���B�k�ޚݚ�G�����o�oUٖ�X����.m4,�ݖ��$j�,��wY�G 5��0}�����َ3�Rk�
l�*	e��f8p-��Œ'`�M9�sNfΟ��p�0�����,��d�.7�����s=9��8�;n����Yq����%L?�����/a�{/��a�ld�<*�3"}X�'1��K�d�#��{�pXŊ����O���:�����L���h�"��~�q�&�I��z�F���zn�f�� X,��+vz@�6eU%�eu�����f�t'�#��`�mxb�V�3�9���MSC��'z���#x�=q^s�6��d`=���|��M��*Z*st��}^
&J����(O�4p�v�r��7b��8Uܤl+0~�H7q=�t�4�����ۍ�[\��G��?���J�:4�9Yj!���Ӥ~���E�"�$������n��e�R
���L���<�|�Y2��5��gy۰XTGb��q.n�9�R���K����
��F�q����b�X�S/
��rf�<�** �I�U��E�{#V&ǀ��<��I4
�!y�������Y��!����.K����OBy��0�F��W{^�y�iH�����Ͱ�A��m�ߟo��7�a;Ҿt���Gl9a��A}��������z���vK�b!
�G��G"۳YW9r�o��Ms��l��f�����&���FP����#i�T�d�c��	�~�
�>���\�J��@6��2���?{k�TZ�#W�_Bj����	�~����`�F�C��	�G��F_���v�_+�Q%ye���j�~*KS���^��}��T���?�~���T�Z��IEa �	Y/?Lq�^��Qй��Sz��[-1�3��D&B����O����2�v��Cq�|�>S�d>�bj9���RՍڍ��$4�b�+悰|��ZwH�Y���ȧ�L�O��=��^�8����k�k6�A��Ft�t�P�`�����|����xv_�{�_�a� ȍ_#��Ϙ�9R9����8{q����0���T�����֝u���^������.@b��xM�y�hP؎\P\�T�N���.]Yv����#�t��f�G]�U/�,+%�J[���j(�I%i�C����o��阞�?X�iӌ5f=[ģ��iU*�֪���@ns,]�I`��`q6۩/�5�����Zk�k�T��X��A��@*w����u�=�!U����!"����ġ��F�|�[����39���ѣ�=���ɮ�/7܅�i���Y%�,f,%g�e�|��ER���1��~+���r2�e�UT���d��n�{�\mCDbe��.�ڶch�Ϊ���c#���!�,�@.[Μ�B��,גb�ﱄv��*;S!p��ս.{�ަy$[<R�)Ω|EK8\��Qm�gV��&Ҵ����ʞBmAE��)��i+��:VU�sFr%q�K
_-�(O�g¯�����ԑR��L�v�Ldp�草�h8W�q��OTk0�Y�v+��ͦ�wC��}<`����V*Q��H\�C�qL$�=��/�(g�lC������{�Q��	������*�?�tq]>�F�`fQ\����;X�=��cV�P����R*��Ɣj�/ߔ�ё�Bl��.�U z���5��S-��G����hn��Ufs�!P#OS��g�0vj�	6��=*� ���˒Em��:�F^Þ&��췯���֢�@��;��Be��6���BWyo�zs�@'ӯ��B�h�}��K��<���� _�a00���멚}�?ƌy����v�&�
Ɏ&�{����xB�cy,R�m�#�rxn��ӎ�_	���7AC���uq�r`- ��X�{-X�l�c�^P����+2��R���F�f�I�n��o;U�8��յ�UK�("�t��6$��]�'J>`D��w�ȡ���z���Ȕ#����Jg�oTm?��_�P��vZ�F+��T5Iv A���|_���rQ�Z�CN�=[-�i���}��D��/Yk6���"Va�&��<��J��g�kT�V�|3��]����������$�����y�A��[�����BX_\�sX|�x����H���خ�a�l ?hݨ����-�h5aq=șEh�6F:mQ�ouL�N�U�'����� �<�8]^����nOR�;�دe�F3��|���US�ן����ѱeQ�Z�w���bi��Rl�����e�Z'����ŧ���?�n�<�d�Em]�k^O���E_W� gIu)%	1#��R���M+� Hԡ���
R�>�	�4b�Tё��^�"勃��`7ELg.�q|�l"0ٕf�L�Zq+1e^���(�qݒUv��#5��m��V��]�o�M7��L�s�%5���ً��#���{����;�
���ۏ��M��>0��;U)q��T��[�����KR(D��-P�,o5ݐ�-�6w�Ya�h�l,�	 rv���:��E:!>4k�7���	��P�\�OqTs��:xn�T����iw�3:�tMDs!L�ah�*���}^�Om�-aÖ@7��
cH{?fb��l^Y};O�=>�_}31Y��!ԫ�}\޻;���ަ�&?�_#��b�۳�H�!�Օ<�a�O���ˈ�Q��K��+�u�3�'�ql�	x*el�W[<��=��ͯ���D7Y�}��Fs�Am�������J_B�:ݠE���+_x���^�mk�G��� �[<+8�J��I��"3�,�G2���c��ӄ�e�1y���[x�r��4	#�s�*l1��^�Ӆ����5g΁�	洯_sԶ�8�/y��\��.BV�6��Y_�N�Q���츤�`s�4L���K��*zW3L�(��ް�
.�qL�	գ~|�eS/��H|�#G[�����M*��WX�e'h&/�/�r)��Nݍx߀�tw9�<z�$e���Gic�A��ء�a��CO�'����u�86-~�7ri��͒;��'Q'�dڭ#���Qmט�
��o~r
�+�6�e��A�.��F>��k�A��w��H��_�;����֘��'�o�8���u���mZ<A�I�!�J{s�w!�x\�?���Q>�j���N����uZ�!;\!���^�b�}��%��R\�{��{��{y,����������8�X��Z:����/�J^D+6��@��(��)�[<y�p��7��T�e0���dBROg�R?��r�7����&��N[�2W����̋Ϭ}�i�+/���F���x���g�M�����^!�����g���w����M>��#咐j��Zo`|��W�n�,�Yf'�	�o���H���>[����g�3�-�*Z�%XI\�8���1���JL��z ��7|Ѳo�~J�O��_-͘��=o����`�$¹��$��r��O�\��9���C�ª��T�r���7���	ķ&��f�|��%�����3��8��4�F���?�(�߿��e�L$kP|h����}.@(���9nsA�cD�<�C����Iا�(�'����n�W�Z
���9<�!�����]�KdF͐
>x4�n<�}Id�4��t����F������W�:�,��{���o&46L��2�H�����i��]�阵�H�E\�%��+ƷE=��� ��3+ф	&=\�2��(sR��IB����0��0�v¿n�O�ý�s6�MV27�� KGҧR��|�`���H��z̲a�
 5mu�~�0�s�sJX�˳V�1��dtE���9ļ,�6����!f	����N^�5�)fS*,@����W��x�����Z�Z�.+�w�U��ES$�#ix{�|�.�P_�\W:� ��39fJ3��	�"�k�A?=�=���"C_��V�g��L��,�=CD"Kw���,w�0- U�X�O[:�[���wSqSdb�^-���,R]]����n��C�qy����ˍ���m"0.�iqVAL�o�T2��z 
"�A����#���&�A���Y ��1�sYȱ����c�#5.=�[�Dg�bt��*V+v��s�1���ڋB����vyD<`�	i=���!�Ĝ)���`�K�[�-��ɱ�X�O���B<F��>Sc�;9�1�M�u���(�H���]� ����3M�@�x���W�������/מ\շ�%�@J�;U�8����T?؊C5)�� ���h����#_H�L;ԥQ�ç9�;��1�3[�֫\�k�� ������|�^����3�{��OyCu���N�����n^��
��Y��K��'�*��	l}�g����*���n�J������w��tx�6��rv�%�J����=��nn�UT��D)�����ۺy9����wɎ%���˔�\��;�2�9�< �0�9��KK�Dݘ�f�؎��Qc/�ݺ�cr���Oa!m*���Mٰ7^����Q�Z��F)��)*��>0R`�Z?	����39"O|��:@=N����y��q3� ����1W������t�� ���6�m#	d��S8�3X��E��\W�"�2P���:�ߌ�����2kh@��;V�jT�.j*�:��^z��gqi*ܺ��30���D|o~��KM����o*ʑ�w(�&��(�X��!e�Q�S�S��'��{d&����,��W�Wf�=*5��3�rʺ������|��l�~{���<��e���]���m}��񳟁j�k0�+ԍgc�4�:\=W�u��S��sݨ2t���Y������-���"L��{s��D�3���Yr�9S�9����'WwN&��G�g�l�RREN��}nA2oE=�����x=|j��W�j�Q�������<Դ�/*D��<�-F�j~�جM5�.H]\�?l�5p��a��,w�E���Vez�%�^'`��ڊ3���&�@��?��ZM�2���v����f��M�SF"���u���X2�M]�_�Kt@��Fh�N��pb#D��/ � \Ǔ#oE[	5�EfO�ԟ��y��f�Z>r�1�D�l��j��eļ�w{����������2�cZd ����Wv�!a��`Kj����T+�#�fqA�7�i4�\� Ũf�sf2������6���_��Ԯ��)	�����AB�I_��B|��<���;�A��W�M*h��\�Ѱ��yV����8x�{�+�CЖr��>��Re��Ϭpo�\�^Cbb�A�8#�d�9}�q�\��
1*�t吢k&T
3�!jj-����h���>SˀT����S�;"�8C��.l��`R|>D�H3$�>K	���N,}�[$?GtHh)��I~2����wОn�79^ݗ�;8;��q��,�']�5(�"*=�:>�"��*m��F��V����e��ZMz�a����L���2N/�a] ��W�����_���eW��p��璡ѱ��7�P�N��
���{��������v��(�:�;�*�UcT-;�T���wa�b��H��^Ϫ�*3�G�`�m�CTO�ժ��"m�L�hu�Ked����W�k�}γ��u��ͮ1"[����?|��F�����/�$��qѥ��j��.��+��
6��_�c����}��5�� ��E��X|�|������4��e��"�����my�9�9����Y��#�M�Mj>Spp��%/��8T�r�UZ��>	�~$4@Հ{���;cG3�Жd"���e���9O=�-ߟ�t����)���Z`��`�Aaٵ�4R=
��<����Ƣ�F���ڎ�����!-��U��Q��M~�xg7y�wzr��zy��	̔�sd��KΝ˛l�����q��)Y��E#�|XA+dר�(�'��6'�DL$]��e���v`�i�$����30@z��>� Ҫ_ʻ��>ʯ/� �������,i�,+P�*��j�J��a�,:�M�b�"t)�y��0Q�m�6��T������]�K�[>��^�����T%KLq\�,P�7��y��q���"EV�8Uf����l��8
NVɺ�u�+�㠧�y��;x"@9���:��-3����v����p�j�@���k��!��C���A51�svWE��;�n���Jeǭ�x6�+o���2�+&�X�,�K��fi�Y�Q�=�`s�����#�$5Q�����?�	���@/M�p7o��(gEB�[w�� t���[9x��yF��������.�8�7$ٽ\r�Y��O��h�����RX{s�yx(�qX�:���bO�~�0�����G��Px��Y��&6b��iM�`�?��7��4-�F8P!�j9�
����Pj�8	@���Pz{=$,U��a�F��B���s�l���c��V/+���|\/���u�[Jի���u����ZU�Em��i��[pZ_�5���+V�
i1��b-�Z[c��L��ִ[��'�����0Z�!_F^3�G����g2KY��1,��>�<'㎆���@趢ƷG�`������1�y���3/�W�a�
�j�<����Z,�;Y��⺏�Q��y�E�o���Ctu��%ـ%����l�bR�Q�`n��G� �!YR��H/9���jg��>}���:��a*������rڬz�o}���%T��?zǛj�d{�/��G7��,���^�xa��:y���-�[�;�6����S�%?��Yr�P²g &-$՚�;M�$�1ꯂ���	5���i��-�f�P�
#���
3¼)��f8� �V�V�,�j��1p TQ����ןˁY_��S�V�����R����$>_O�Dƅ0�}Z�y0^~W����.����yr�B��F6�??1L}B՚Ц\s��X�۷	`!�9��֭���;����hD�7�.Cf�ø+���<y��*>`a�$C!@��u¿�a�Zu���$ot!��I�A=AO����
#g�@��x߂���P%�^�3W��k41D�B�u�hV2��o)J�'h��q�ah67j�윧���18�x�����@9L�tt�VH�*!���p^z�7��t��|�Z�uH�!��Ω�et�P�0M��x6e0q/ɷ�K���q�b��+��J��'�t>G�{�� 7�R�#37� 4�A��$���!���&��e�P� �v#H����49�������X0�>��D2���&�C�D=xU���$�Q>�j�~�i�p���(����j
I.�Bz@>�W�y���B�L3��X3�};�����>�$���1����c�f����sy�����⭧�[�Qˡ�!<Y���d��)�"Af�������\����j1�	=꾋��A`w}h�,3�tY
��Y���-����j�z)������hh&-�1��d*y�
R�zj�{��-�Z7Fۮ�&���N^�[UayŌe�*��5��yǬ5vP�0�޸Ӑ|-z�� 
��E���[�A���V?� ���o#C^�sn�y�O����⧵���Y�c^%��K�ȉC�QE�'��6`�k0�6a�;"��+�ԣ���)�3������'(�72D�7��� ���s�P^*s)}F�v�c�U^x%��QC���'~�Ռn/3�ϒ<�5�����M�Biѹ����>����3�W^��w�����y{�J���CdC�I��-�?��'ʴ�)#Υ"C`'j�U�����Y���F	wKL�U�]�� !�T��� E�6O�����x��:m���n��.AL� ��0����whC��FNL�洩��/��≈�F���e^�%w�3Dq|>���MjvW���2&�rq�G�v���\��j�t��3XFE�,�S�a�6`�?�&��^�z����a�Ȟ�l]6B�ZD�XŽH�쪩{L�%o�Duh�I~�*���6uf��۬�;���M\�p�!{�ײ��2��)E��^��K\�0�w�yn��͚_��`��A��{ؿx���HO�h�U�dV�[+:�����_�������/�Vr�Ӈ1���Tu��x�ºG(	����{�h�Y�]�>�;�������T}�\�T�t�7z�֥���5I&��r�Vq���}s�E��'m��>�J?M;k��^����3�<�W��9x�b�hv <NW��
Q�����=�5ÅsP�&��Q�8-��A �䎠�q���lz����Z�آ�����x���A��E�{֡G&t,�����-���E��:9�F�Sa��e��[���A�����}u���U2��PMG�/�����s1�ْy���*>����Aw�F��;���z�0� �n��Ng?Y�5;�u�?�Yd�$��@A��F�w��-���f[S�V�఺���d-�z�Amq���[������r�Vj����$|�u���cX��Uq��p1-�#���(�[8]\�,7`��T��*��:#�n(H����MuWLo]�*��V�����ގ2����v߫}�ߖQ��FH�|&}h-��@�	�#5&��Zϲ@a�,���r�(��C����@�=��+�?Z �M��LF��]���V�ܳ�o���c �H8$�֣�c�CWe�m�
���/Խ�zE��=�&h�Zv�,��ね�[�i����t���ƴ���ܫ��\�s�^?J$��Ǟ0��Ag��-�z���Mfo�P������!��TH�q	�O�O�]k�@�gy�T��]
�(L��KT���ɄA�/FA��\Rݣ��P�S��.2��(�i�o&J �Ejg�=Fa�\����u.��Y��ӧ��rb�K�A$]vO����tۍ��L�鞚5�1��`��n�d�+��Ӛ�e�،����8>,wr���!m>��)H"�e�H+�%�^
�1)����x�Y�1�5?�#���H��$F�uO@��v�Kק��s@����kj׹�lh�3C�Aޤ�*xog@���^��i�6��"�ȫ����44��L��v~�È��=+��;~_��(s���)|(6����-�X�}n�]O�4� ���|S%�)�j��k�}�7��d�4�#
(����G(�Uy�q�iH�,-{��IHs�8�t3͇	��}A�A��!�Ph��R�2�>�����V�b�	M��2����K�!��̤��ma�g1R�D?��2ֺx">�!A��4�IP�|�9�4]褈׈�z�J��bpOҁ^��^(�;kjCGE��X��B,b]:��25ſS'�R�:��xR�w����.x��xc���T,� ��}�^��]`w�W�zi�@��94�";�gӛ���\9�&��BB����[>��{)�-����A�q���9�L��]�bVje��m����Ĩpvc-�������%���&�V�s|���\�A$E3��sX�.^�]��a���L��ſX
�"�aWrT&v���Fv-�ÔE=mŵ�r��yg�-eͶN��k�h;u�+�N��.��M|�׻���>B�5�S���6�1�3��dM
���Du���<�{e�/D��Ϭ���Å��Cc(Պ��U�/�/�/�8��	���ZL��J�I c�`��h�z#0��n&�Of�cu�� ����#ʥ�~h�7D]��O�8�4�8^��X,��}`vn��HwÚ�$�J��c�Cܧ���8��T�_�j�~�9 ������2,��F{�x
fa���8�՜0�B����of+%��L�w�'�� ȃ|*�gy�� &&�w��+>�+R�&Ek1';��H����I7Gi�3XD	0��O��q������M�]�ּ��-�E���yt���!z74�N�5�� ���yɀ>3b�B�k�S���>.ڗ3	��! g�]E�@���͌!�u6�)�ĨȈ�Q(��|x�p@P9:�[oC���р��>�,D�!�_!�&{2� ��<N�m�|B����;�[���]�9�b3�HWg�z�}�v���7�Kb�\�+��Ȭ	p�����b��%�\��T��R�����x<I�N�~Z�\�S���k�$.��GhM�>�M��b�F�LGSy�6]���m�|��*���?йP?�W��R���ms�|	�e�o� ���1ٽ�+ش��JV��Q""gS�-^����G���1���2N��S��ʉˬ1���	��:O�
T���p�<C�������LͰ�����#'Z
O�eXz�7��1g�=Vi�U�wܱ�Ц�v�v�
�r���5Ɩ���D�+%�;it����`��R*�eOP;���P��d�?楦�0�����Rǁ�uQ�/k�<�@��.[�=U#�wD��.��Ѵv,ot\��b?}���%O*��jͰ���V �k�	D�C��d����mm�d�}�W*���#�� D0*A5��֩�:+�Ñ�+V7�?@fln�X����)�$N��
�m���kѤ
�#_�i^L�}���k���,���A|�����(2�waf�p�s��ג����o��((Ǟ).YP{d�i���m�ڞ���6�������8,1x�I�>��j��D4�ծ4�Z�3#.�����g��3�6�:�>>>fU���'�C����Y���=��H���j�m�"ʯ�l�����j�Ӹ�YR:�E��\n�Y�c����)3Z��+ �q�E`\Hv���Z�,T|�t�%�n	Vz�V�A1�/��vw�`���l:�A��������g�O �H�q��^�y��o�iwо"���tJT�XU��P��v���J�j	�@�_�lΟ��	�ONF���tߙ�*��ͦ@�uF!GԋR+��� �A�q�3�!P�f���G��H�����$�c_ǌh�qͤ�v���Tα[+���'�����P.Q�_�UЛ����4/I[Ɍ������l�}��ͩ#�8c2$��֌�m�Fc�G��)���H ����$��k� '�0���SBɲͮ�+����.)q8�~���$7asj�C��oҝ����݌��`���Ų~��n��*�b0vF���J�>�͖b��A�����-p��z<�Ay膖�n��+E��	n�ض����Pu^i���(�f�>���uo�=�d�H<��2���m,R]�<l�%m�����~z��wQ�+GTE*�d�^;,�z�qT�EL�#��+�i{���͡�c/Tٛ<~�)���d�n�h��["7����-����҆��K �z�1�`��&tK�F)����}��S��p�f�y܀�Yg���H�'ß�F�f�T�߁ys�\ɖ�5�����ܢ7l� �9_"�u��X��!^� �lՆ��M��g?@.����Kl���I� �y�m�����L�!¿��YGYY��%¬=�<�S�+�̜<����F63�X�^��u f�K��M%���v�/qeOF���)�'��FO3�{�OEƪ&�?.	�j&��~c�2�g�����SP�`qM��fn�T�t�����4K�7g���_�0��z�A$%ޑp��6�˼��XE*`��mLx�,�cra<=AsԚo?��,l����xV��=��%>2��ƣ��Ŝ�I��%��]��@Do�ȃ���Ub2�^�+���W7���z�0tj�M�6f(���䩻��S���͉-%1��#DJ��F�E�.��j���X�!�VW�r
[�껠�v�
��e�����!Qw��goCzW:a�ءHL1q�ٗ�ɛ}��x��2�ʌ���[��X�v�m͂��5�o+ZҮxf!#8饶���]����Ts�BE��B��k�X6o��[��H�f�tO.7|z𒢐�1K����C��~6�^1п����1�x!n��_ IH�+_1p0���؁�S�i�`N�뒌��eL 6��VN�)�WM@u`�
�s��i��g���s�W���B�䍎�+G �fI/�ځR����yȎ^�EGxc���cҪp�l���e7�0�ǂ��Z\b��[�O>���2�ƜS�)6�랊!���U]��$�4���>��36�?����K��,���DA�Lq�}�;@9{�B�+-e����C&�-���*
����=ܩY�6�X"�3"q��¨�Q	R����5'���E��)���Y|
Y���u��qx!/��. ��=N���6[���q�^g��j�G&Zxx�!�:�W�K�yr�cY�I�R����^�x߫�E�"O���y�q�Fڶ#�@�;�8=�%��7�����d�NO9.ӣ�"п拱�C��τ��M2�� X�QL��{ 2^��W�.}�-멂u��������j�[��ۇ��9ŉkFu��;��Ň>�e28�� �/ǔ�ĝ�?���@>�&j�EL�N�,�޳o��18�=y�* �5T$�26�7wH\mL#��M%n���<��
ÝV�ԃOq6������#��.`��9���\x��}>�-i�dͅJn�W��W�]/��jm�ik�h��j|O� f�Kޚ]4Ag������v�c=�0K�4,���gt�������S�����`�ՇX2��+�x����Qc���0��R�a:ow��- �jLF	�N"�W�IB�m8G�G���VbF锖S��esS��3��/Q�{��_��Y��'�������%�c[���H�@܇�K+z?Qx���s;��F.��ߏ8�ޓ�����T���=����Z�טU4}h��1(L������k�ut#��0[C����7�S(:<���4R�R��%�~C�IY�=Q�vWĩh:��1�Ҫ~�����I�v_o�k>��΢o5�Y5t��N��8ʱ�b�E1�G��=�xTaڋ�|���Ĭ>�x�����q�4�!<����%���I�\�b�8�e��l�1k��h̑РIBQ����>o%�s��)�G�G�hp��(ry�R��Ȳ)�}�.V0���n�pS~�&��F�^�1����.���6�_@Y�]�6!�}ߘ��*#)�y&��:���[�
�v׬�9[28�A�dD�QVh��-�Dǫ�W� ��뻽=�5��*f�#�����׻��,��].�8�9Fn0Pu��Vnv�\�3��L��G/�r
_�E�XO\m+�[IQi��~D�Q3��0Q�Wm�R���]6Ϡ��$�����?� v�u��n(�e%�,�X�	K������>����J9Rr�Wonh�������j���K�{���<"Zh�Jd�BBާ7��X{� �2C �)5�,��G�/2<K=.�=�,�?KQ��X~��]�!a?c}��-P�/����å<�������P��8�ut$��T�t�����a���j���5��4�E�i̝ȕşn*�0pkg�1�9���v��~@Q��t�
�v�@}{��>��|�^X����ZQi�c=�xW�=�W����`H�7�kpq�\�H4� ��-bK�)��lmbiY�*�6 ��ˬ-h{�G��UpڶZ�o�g�X�F���5�_��I���)"�S��C����E�D�y%p>�����2ʹ��Z�$*�g���s��KVU�3Ds����y]��rH�cl=\��3�K�K<�wK�i�Y�?-����3eE��s���D���M��ɹC��,?Z?tOns��c�#�Nģ��N�s^���Ŏ
CB�?J<���>BK�/_�� }�&��K`U���2&�w���|�ﴅj���;��#�\~ eM�R#Kv�� ���N}�{n�S�{?��)̪��8l,��xjy.�ŭ�>wE������Y�B�H$L%������]���,���w��<3jH���d���K���0�ʕ��>
��YdOq"so�ɑ����� ��h�D�1�joﺤ��y_�Nk�,Ԍ���s0������� �(�n�r502��t+�>-��*r�͵���������f|�J4��U	�k�����1���w�г]��o&�$���~^p�&�a 6��OI���GS��l
�̣���՚	t"-�����Hb2+����/B[�ápS#~�h�wh�g�	�;�ӵA[�ހ�x��ίu7hɥk�0�Kg�%�g��v�<s�ߦO�N��*u곝 ���R������j�0�ў7��1N|�
"|�Vk��@:E*.zh��l�9@ԌImc�Qx�Q#wTz�OR6����@aٯH�rF��a���4:���n��(�XJ�mɳ��E(۝Z�EP��N�)�?҉�m�G�����@�ͧ��
T}��.yC�N͘��7r|��vA;�,4��4Q��k���y���ȭ�>46�/�[xHd� �Z���ga��<U��v��T|�]�(T�^�����;T	���DfJZ�Ǌ��<6���m7(n�o��T�_݅�x6�c[s4��@��� ��e��	����?}{_�@0��޷�d�g���)>��<�y�2�u���Bv	/ l]J����6e7�E�ղ��������v��s������;D}�lEO�B*X��h� msBj|�~0q��A�|���}j���{A���϶�!���L�`�cqGP�ak�꫈}W��ì�3&�f� ��,�Y���*���Y�`⦶�̠������)Ii�k��s��G�L?D�o���q�l#����>U��CT�q5�#ad��ޛ,�n����Fe�Ak}�y.�<�|h����������Ǯ;����ȫ����] ��E�@�>��8FZ�{G�g1�B������;�����b�N�N������j���Jl"b�S��n���tl��֝K]����&U�X!ZO(Wg��$���A�����
ʜ�]��v��XdSMٛ��cG=��Y���yIA�����x�|p��S�j�K?��gJM,˦�^�.Z0��D,�
$t0�`�}��
�ͳ���yT��nLŔ� ڢ�4Zz�	KU�o��:�\�y���q������t;�wZA(����z�Ь�}�=�
���4�c�����ƫmR-{�%���دE�����QI�ekhT4Y!�ࢄ(���u��ı<���b��pZ�8��;bc��X���63l��3Ib�R� @�"ƈK�$�Uyߐx�[�pT*��Z��>��0�aQXX���Yl�Z���I��'�J+�Qk{�����j* ��S)�@�Q�A��.�1fp����tS��͊�\N%;�#�4>wW�/��%|2�]e��p�Vv�.rd~m��j���%=
��l�]\�I�=�OUh��t*�Cw/a}o��_�uR�
uC�$�-��xZ'�G�T��]nQoU�<`=�3z�)��7?�=X�a��u �����I\c�%�v�X*G�J���>6�-xٹ��9��^�|�������٩�>a������~�=͛��	���{�}a}�=4#��7��o�}��WX��9��t\øQ���рT~u哀J2��Oq����2�$f�ƴ]���܍S5E&Jg���
������䩅��) L����Šú*��'��w����C�iF��l/�b�"��*/e�i[Ա�*H��f�L�Oȗ_��Q9Z�ٙ-�� ��A0I�H��?6Ud��hT
B�k��A�?�s�-��˳�Kk��(�� R}Ѵ	xied@ذ��BJ�0![��NfT��������=M��u(���I�8�^��iU���|*���޶wP��^���z[O������,NS\�AgLBj�ˇb��_�ER�TrY���ɋ4!�aB��ϋ#E�� �Q��\.d�,�x���Z���۠N##�!|g����h��9&����l����Cm�~^n���r)Qb���4��f-��7	Q�v����
��tG�/���/����'�J)��㊊�϶�����]������c���U,MɎ��p�R���"�b\F���U/��&Q4�@�/���e��͏�M����T8�rp�f˴[M������M�v8���2��]B��;�s�zY�$�d�.�����c���{��m�Pp���Iŉ�{6�����!����XK���r�S����Z�^#��y�PN��%i��艎�Ѻ�6W�S�������/|B���͗��x��KW�W0�P5_�g�BJ��_1ŕ�5.�N�+Ϝ4ci��;?�p�5Rrb�f�Lҏ�v�bn�P�5�%-<\��)��P(x�1�{�������"DSW����m��:���w+���,𑊱��AT6"�0�_ʼ��׌�?���Pq��E��Za%6A�$���ȽeM�S|ŜA�?=�X�bf���p���>GG�)����g�a�XM&�n��m/��iQc?T���8���k[,�Mz��<�~����$�g�J���Dl'�.�q�`>M)ۤ����U�F�{�����w����^���eJ�|2�֯�i��Kb��<��b�dǇB�u
S�Z�쟏������� H�~�f�U����<�G�1�~M�i]�`��g�o3��,]~MK�ʫ\���&c��]��! %�A�F�<*ādMs>?J�x�3��cA�:le��L�%u���0����B8`T�b�&J�m ����S��TI~\2u�Oz�a�>�%w��R�b^ ���x(��k(�M�EGEXdI�"�ҁ+���Z���p	���9g��/���&�vޥʳ�����Wǆ�#z2���\�x�"��ܕ�3�E��E�W,XB�~�`L�*�7�ӑעAjY�<�����dy>�/H���Z	f���j�>�`ݦ�?�'�t��ԫ��k�}ڙW�T�YR����$��8� *y��=)�'��U��d=�;Qwz���/���f�nߗb�3�-*�ZnZL��0��x)�Aܖ�'Cf�	���U�oZU��E�S��0��$�u�����8���'.M���v/xv�-��]��K�2��NgQ��ee�����;މw�,�!s�[Dʁq�:��aVU��A7��j�d��S	jE�L>��*h�H�t���k��8�k�R7�v�Z/� �H��@���,z\Ah����I���6n������?V?4�r?�`�����cy���v�_���J�����	�3�	��WW1�o�H�/��L�˖82V�Q��}�GA@��b�LP�����aҫ���F�?�����W�F��ӆc�ЧS����WS��9Ѳ�>QQ�>��)�iw��A/1�l	�\�u��'5�-�ڣS�U`ݖ���T�q��>���kdK��Qvʮw��Qd����B��[D�Z#GDc�>��J#x\k�o3�-����f�Ï�0P-�e�o	:xy!c��z�����|�:�*4��B�w�~��Ԅ�M���sm���?��@�l ���N^�6dǇY�m{��1���i4��n�hKu�w���쓷��������y3���Z�<4�/��9Z ٛVTP�O����
GZ�]���I��HR75�"B8�y�}�k��s~���Ӹ�_�����c��\,!�e��9#��K��d\
�U�%��#|�w�G�n����'������+w�휦={���rc~9�t������7/=��G�?Y��WL�ni:��.��d1�\q �D�!Ѕ�6�e��� {r��3�:�#I='�x�ƭѩ�>�A�d�����܁�����6�8�̯,��@Z��(�䟴�T2\S����J�~P����6�3扨W#X3�����^`n{띗��ݠ\���&�^����A��Q�g�����]-в��)F���r��;�0�x)� ?�2߸-�����E1؈������>���F�bP������ä�wL��#�9�,��hJ�Cdz]85�(4՜_�!簘��a�+�	̓��m�=�^�|ըa��uO6�@Iݟ�=Oa�.i�i���h�H���\:���%~�;%�v��&��bK�mD���d%�m�5N�"9P���Ky" �����)d�ц/�U�-f�] ��:�R����) �Iew�l�(����\>���� 8�4���^ xr�3����[�����4�F�&�O~A#��N�#�91�E�!Z(�K[����E��4G��db�;!�5-���]k��F�Nw�X��R����M醵���@�4M+Y��[/p����Ʒw�^ػ�H U#lcL}������?�c=v�*��jҟJ�ҍD[E���bQ�gR�F3�"ʓ2�w���@��&�z�m�o�%7����eR_F���@�E�EĢ	�x����I�~mn���@�C������J�r-ǃȧ�V�l����A纑7���18bP�f,j���s��܄�T�Yg.����a��c��x��i���I�gg�슓��ũ��u�6�ND_��v����[���xL�� ���l���%�K���E=x�<����U�[M[&���䝦��T>B,m)�*������GV�vP�=��Fv����!����S �Yn�$�� �?Z��MښX|��6��{<)�m5��F�x7�3���~�>\�a�X%���
�����BY�x-��#�y���Y��I.���惨����Х�Jj����J:��|V�%�[�*�^������Q�6���I "�W[�Baw���� C�#��S��Qbin�G|�-�:��_*VY|����)ZhO�!$G�U�e7Ψm�S�m1�en�d��J�&�,�|a�xq�R�=�]�a �I���J<�+(Ut)��`��2����c�@<�e�ɨ��i������aXw�/+���8�5�g0 �:��0�l��br���~��ʖ?�B�z@���h�
xکr��L<"������9�o���!T�9HLۚ^U��-�"ݑi�o�-��CęF����W��V>[��r~���ydH���P�[!Rc[Q��M�ŧ�ɓe�*��Wd��HC�������!UmB�/fΝ}�����H~8�OR�=~qW����oP"G��t�h4�a)���t�wN����Վ�5��[�@%NݨO�XdƉ���y�vu�D��z[FoEC�9JR.d���
�!� �5@���\��t��|�j�,-L� h�Fu�.M|4bY�v�׈���Q;'� �m��)�?�0*�d��G���2�0��jdW7;�	U���������cJ��bY�d>�K@_����~X�<�0��R�1zu�/z9$����H��#~�|ʴ��L�{c�,�4h+i��yS̯L�vT��j?[	��:�M`�oK���#�;�圞�k�B�\�Voeq�J��5W�[��~����}��}U .����zRW�L�:�x��>�=e#����T��@&��6���%��}�;s���}׌e\�D�� Q^���1�w�u �*O�j��<�H���q��H<���������俍��]�*!��zw��vC���	ÛwY�ވ���Ω��w��vQ��W*�2��M�/)��X���2��]7�ԭצ"�`xv�\�����u�(�䏉B�����O�����J�ؤ���\a'}�q6�)�q�����ӵ+���S�u$s�sk��+�~����� c]���7��[��mί��\1����[x�Z�2�4�y��n#�?D�B���Ԛ��|�	��Z���t���{�Y�'n�����cAF�lr�wa=��V���G�`ׂ��-D�PY��fEK1Np�l<��#~X]t3h����m�^BG�{:�Q��@t���D�/�t���y(�Ӻ�X�K��,%m�s����Rx���#�j�~1<�2ڕ2<���m9�L��*t#2�j�T���P�@h��3O� ���Y�ޱ�g�h�kqe&G��q��J�E��YK�@%瘉�h�?�DD{�/8D�����P9������>M��4�M=�YjZ���y�uGew�p�ƣ�6n�����tsY�;�K(|��v�^��wB;
Ȼ�$ 3���;�b��.⏥t�E]oBu9�A�.���b��X����h��<��w�Fs��
M/�C~d� � ���'�Mu��NL(�k�I�W�(�[��U��\�r�^?w*�H!��9�Q��4	�J"�z^�YGm�.ݎA9�o��o�]Q�_��zԛMg���9P��Y�1����4N}��Qhm�����>=�W>
a�6�	�R�=��,�|Tj�C�QET#�q_ʚƉUE~=�XB(�X

E�"�Sn��0�qR��W��\CGQ��DJ͜��e��dܾ���'=��:i7��F�y러�s��m�d��һC�%ӴS��h.N �Jq�!�'�5��sp:��e5�X�?����<��:_dC��nL��%������
2�e|@��IL���Wq���*;�j#�cv�t��?�3яM���[��EZ0ev �z �� ��/��ԺK�Y�P&����%�:��}�M/zX� ���2J����U�aҙ:�:�(O�|ސv�SIī�x��;d�,�z7$�D��,�JT����VtUg�e�;��������n��=�7y�`���糧S��kI@���$
Ν�����$���t��C���������@P��*��o�o���P<ɂ�8�EIS�1�u����b6��/P�ڽ( 7}Q� �[u{�E4(�r�`_�_�����c=�x����p%��I��go7�6�>-X�O�J���`���ڨ���,�|�8�v��	8�m����(�>}ϳ=G6r��e��"���E��^�77����'[�>g@�A�E��{�D)�lZQ��Zzz�%�A�b ֯<�<"-�Y�֓���0��	�z��>>��<62��Y|�Q��hK�����,���?.ɘ�?Y�'�+��9V ��D�W�͍}��xS�^W� P_d��OsB��@���ߊ�Ad�߻�섒�`^�>��L^�y��A,�0�*XYb�����߹j��#gC��>융<��x2�����RFT���TQg��ǜ��B�zg���4�']��ƫR����r�ݚ���(�����w��\�J�Z���yQa�B����Z� Z���<ۏB2q0�E�h�ǧ�;d�_#�8�/�V�ha!� ��?��C�ڿ�m�F��_���w�2W��Gɢ��F����>¡#�U�Dx+�z7��:��Q&"��t,A�#?��Lc�@V���C�����ř%���?~~�$�r���0qV�~�3(`�2�\`s;�����D(�ayߒ�P�&��7��D�tB��#c]7�o�AR�K�x��?���ꃬ��M2t�s���g��CZ�W�܌�R��an�,uA���� [k��|:)+�v��j��p�l��2d���$䟨-n� [�:I#C�(�Al�QU�M��f���R��|=(K
_8!$�*yϖL���ɒ���0:@�p/��Pפ
����B���� �wI���oU���0�������FXr鯺���4�],��$x�tʊ����/z��
@A��r*f6J3_+O�U�eCX�"V��(v������
�=�H�8���
��>�wHUA�t�͙��VM>�?��T�1��T�Da�^�3��:����^��SI�f�NpOn��GS'N���G�{�D�bBO�T��:V����K*�s�f�L4OD�&W�'�kz�H���G���j�R���8q�O?s�5Pf']�>B)ffEH���h����A�^pT�4w.�3dg�����Fޮ������^�sc����A�Dj{�4v�����J�����H�`r57�)�	"�Vg��dgvC�D��1�d��!����vP���Z��Rt��-m����	�&�΂T�QO�bl�K,�|h��[4�a@ߵs�W=+R�%Hq�B��Jc�Uԙj|-��^^, �_ǝ��>J%0FBq����{.I��N��8�I�|��Җ����A4�z���Wx�Z�>A>�gT}c��.6�\�WRi�kg'QÒ�/�]�Z�i��U�����{֗�rRY�Hv��d`�4�Vԕ�_>捗�^=!?�(�6w�X���l�(���Ob�s�=
�;N�$� @��ia�ԅm�ph�`$�Z����r"ym���V�,�/�6`q��Q4k��K �a3Fsn�i8��
|=�E�֓G�-�0Q�r���w��Ko�^+�r�Z���^�
�*bH�7������+����g�W�<##�&�I��J��t|�U���@����zooľ#[��
�Hw\�i�:СA(�O ����h�׍�Pp�  �?T�O@�(Ͽώ�gcV�8`��c�c��#( ���x��eZ���ǚ�:{��b�s���x�JB������Z�m��Ꮮ�vjk^��`���)U3�8���mN�*4��,�����H�m-��cx/6�	�6@\墂5qrΧ��D���s��K;�ߦ���t����&9����]�N�N&9�������8X���F���o�@���| Z����@���3[�12+)���ɢW��gK��M�h4c$˄�xTVPv�ɔI|����L֟֬{^�Y�.��2��,�.)�W�/qx�?~���\�.���	i���g�U�Ľ�3@݌�2��?��k��Ҝ�!�T��U�v�j�-��|�n��Sw�ND`#�;b���4Γ���E�"���߫���袶�&�W�����H��ZHVoƠy��A��h�7�Y&�f��P��d;�m��+�kU�AZ`��I�5O�;N��ƻ��v������sz�D{s]���H��}��xkl�z���6���]��Hө=٨k�1�`��4m��'���(g�Q��8����"�s�k��vn:`�����y��:y��eP��l;��z��:(CƂ��:1���GD�&�c�*)�Y�c9�Lor�4:҃Z4�YP�Q��.nK]A��j���X���F����� ���Lx|M�?�^~g�Co�(s�wA�ə>%@/�� j���Xmj�`'���@P��G�9�dn���hI�4<�/���eED=Ͼ�*֭�e���x����?��*4_�@u6���%P��P}��Q�Б-����]�S�,d����:$�ª/vg�=$x9��A�_�c�b�{��c����燀e�ew�3���z�Rk��K��?ǫnW�I��ί���#_ԇ�
��ԢZ!��3���K�߿��SE�t�,~C��\W�ę�LV�VH<�F�6�Q�혥���4m�M�#�ߏ���4dEH\���4l��l ;v#��%����&� t���n}�eޯ�
i=���S/P������Ӽ��ζ��\�`�4��k�Ĉ�f���4쮠5�M6�JZ��s>��X��T0<J�j:ANa*bzݙ�<���ẀcRiI�L�2���Ҏ�Ѯ4(�yv�OJ�Jq3����� �(�S�a11@.����וX��7���F��=!�B�-zo�;�y����O�+�8F$y� �8{8������� ��g�<R�v��b��ˑ���n�i��tƹY��e���ǈ|���,�Y
��c_��dF}U�ل�5����t��v`��s��V���.�et��Ӡ���J^?����d�Щ�(g8�d������s����n�M�]�d���<(��b�=&�D��ޢs6:�KI���6�S�Hq6������ƥP�t��X�Vq&�)�a�ç`��c(�m��[x�����j�1����D�`X�7y*�uG�ݰ���ס�j�L[g)� H#��JN�=:��5� F��(7����� z��[�m��3�)� F� R���=���yfʶǃ�c���W�Wp�u���G0��CT2K��i���z�̵�҈}��������s���5(���q�ie��|Ӝ���-YM��7<�zj��.~�N�l r�Mn���fH_�#hK�����ٕ�9A!?���dxTM�x�|�|Hy�j��Ղ5 ��,�_X�����W�
��-� T�?:��6�+�(�J�����),q��s��I��]�F��YQZ�:����]g��a�yy�K�P��_�~&�Ҥ�;7���	⌛3��_���d"!A}w��{��<D��T��ԄF������e�������,�03����d����ҺP�9�%�d3fK���5���e� � ڄ���q%_CC!=X��	_<�mᏪn��Pk�M`c���)�Ky"�j�b%U��=d�
~}�&�c��| ��4AO�[ّԾ��np�[%AE<���}b[���f#�q�����5?[f�!���ɭ�,�m>�-J�����-\�}�D"ܦ����ig#%c~k��0;S�"3�w�I�b��ց�ȸ#��SBeO�\���ב�٬``��]tNwR�|^ipz����Α�'A���X�F�Z�l�)\A�=Zf%E�������M�I��A% 6�n�;�{W�1 *��j���ߺ7�4�w=?��j�g�Rn�=���	���!���2w����qr�o񷃀L�2�ַ���E�",�⧶�|de��hvO��j�A0 �7����t/��2`4O���\�!G�OLrD����s�fB^햽A� o�\�$_�k}@�PrE�[�����'�	`���O���0���0�.�Q�<z!{���@��_Ѹ�[%ø�ZI�P�U@W���D;���__�k�%YS��.��`�]����W�d8vPNW$r��RUY�$9�
DO6!��Xr���5oX$m����㎪�Ry��_�݁e�ɯ�k��z?��h���lgHP�l��n���vp"b�
��?zg=B0r]��q��J,��C?��Q�bZ��n|��q�)y��<߀M�߈dfB�
�8����.�� ��ê5ӹ	R8�?�����V�8�A0����j��c4�(m��ĵT��ɪ|��p&1|m�{�f#��q(�z(��/�9����T"J��f��o��P�:.��	�p܌M��/�w+5k {|�j��ֳ3cX/�7;�(���E�`���}�]�L~M��ݳS@0c��IL�e�X{o��T\��y(yn��=��'o&���8[%>�y�f��52��.vB���۬��xd��Ri�i�+��@4҂�UM0퀯xه^������ �Xq@i�-����	!	��?���!?s�����mF�Og6�8'�쎁�P|�Ή�(4�~o��F����χE&S�=�����Wz��(P`a�P��� `U\)��ꍗ��n Z���U�FY�Auw�s7ن��\hCTr1W����&Y�TW�#Ob�;w�'C�\�YN�8v�p��H��>9\�߭	�^�.�#�Q6ָd�`�|�̚������"�r�4H��,��RBM��(D�-A[��K��'��d5���M_pxS����oܧg�B�l�ze�'2���
)moЈ�]7'���,4�/2��b�����aA��Mo���!@���W)L�dW�9�}�]h"�1�v��j�k8�{G� ���Iw$�wCR�w)�]~o��v�\sk�
{':d7�e>k:���k��ۧ���ZB����V%*#�:a%�i/�ʾ~���8�R� @F:Q�}0���<%fG�U���Ƕ�}�v�~��s��f�
I�� ��2i���̼e4����ow�u�a����`� �>cp����|��AB���	I�hu`�7;�k=gռ7\�\��@�\�G��K6��c���8��?@^��/̧iʿ{�V
�o��b=�!����x��9������AE~��>�-�?x;�A����	]��^E�ƾ�N��˷r�@%��Pעٕ8۸����j=*.�S>@�mq�_S-B�^i��-_�A���g}S+
߷m\�vh�8��ҺG���^�\ �کB��M��Z��w������s�4ptԒ��Ͱ����9��������5�y�2\|'�F{K3��V���+#3��W�@7F�9�Ө��4
��e��5�Z��6�����B���Uք۶݂,-�g#c�ˉ�������.����?\p�5�r��X��3�I_�0���_�dO�ic]!Uo�pXz� Ow�r�i:%���WE�6C���~$���5s�Nr��W�',Y^$c�ύ��������TS��R<����~=~O�����H�A��fQ�*�趁��e=��d.�DN��%���M,����E&��F���Z���as��[AnC��%|Z�^�t�,�24.~����ArF�;�$�^7t�wKC�tV7OŜ�L+�*Ko�)��q��>�JW��#F:|A�a���e+SN�u�N�ZLU���w�r��C"K���w�9C����ByZd��r2*=w,o7^���K'������Y&C��������4�U͛y�;��:����_a��<��l��9�b"��3�q5CB��'5�wL�Z ,v��ve� �$�!bp!�uJ�ã$z�
v<�oz��@��Hy��#�6d�N�v����b�W7�Οz��	�Xpm�:o��搯o��˝�ikK|â��Z��'���#���1�H:f�p��Vјd���Od�]��C{����e�`�����ڿ5��OݸR��ca��$�hGNq�<��們��D��\���}im*!c�!�Z�&=T�tҾ���P6����/��ª��ڱ�<�O��Sx��v���6�~+��:�#�%�&�8�T��_7��.�eB{�7B'�n������(�l�^�Tx��{��.��K�6�;����j���e�9S��mm��cDm��'���?��V���A�Ľ��59���8��N�1��TBȾ��6#ڻ�K ����k��������Д-�a��T�&�͚��8u�8�]���WO�1���h�Ji�6ֺX�[1SIOE;{� ���x�;#��Zqem�B��8���K<_t�y*�~j���g�r�QA��\SI�5v>����O��+���%)	
����J,��1f<Sc��Y��1��V"v:[b��ϳ�9�J���CŨ�@�ºJ����܎D�E-��D[s�ZM"����-}VV�s�:�I3-T�'�W�0���x��Jc����z�'$��%�b֎�a	�:����W���J�"0���6\~��]�p��X�[��/A�\=3o<q�����i�(mO�fo�A���}h��<�*d��/�]�-�Ǭw�/W''� g�-�P�DRu�p�CƣF	e$@I|9�b�_6	���"^�SS�:Q��ںX��䌿Z��1�ʜ���_�C�ml�����ׅ���&۰)c+��=�e�an��Ś�>�Gq�.���H��f��
����Fx!�v5����\��"&�P딶� �\�O�5þBGF�$��d P�B�D��1��epG����b[,@�8r����� �	�o�cv.�W{��d	fy�K���S���A82��ٳ,nNY���+��$\�8#�t�'�a��y1Y)�=5_	*j��
��o���54K_SJ���˞�&H{��ø�U�l���R%y�RD�:8�3��@	��Nu;:�;�mj�ޠ��p���S3�?��3Ec�1� �:�	<�;�zH��Յ�u˯�:�=�A��Z�W�l�2Yr832�b�����?�#ӍM]�L���,�Ԕ����#��P�L�F��w�|��*�6r�H>��:סc������;�ZZXOdd�����OjZ��ٜ�u�t��`��^ry^t$bQ�t�5֜Ӑx����xtZh ��ES��S/��	UbSq0� !��/v��	�Պ�����7W�qTk7�0�t!, �n1 �m�3!�X���
:��������#]$�"�E{#��ـ�)��<�M���	��������V��4��'��}6��~ �`n�݊34��0f����H =�8t�u1�Rs	A6�:��~�l�����k�Kv@:�e<�ap�����7\�TG�C���iy�������男1r'�@���a�9�x\E;r�����d�_+��sx�iL3�H�!����Q�n�"��v�u�	���>_� �oYF0ah�ݦ����2l*΄`�a�����J眜H<�X������Pq��y��G48���5 9&!��+u�os_�:�]e��3$!w�"��r�,�p�x=[#����n��JĚ*�; ŐWp�IĻ��!��7��S�|h�Z����b!-j;�b��a_m*c��m%����S�ggc����h]�>R��*�z�C=F����?��0E�CT���A�����{��#|�/��佀��*��:�\.��y���m}�y��a?�ٖ:��e�e����VF�S�2�/�L�~[di�0�t��r 3��/��9�q�c*�x����90��j�31��\Y�{�-��놓4".@K�̥�?vaw�0��9������8*0�����QAp�4_�BKD���0���=�V����ڛLA�G��T-Dަ]uﲅ'`�&Z$��R���C��A��N�*�u�f�i�	�]�T2v�K��Ѹ2]��!RP�&��9�!�T9�a:9�YcN��C�k��ax������IQS����`{@a��C�`{�[r�''�Ef�!��/�8L
��s��٘����b{]��� L��������
���"{�ZN�S�ۯ��(m#��M�F�h<�y�KR������u�kl�
Y���R�\ҕZ�nnO��<[!�PO1(���8㮫nZ6�]��
��,�aH���h����]=����Y�T�ж�8�C�{�@Y�l�H��D�F����׳�h,�����u����T�\��r|r%���K��_�}�VB��f���78��:6۲�H�G�ٶ֤J"�3g{9w�������b��$FU�I~U2̟�a;SY�8D�Y�1%� ۙ|jos��.
�w9)��S9��nM�W�s���]�X�߇��k�˘�
�ޢ�g�����y$`H���M�m 7bR�Ơ�'��i=��:��ׅ�F�t��&�����lZ�a������G�Ua�C��OS4D;a)MXʗ:�q	�]Y�[ �*Ȑ�Ș��r�'���Ĭ��(e?�6��?K'Q���o��j"?O��K6_-���;�lh����?~��|im�5�3�����
�B�<�i�RV��o��v.F��}ȉ�go��p���[�����qL���Z$����6�|m�jM�Hj����O����=�3^��:̶q����p�����ty�;�{ ����fiF�|��+�.̀����\��	9�T��{pHQFf�4�J��uM�i��z�~z�����d�Hp͒�1$ƈ�]Q��{�Y"_�{j������;ܷ�(��έ�@��j.����l�?��/���t�sՉ����g[�����g����e�9>[�T�x�:k�@�*�Pő����_	��i|�/Dh�Q�LzG|�"��gu��+%/ȴ~T��Y1���b"1�0VJ�'8��cT�O����9�l*L��I^�ϊ{�����	�@x��$ɋCǡkK�cDg������Y<�!�HӬD0���'�O�����B����R$u���O)�Y�U��%������*���ȟ�j6�	Fd��mE��}Ž� ƛRO���C���t) b�|�0،�=Κ��x��<&2P�Ŷrck�f�bW���?l�4DŤ�e�']�Ly,g�$����K�ENP��KP����؏�Z�H�H��oa]�����	�V����Y�ie������v؆;�p�/�X��.���Zs�
��]��nHH���-c��ݥhs%�P�ܠ@˶�x�@T����<r��OsٓF�#�׌�o����)�>��;����5����2��Z����ʁ1������ Qⵤ�KONx,�C� J��)�v��?!Yg���RN��}#_�H#`?�z5DC�����x���8k<�+�ƨ~���=����γ�0���X��y��!%*�HH�F�~:Pd�>�������cAŀU���7 �+�F�ө19W�8���.j����F��q�5у���$�N¶C=�FM�F	���/6��ҳ�eU�����U�>�xl_��3i��S��b���<ŗ6G̍���M�	�|0�^B��䎳�=bV�胀�g��ƬD�bq3�=��/�/����]τ�;�$�L*�d�����C;*�t1j$p'�� 8����Ё($��ߜ��J����nGV��n{��aˋ�r]�d�X|6y����E#d�햆���M�3s`��:ľ[;@�~�m@���#��*Bk�����)���vK�h�;W��^b��g�-����~�,V�T�i�*�U�(	7�T
`s_�����j'�7[n�&j{)�g��b"�i7�6�P�k�� 
������
/dF��In1fOu�k��JY_bOW�V��3��21�� ~���v��>ч�-]u%���Y����=·��)�¼�ь\j�M������"�J���1��%o"���g���?u��^���z�ٹ0����A��G����ϖI����X�����IU-�煮���/)M�t�D�HK��墒�1/�U�odg�ٯ��M[U��!\��pu�
����!��t;-��0�e0��LT�ȺϦ�7%E)��cj�!�}��U�%�ŀrk����X|�G��({ߘH�7g���QDdzM�2���������^t���ȁ��5�n���!r�4d��\������J�}q)���C$`@�.\=`�3Vy������Ѹ�)����E"g�+5IGN��c��zҷl��`�+r�Cz��5M�R=e�=�aY1���|�sF���)��<h�5���'�[�`��CS)������%_�3�v���iZ�5Z�W-涒f��%j+x�����Zu���Hh��)+2m!�N3�q-��Y��*o��:ߑ�b{a��*�`�"�W���E�����HeJ�	�i���}��Я��OC߿��h�o��H���Ƀ)!o��[[r۰\�Y6u��cӾC0ޢ���ꦻ?s(�e={�����͘����/�ٱ$�c}�ݭP�H�)��_���;�)"d��di�t�d���:c�l!��:IUw-5e��p>�*�����[P,�!^�5uZf�H2�)����J|��b~b��[��^��-�������P?D1�@W�+t�z�V!�}��G<�- zy:عw�MS�Ꞥmh��6��h[7�ޖ(O<�T���{���j�@��4��1mc~XO�|Rx]�]<&�:�;�yv�oٽe?Άn���Q���3��l{��"M����p��7�P�-�̎k�W��7����q�N=��^ߪ���*�l���)��E���l�njkH�V�6����H�L���� �VY���C���N��S_�6�Ֆ���C���v�ǫ�{)��b���|���	B��G2P#�W�h��-L�Qt-���bUc�~2��H��T�s����Z���Y7޲��@,�1(����o�=�%N$
";�N��j�]+�k@z�e�� ���8t�YɶgV o�aS�w%�[H������.��
���- X��'� h�Ή�Xx��N�eg��\̼��2h��vg%�����V9�O{k�	� bن'A���5�i�[���1Ғ���F��� ��w���On�6m4ϱ����h48��_��� 9��m甽�>�g�~���Vn�6�,�*%�*/��x���k�V+�Y���t��|��R	) �e`A���y���(C�i$$,nlz͐b�(D4�M�]	Mﶱ	��o:�ч9$�?t�8�6�y�z�-�	JZ��:���F��D��ã[� }��P`�%�b��g�V,�J]*_Aܿ��"{9:%�����#�{`A���ϸ����j�A�sx�5Ϝ� *�̾ya��Ani
`�W���9ي
ֈ��UlH�E��D�MP
lA�2�'�Hw�+���i�RB������ڻ@��#o_�� /��/�I_(׆$��(����/'��A%5B�rT?�\ӖQzt3U�-�K:�"�x`"�ػ��
�8(�Y�ɿ=}��h%����m����U����ܑ@2��S�@Y��ߩi��Ք���;_�E4���\��+��=���k?_�
>٪"KdX� L�By,��/����!�!J|oN�Ӎ ��(���JJ3����LȻ��F ��v��C�"dڝ�֩���y��.b#�A/��l���j>�#h}�r�T����������c�O�pͤ���!�<e�D�nD�mB��J�f�.˓���UՍ���9�j)P�C|���C� ��k�3�!P�}��1�B�`_�����l�U~;(^B:XɣkH�c8��pY�������o*��q���O_wz�!�˛��әm6����%zc�O*[�E�V+�A137�i$%�,1# �Oу�+3�ٗf�����U�f+��&�n�O'��;���.�������C�;S�^��d} a��P|3;z��wӴ	v�R�x!)-�X��a:��x���7��
�[�3Ee(���A��J!�d5����᥾��W&y�g���~RD�S�d��̑>=��A
��v�Z�r�-�-��ű�5�2܋��~�&�ÝPQr���� (`Ȓ87Ϫ��C�I'
��V�o�	����~((%ő�b�إ��O�����c3�-����B�%Lqg�al��޵Z2�u�~��α�¹�.F��~�oe���WR^���X.��.�	u�)�)X��	��zx_�	�uQ��C���0���(R�X�.[��.����D�����НX1�t��Ӽ�2��P����X����}���J%<�S�����ٞr�o-.��ؑ�gFxn���y7����WM���-���Y)#s}��RL>�G�5�^��1���UI`<��|���D�Y��O�Y����=%�X[��7�d��掠�0.\Q�KqXh�*բw�����9�k�7;h�P��[��Lm�;oO�4�u6��DXr����r4��ψ��l	�8���rk������C���AD/���g�&�P��mmǕ�k���|mú�E��nk�/�& ���E��~�~��9�����3��&���*�l�clU�
(cӊ��~|�k�����d�X�F,�2,cJr�A��}�21=�$Uݠ�67+���������ɴ�����_�9^�xۼ
��%w��Qwck��fh��}���-}�3�[��Yb��$0�j��K��=�	�D��;�Ѭ{e�Y��)7��6~�����a�/6�������\����:8����0�[x��4�H��Jl��]���S4a(�t���>�0�Hg�� �l����r������;�1�+_H�L��=4��eaL��|��ʷL]����KR��9���4�銇������`��[Ktzs�bN5+Kj7�P�}�}:g�=�DG�*�Q�o/-����z�Qb�F�*�h�QOБ���b���D����a��\M�(�9�0�+:N�f(Y����.���&r���"&�V�t4��$W �j"�:�1Ķ�9N*�H���)S�Ռ9^�[ǵ��#���A {���Bgh����D ��Yr%��ƃJ2�z�}�p��3�&�X�f��@�N�μ�ö�{�ߌ߁��&$�u�O��4&Կ1��q��e-|�/��<�Q_��x֜"@w\9&��i�b-}�@h�E�ds�ӆ�y�Ꝋ໢�%�f)E�r��xR�a=��8C��!���wjR��t��㢭��?M���N�LB�Xa��j�s�ywjL�V+K~ʆF����v�]�C�G/C���� +I��	�ľ��i�t�O���iZ�~�@��$��ʦ	�V�=�<9mr��彀5w*�̨1���m�/'j8qj�H#�[��n��u�ER+�pj��˃`?�������O��T4��8�X}q���`�j�M�'��4*�a��Mb���}{0�Fk�`D��4�@�Z��f��U�8�p5��ɺ�6�}ǵZ�����!�*ɣH����Sd�Jҭ��	t�	�֡zF��=cU]z<!�{�r������a(nt���.�2���$}�������NB�;@b[#	mx+W&��!�.�v�1r��4<�o�{�����!�S�jܑ�J��ģ�?>�#,N�l7���`���F�t<@+�2E��gw�Cbo"6�b�;� u��̃�{���ː������������;.#���_��,3�ԁ���L$��������]���0�9�4���<94���{7a[^~���M�҉n�=n�~�q�4�����Nj��M��X"T",��<�"�h���>����>H�"�M�XS? :�D;�_S*P
��7�-Ĭ�K��E�3��V�":���4�\2�a�'�"�%"����؃�!i��#�`�RK��d�)2>#R'5y���
�1x����O�#v�7dK��h&��oV�)�'�;p�3�(*���ZN,Z;F��7�S�@�A�ۮ�l��޶o��&��2�i*�9|�'��C7�`_���������;���P��1��u������T侠��V�`��6���W��Kא$����Ls�1�F
�'� �qu�u��L:[�Z�ܮ��.�c�G*��	�Z��D�����$ ���>j|)��&~�+��f�H`�e����uw	��܂�ٙ��0�Jg�/j����.#֖ג�r�I8�?@�`X%P������G�8���7�����@���@x��\A����<��&�:2�le/�I̢	<��Pҭ!��g�͹�H=�1����=6�83�\�s_�[�Y�DA��jkC����P���r�^�l���/�dKWF�~f�r�&�B�h��)��4~],�m�C"�a�]�7D���� E�٠UI3�{�P9#U��y����E��fkj�-�_��� C�����;4���ԇ̣���s9��H�,KpU� ��A�L{��+�zW_�3w��2M+����\˾;5��tA7g/]����W%*�g�8^ev�]��pa���pRk,�0'�%hW�ժ|���e|Ɩ��;@K��V�X ћ�$�+v_ŗ`7>��"�q�SΖ��T��"��x�u'�+��3�=��``w����Q�sĒٰ1z0�Fv�	>�$�_x����m_� ��e��8��M�	E����'~��
Q�E��WB@$p���ە�@�R�gkbJ����4Yȅ{�J�ڷ2��.� ��u�D.wGubcU�`���P~w���W"���kIp����3�{���aa��NB�9��7�>lg/I��A?�7[�S3����χl_�i~V��d[��п�riٮ�r�Txڞ��ŵI{���;�ۡ�~>燿��u��/���MK�S�({�T����mI�0�
��UqTN6�{c�܀��.�}�ӫP���Z�q��#v+'z�V���~ã�O"����5�n4�AA����l|�ق��s����0@u"G��w:_����**��izu%7.�c��#�`ZhKw���9��j/�x�r ��P�t��>�#>z�;�j�K�%�ï��{�`ѯ��OUqo��oO�[C�����@',XJ�y�ЄE��"k�8<A4|��i_$�z1��і���9���a��RYu�Ӛ�>��~h��U<���h�Q����;�g�ކZÅ4�i���<��y��=N�L�#4w�_a��y��$o%�ukɮ	��m�Ss�JI_T�?�4�b����[������������[C�}^�Y�b���PL���7����+�+�\j����G���QhE�2=`�)6-�V"o�\~���
,m=:CL��WH���[�a���-s�@�|�0�׆sA��u)�����G3="z�L���i.����Ы�_U�+n��3��
�s�=^
I�d�R��g�.�u��%��l~�&Mrz��]��Eh�ꈍ/Ȑna[��(��N��^��TqLN
��R���I�R��C�@z�IL2�VXF{����)�Z�����:#�\�H�c� ���9aES�!���	<Q���&x���	:h�t\��C�V�l9F!n��T��<;�0[��k�7s�����O������'N��"b+&� '�;�y������)�#���)��
��ˎX^�o�K�#ӎ�^�|C<l���m7A5Qс���^v,6a���Œ"���=�)#̕q�n�<y\�)V�zM��f��\<��Qf{��/?����E�JX����hO�ًn'r�C�� ����5)��90I�F��W8(@ʮ�{�����)ʮ��" DU���o�_	'
�~�%�U؋�V�Bn���(͑<�v;�~�����6���(��: ��=|a&��4#�#��ny���U@��kB��)g?�J�ea_uo��`� �7���I��&��a��~�$��a׎G�W���D�r`���#8l0��ތ��s�"�Є�4U��I�ܰfL���*Ԥ�j��dH�1[t��Ɣ*����]��%�����f����D��S�5�!n��|����TRh���\����}N8+����������WE��#ۮ>��2�9�B]`��i�I��2�j�ۦ��{f������33Z���� (�O��sU#Y��N뮕�z����'F�@���E��8�\�H�A���?U*to;�q�����B��Y�e�MC�מ:��J���UVx`ꗕ��5� D�`��eչt\'W��Z�M۱���FMq����s��T0A]�}g̀�E3��'�7a��ΉFKh8پ?z^��JzmDu��@ѱVՐ�⾒I,���*�������I����2�㝑���À8� ���T�b.�݊�N�C`4��}{8�;���������T�b���R�Q�v֦�e���O�$sj�V����2�_��XE,�Vo2���mXrVpv�l9!�ހOT�D5�L�̧y�t���DHoĜ��
cU|`#�8�R
"Ee�v/_;� F�? 1O�}�o��67%���q�Z��|���Ζ��	��`ٕP<-��(Y�9��	0*�r/hV�׸/^2N�?|�LY���7�6����}����s���!fD����0�:�:�=*)D53�X�Ԟ�4��{n��Rh���r炼-�H(VX�݆�y	MM�H@a.9��Cd�S�m�A.ɥS��k`t�<L- _O����e��	7��ۨe��/��|�p��m*YH���ˎH�[�����iVw���KiM�UΓ�P^�熷��n�{+�`0�iBD6~�Yr��_r�	��N���ai��Ý��x�Uc�� 窪bX�J� F�\C���{ǧ|�ÜO��m��X/�+�o���,�߁���s��N�n�:��Yl� ���ҷ��Kό��pzi��E3�
�Ra��Jng4����E�`�_�]����ڂ��:#�^�$�ͪ�$P�蒬��zx��l��X`��ߧQ���կ!�OfO�>��!��=�1{I��3����8�r���B���Lyn�Y,�#dc���	`�g���%*�kB��Ⱦ��R�?�q�6�b���
[������Q�;�7M���G�����]cO�1�w�a�כ�����q� �dx�"�;S� ;Tklj��0���;�+��I�6Ii��#���Կ�v�}�H��~^6�YR�,�꟟g����ҋ܈���G��]JsnGu�)V}VJ�Y��f���f��Z/{*�b4�,�����\0Hˡ��Qw��G7R	�H�u1�٬^)��;C�ӓ[
���o2̿}�$Zfi����q�<�#bZ���~�%V�@L�Gi���t����mf����l�(H2^Nr��q޵e�5^�5��cI�b�R��ÁcW�T��E��ԭ�D�^�j�v|�H�D���nJR�A�Z^��%X!x��b}�o'+��*�;[cl)�D/22��\����?s�e^�nq�c�iJE���Bw�35͸�ݰ�B�i9^�:�P�+���w�Gh�_�Vmd��ex���Ƃ�ҍ��Gl�x",���g^Vܣx�ټ�aR6�<���iNr�Q[ q	��q���d��DK�z�u���@9��i����-Z���1ꫩ�|�Y0��]�7\��0s�i�� W�����(>��?��i�<�Y�K�j�ubV�d6�]=3�ی���ԓX�g��`<�a}){��1��g�2�4��N��Q�p�l1N_���'m�4mŌ~���Ng�P�d�#ۥi�p�vU���.\%JX׵f�����h������[	�7�/�߲���UY����X Z����kL�:	ZXx
�m���_k�c1�?(i73+�>'���Q�5���ݿ뎑� 킠�Un:틍�Rx��Ë0��`"�|T��	,�'�jB�����;�����L����jDt�ޝ�%5;��?�ܯOv���5A�Q\Џ�݆Ԏ���F`T�N>^cB=:jv-E���FjY4y���8��V��,!'�$/�́���&��MMW��\4=@�a��L�D/�O�r��ʱ��P�^Ͻ0'�
1��b���usS�2�P�q�tҰ_�9��ϰ�����)�H2YCL�uфpT�����c�#��>C�z$Ȥ(ڶ\�8nn�
3G!�����/��%V��i�~d��sX�y[D:������)�l�Pz�\�T	�:I�S&���S� ������uk�/�Z��g����(��u΃�T�Y���,��X��Z��μ���� ���ԉnuɓ	uˋ{����:�xe�{E�=q�d�su��޳��΄�{ڭ|���-�/�W._�M8�x0J�;�P��s��xrH*�����jh��H��D��Y#(e^�2.����d��TD��$����.#�ɚI~w�n��=2� J�$S�X!jIx�������oHD���4�-��}��e��j�+~�jV��HeiW��'yʍ�h�EX7h%3�DN�+%����ߓ��uo�2�zht���T����W'�C��t�]��4%Ơ���$�����Tوo�{8�)Y;�k5��e�a���Z�;���_7��~�Xz��W|V�lXT�%k{2PD�%��}B��o�6�i鑫!�+�\�`XmP��K�U#;Z8L��=ZY�T���POE��mxk��G.�Ջ���'B�J���*�n#A�
�]�Q��y> hz��5ϯ��e"^���aC�	��c�h@=�{~Ё>)m�Y_�v
}����7"D+��@ ���WK/$��&ݏ�314�	�eI(kq�+����#c����@P�@F�ȿ4 �k�	ϑ8'��7�4����b,|�F�X��	\	�� IS�ຒ8�5�Or�/�y���nM�>����|h��IIg똴�FJ�7,���}Y�]���2?3
����v�a=�ur��\��4J�ꗈ���vhY���*mV��1v[��?�ܵ�u�f��AaTB��`&Xp�F�F	�����1/'i�cHv����] �p����[�����M��#�Z�܎F����5ɷ!O_���=L��\5�PSfd���2Tsk����2����Eo {�ì]M�5)�1�+�Ǡ;LNQ�U����p�j�T�)�^�	��=�p�:����Bb��:�hKk�vB�7_a+�l���,��o2o
�'Ł>���y��%��x���Ô�͚X�#\�	��N����fV�=}L��������褋���`x��y��>���/Q��A�O��A�%��O�!���������L�E�G��Ӈ��6G��]uW67G���'&�V����3��<���+du4����5�-�S��͢뉁�ђ�ʼ�,Y�XA��g�{J�4w�
���&��BzS+� �`4i�׾��s^Σ��p$IL3r�Yn�U��D�ڨ{�ςx���;�u��|�r�z���2>�|]Im�H8~5>�]r���d��̜�-�
�K�e�ETXx����Q	�
<[wq��L`D�a�;��쨇�.?ߛ�j��>�PzTC/���9Y��e�v�[�2��Xqͫjlm�&$,v=����~�h������kܛ��~���8�C��iL�UEwLʭ�.+�u�����N�N�x�qk�<ȝ�4i�
������i� ��$�0���uR��An�aa�p������;��0a��#.�<TA��r�D�ƒ�9@�Y������h�J/�V�s���s)蘟��vzFEX�=([�D���n���)���Ċ~P��Z��r���P',��=^��-[ҷD.<hz��AH�g,a���/�^�靍��fp��*8;��ac)� �t`;�鍃���������t, F�zW��|���m�c��j=V|kƥH1�W�r����*�쏨�$-=ᢁ�mF����,�~8�GkPԉ�I�r
HGh�_��P L��J�^�*�W�zOMd"_z%������n$As2�k�т.�_W����	-r��6��C�l�7ff�=.Q �������|�Te���(���|ʟIȓ� �U���yb	������Y2�k�Gk��:O��o[B=x :��k�щ����N�|�}�	�&d�6�L~�%��,�����(OA]�]ڂ���19�1��{���>�#`e�����K{ߛ�'$&�S��-�Gs��@�x$���,�$k�,eEk��Uą�7q�ܷ��ľLâ�`&J�g_���	jδ����*�������;g�P����(��%����R�чePQ�� �O5�2�x�_�9F@.?Y�V�l�R|��3�M\B�s]/9���Q���㑕���r��������J_̽&���D��Ѽ��U@�ڌ&5�B�~�r9�wsNn����,M {N\��m[*���T�����PF��G-b?¢�<`����2���f��l�7D�C{�Iʼ��T����3��~�lt�>m�?��Z����?�+=�����=^QʓS�lۙ�Y�a�~�Nq8/�.�D�L����,�*���Dgr��S�s�Rtۯ���5(`Gg�F0U�:-���
41��ㄕs�z�ej�*�}�0�-���JS��6���4_
5�FPc!.������v�ӛPz
S����B ��o%�T$�7*��U �ږ�9���N�2�?����|��h�@A�W�pF�D�(8���c�����n4���@i6�OI���ɳ��ޮ������S�+�b{^9$f��/ZH�E��{����4$�CRc/$���~������ʳ��!d3;R{��wk��U+'Ǖ��<�i��d���-Ym�IuE�g1��G� ��DQ�O�VM��Ql|>��]�m~^��g��S�� '�.B��&?cBo4���� "6N���"�IeAh�DEu2=F7��M����/6뷦"/sq-�s�K:☕��ڴ�/�h�~���1.��?d�wV�ꩢ�㨻tl7 ��dщ#_�pQ�ᰏތ�8�*"mD`K3��E�K\�;P�QpZ�)kK��D�;�tv�3�׵�M��x�`�ՠ��ؚ.�V\lTw�q�`���LX���P{_F�H!/kHǐ�2�.�f.��w
��9B'�ں'��M�4�n�@B���Y��y?P�!mJ'"eifΝߎ-��P�Z�d�'��f-m2U��2�I����&�%��;Xcn�b�X�e/�<<�Vd]S�O�3� �w�k|<�Vz-p�ʾϨ=rzk��C���!�c�ܣ�~W��y��ˁ�&��Z��2���O�i�������D��9���������0hm'R+�ǰ\2��^�.uo�-��ZQS-1AAp���I]緃�2:Z���!�G��
��	T�.:m ���9�N��	8/@r#��R��æ"P��ճ�*yf2��M�ԓ�x[������{OӾ��V�	�q��S��:�&�k��'�?��&�[i�&�ۣQ��10V�I(��
�9�z�!�I���'��(��H���]Nt����B2�d ����F���kn��\�`#Y�!,���o�b��/�����Ӽ�ʃL���-����[:P=��W�/.�E����Vu߄x�w|"����~�brN��`ĭ�PR�&�&���"?�rR���P���p����6sA�����ne(��d�߀�O�?�7�1����λO��_��b�~W�b8\����P�kx�.��W�Ѩ�n핳ӗʢ�C׌{���4 	 ��i�0�j�i�y5 /���`<,�܉���|�M>��V�-Z�S��1�7����`߇Qu��C�G�,-��}�f�텠����P�ȅ�5������K0�g���_S �j�];���߀��D�w��o˲8"�ّd@�?�ΰ��V��>��X���R]��O7�v�q1�N%[�O�j:��ʗ��!�N<���"�Ô܁�b�x&�9��S P���;j�r�����A�Ug��NA�G�;T�c�!Am�_�.E���������� ����E/��;��u���~9�GeI5b�x4s��Z�4"u�@���oט�����/���'�"���z	3��^�M�(ǻR��R%�	���|soy����N�����v������;.>��΋>'���WcM�z�e�����ޜ<vŅ�˦�i�Oυy������f�
���qW*C��CR6�x��]U:k�ք96����~U��~��� AO��n݌-5Ď���>�WP�!����;���W��ܨ,��8�Ǖ�m[է�K��;��J�NL�j���[v�b��=���kB�J.�{�(�qْ�����j���U�a�{���Us`k���i!BE�-�~�we��15��$�$�1��(�h����Q�K��i�X��QJ����L	��I� =���������w������Q�V%[��β��%��#_=W<hQ�[-�� ��
��q}`�j�A�L��Q�s@,N	~�{V��� Tį���$8H��\��*�G�����j¯�ñYu4.�AE�B�1Cw?˧�p��y��'�ow��\I 	����e�R�O��j�:L�a.E�ܦ(i�\tʁ��O��G��Gq[o2o�ȉ~�R��R �[�\W��ǋ쯬Hy��6n���B�h�Q�u�Q(!;���<����8z��X��A܋���  �ʢ�E���mƠQ���_��?z��m�)Ka�f�
��@zn��K"3����}��~�)QX�V�Xk�C>�5\��{=�&R*�E�ϴ.��Ai�9q"��.�C�WD9�K�w3��r�9����:d���hZǉO����B�hR׫�%����h�\��;�C��K��C�&��v�|V-�S�W�g���'�BN������6����G����S�+>��[�޵��y?�$�y3�no��4����Y�C��]�N*�	��?����F]W^����^H-���M�$�$q�$�
�̺�3�����_=:-���c��`��Ɲ��~�9'��16dV���A��Ζ�.�}/1��c�����7bA�.8d�����4ڦ -���;�R��K���&�Y�L�]/��{��ctu�¬�?콂_��̑���Q���x�UI����$1`�,G �M4}o��t�Givz��)��A+�X�2xÓXĉB��(����u�t������������NջS�e���\��nP�#���	d&-��R�gM��_Z,ٰ����L�8�$��~:Ż��U;ր�ۊ��V싔N��ɽ��;򹞲c}Ʈ���޷IǊ���G�3����\<��B��X����L�%��ݝ׏�d/�Ԯ$��,�L3��E��B4�av��c2�l�a`��'����{�BOPb�uB�9l�)߫�c��_����rR5��h�������;f��L��|�>Q6�3W�Ǫ{�ky=�t����B^��L#.�hcQ:l'�V�x�i��u5����i�ag�-5��ۍ�ǵP��n�"R�� ��n8��q��/q�G֎���` �BNA�����EE��sZ-&N"��(�m��f��D��BN��1T�O��iv"�|��/hz/E��ҏ�%e�w��i�^�Hg�U_��p�{����Kbo��&(䜗?���<�6�"�~#�s�է.�ۮK�4D�Q�[��d��Df���xHc�C�/9航�Q�l��)�y��ݐ��ݔZK��]|�B��c�h�j�S)Ƭ��#8"��֪�?0Jh-�{�$�3��\,D�wvW�����nH�@ǿ�+�}��SE�v7����H&�ן��teJ���p���͸h!)�^����*���wQ���?�e�p)0WTk6a�4�&�~���{YΫN�x���*b��u����Z�-��:/ͧh3�1�9��v#0�o�?�B�h`�^�M��dr�\�$��5���5u���f9��G|QV@����H�%�|�_۽$�1>���u��M�{�5:�2�)P��y�U�}9h��]>x/����)�#q\�!y�/�p|@#R��ݑz7I���O ���c@.�����4\��>��RJ��އsՉk��@.bV|��a*ZY�1j����ZGX���;f3� h ���u��"�l���f��:��'m�J`��#��RD2���
d�t�|2�M͉Xp���g�:�Bɫ<��Pl�G��HcU�� ��K3��ٞ=�.S?]X��[^�4ϧ�lN!�w0���֠��!�bh���$ehߢQ`e^�X�~oT�o��P��IO'o6Q�#R��Ճ"���a��ׄ/y�>�'��E�Y�t,�(�FDK߃�Ƅv��QJNw}��."���M�Y�W�y|Ob4t������;e]�dS��,�ʔ����%�������DGw��ӆ5�$l5i;ْ	34ս�=���le��yU*)�>�na٭����D��A�K~�BBS�A������e�:�5kX*�l�.���ȢMU���k	������2�:	�@����s���ϪO0ɹ+��\�9��Y��a������FF$w8��dl��I��E���*���A��g�|4 �X���`�Q @>A@�B�Q�!�j���A�i��B8����9�;($�[�h�rᢗ|f��\��y����1�e�H?����D$ 7_�4��.�_���Ӧt���T(t�4�r�d�A��pd��}��\¡��'�\���ET��_B��$*FgFq;��Zo���V�M^p%����Z�o���Ǿ��û����a��D3ڸ��q�N+��[h%|��'��J���/U�b�㔈��O�S �	�gw��STL޿��T Up*�
�����ۧ�?�~]I`Z���u��H�8��_��oF���D��'xf�:h���-�b���yIH��(jی�M�q(o��5?~@_S��d>��d~����HF��(�m�B�5EY�gl�!���6��|ˍ�Va�	Eg�A���Z��֎�&P-����5*VW��$�6��;A@B��c| �<�N&̑�bDpl�i���Jб��O�9���`J��u?���M��$�yt�����|غ�����j��S���$\�w�]�j�<�$����G�$���t�7%�
yʅ�'g���G<���GY�eۨ�߻��=�	��o��(Lxn�YM�|M���w��C��P�B������͈jԂ@5[��R�I�ÿ�-<^G;@��%ذw�1vI� ��߱+�˰=&� ����4�����mk|��^7�l��fx;\��؆r�n����1��-�{4x⼿z{PZ����QIǚ�t��q�[xSz@u=��R򁍚V���^֮�{�HU9�rMg��/�� �D�:���p�.v��S2�����}��2��d-2>���y~/q��iqӖ����e�(�`qb�G����i�\��_���MwxC=�Pӷ	:���¯N?wz1��u�S`
KO��Wd�S���V����^en���,���r���8�����W��� ���_-�5�>Ve���v�ε�c_t��#r�V	"4^�`'-Үœ�c����:�~��&~gG�'ar��v=��ȯ^����ר��nm��l U � ����V7��N�dc~<nV�yacɑ�,�
�ۇ��y(�crFOX\78ϵ�'����K���M�9kʇ�B�N�x�E�4@5>��0}�C'��wɫГ��#d���}-��"M(�N�<���Amh�p*�$�Ad�{��8��<������ϫ�U��K.�ʍǊ����!�1�d=z�/���C�C�DP[�����t�P-��;�֮���;թ��Wd��0{[5n����z.2��lq��SZƱX�Pk���4��0��Hl�
'YH���ذ�&x�G�5l�Q�.��hR�5VN=-ց3S~Gl��Еbra޽�zX��-��E�3�RL�"�� ����~|6���m+EF�{5�����}�2:�P�u�z���vD�B���\F��
�}C/i�d�2x��rR�"oѿF>9A�����
xI�4$4Jy��e�1���z¶�IW[�D��P�a���
�nˌPPPP��S�[b*ڎժvB�Ċ�F'�p�R)�
�S_��=n=�8�����1��9��Wy�犵����f$��$R����SE�6��W�O��@G ��^���4�MEo	e����Ȼ[��ƶ��nL}��ĉ�:�>���X>t~+��ұEg�A,���t��K]��3�O��[���_"m��5��3W�_S0俇Q��y�]/fx�����s������UPF*�j�A��H����A��s���$BU��|�+K�?֔<���3��Xv&&76*���őz	������&�4���ƥ��#P�5�*�Y�SwM�tS����w��|I�6/��Bʢ`&$�r�N���6�	%�;&���>�P�U�+ktT�˲s�f�/ IZ�%m�59�:�-UPlua��m�$$1�Ǭ�B_I�k�z�L�l�w0x3�u.GKSB5�E�r�g�6��A1��jڦ�-uM�o�'"��Db�h3�>�Y7�`��m�aQO�� �$T�9�]@>w�ZCa]��gz��d1��j�>#}�X���.D���IX�e����Ϝ������M���Xjʟ6"?�H�SD��{#K{�@&��^�3�6$Y�`8�[�|��;����%'q���tO�ۅ�$wii�a���D�Vz
*#��s70�=�v� 5<�)��h`.A	��L�!F�v���%�s�^G�C��+.3�@Y���z�@GfN9��c�rR��K+Q�6C����BO+!&�^j�1��������-@3aD����J�Ğ���u���F �X���%�8����Y�$�6^E����D��c�@h�s��j������-��s�(�TL��?��� CP}���[�#�o�W\��}]���SMH���}4)����Ż�|�\J�g�(�l�ϒhyA<�S� ���'չVw�gr��aETܿat�w0��-��%Y���L�T#xFB*q��������o�祪�����HU�A���� z4mO�s�����i���e�Si�wh<���.���+\a�L��-P#����H'�{����p���1Y���������w�IÈ��J�rjvd�v@��v����nv����pjx
�F�������,�6l6uc8�I�I+��բ�g5���>U��t�?�0 �8OB�>(,�ȕF) L2�ʵzGdY��ڏxJ:/� J�$��z�X����X�_��΅���3m�i�^��dp-m�er���qY�'e�P��ā�0�#SL8��ʌ��Q[��_�s'0'�k�>����pB|�O=��a��~�)��aP�+�J���=hť�g�3sW�V�g�X�P`�{����ܒ�jC!؊6;�p�����
�Q�C�m��D��7"�m:�I"{6]��Ui��+�``�.X��_D!��W¸���f���8�)�s�ۓ.78��w��%�j�P����cNU�S����2�w)�F�
[�0�q>�J�nr��c g���:(���+,w"}��V�߰4ڎGw���_&�y}T�P���d���ҥ��F�������
#�V�Vx�We�$��Ѭj�����$�Ԡ�Eg���S?y��w�d~�x6@�|�K8���zt���,��T���%�ch�[��E�DFgD� ���,㾄�uD�Ld2������0Up��:�N�Ԏ}?b�%9O���sW	ȯ��Y�uo����-�Rv&1޺�C�w���8�,j��'M�r�ƑգG�m�TQ��&���W���<+v�*�KKf�?A�}��>�WdI��5�p�+�!�%j���(d�~^��RI�����w�^�U/d��\P�(؎gU��%�x�w��Fa���e �0�kr��"S����GD� Y�3$�I�>Nr��O��@�����]ᎎY��{����Ee�]6-6To �khd|��7�n��&��L��s�2L�b�뎨��VD���W�{�)%Ø�^���&N��������]�F�y���sm�g�[���>C�
�5�ѭњ���
���ȱ��tk ��З�9��l
�j����Q&� L�Y)����}�,�jq>L �3��$*������P�ul���W���n'����;u������'�����aE�mѰ�ze���K��jV:ȎW{>��i�P�����	��dc�f�I	w�M
-�,�d�-�[h�����#/��k��Ġ��p)�'����o�� �,A�sj�����1FV�(

ƒ}	���/%@-��yo8�MJ�#�>Y��Xl������}G��S���%�Xs.H�u�$�z�k�c"o~�d�Rv���r=�*�d�#����ȫY��G�,����m~�%�.�B���\"��l���0�J�q���ǝ��{��\��U�- @����zA�b�x���4%R�<֓�7t�*%�y��e��$r�K�r���qǭ�����m��<��b8�8^l�
�'�y�xGƱo��aS''��P��Fc��!�2V��������.�+1����[�G@0�-0��O�o�3�<�j4y�[a�'�#a��'a ��,���sX�=�ȓ0_d��k<��?pr*�7�@-�����β�*'���\��8�h�
�>T/�yZP.Wоy"�-$[�5���i�c��Za��{�|c�m��l�(�Zb9:���0kvFL|�F��t�B�\O�m]�Oi�G+�Ȃ���?#�H[$�5݄���VG��C
�-��[,��_a��=F@%Rw��n>�+��}��o�R$Ě�@[r�o�l�T}�9�.�5Kmh����h��<������M��)P�f6�Z�X����|sL>��闁��<����߃N��[�1j�/���,�,��Kگ�D��R��8�={�v�8cM&�^H����IᏨ� S�t�B��x�I�k_t5b_l�/�����_�^2���Z>f
̉<�m�r��HC��"_{�G
�X'���2��J��зb���߱)1E���D�����w-%�˸����;Y�ն���=�Yx��+���o5��q�7m<�(��2�����B:�P���~4K覧�>��ݲ�:���?�*i�⟂�2.V-r�S#���� ��#�_A9�=T�Of\?ʀW\�̪�Lo=\nX�Mm�a���M�i.!�4y�W���ѥ���BK�m�_`��F!���X����Ս|���=�4�3^g�9
x�������Q6� c��x���.�#$Ԁ���o�D�����ٙ`��\� �ڱyY��6y(�)�h��s<sq��oeV�ٶ��KP_s�?��J�ݘ/�=.W�*|�v��j��n�ӏWP�x>0b=~��$=(of׫�����1�B:�VM��n���rz1�GG�z���%������u��Aŝ�#�� EK�b�W���/�l⍁�Z�i�F�����R�g�����>	ɡ��y��0����{��2|�Y�=�04�q*�	I_x�p/&����8B�����"����w�"�K}xH]�h͞T�i��ׅ�p�㢆�\�8T� ٽ��n�1uQ�f�O�!�-��˗w�(�I&#��V|�R�v;l��]Qē�a4��aE�v���礿*,	!�H3���d%e�p_KE��J�ySWݓ���UOņ��>Gmܕ�H�qX߰q�2#%o��:�Kᑐ�{d���3����18.���3�B3W�g��xd���4ыz�]��]������)ź:���Z����6��_����^z�����c'&�A�z	���ŖS�5�Z�r�=y�H��n:
G\�˄EҜ�H��`�qڗ�m0["�����⮁ݼ�%ƣ۝�Q�8�)a���Fh�j�	�*ɬ�(�p��}�u1�� ^U����s�]�JgYvR�Ry�c�[�da�d�	�S�@
�Ҷ�^i�UX<sm�W��qS7��GEG&_S�5�gq�Dاmrz�b���z^b�y���F1װ���;�����3���fJcձ�HA�h(.9û��f�o�����7bٰ�<��#	��pzܣ��	~����کoh� ���5��f�q����UX��0�8���T��@J�AWߨ�}:M�чQ��`H�:�����We�"Y�\��E���@v�U)-~�5]��z6x�V���Q�؊I;7T�a�ج�;���Ԝ�&(�7?IsE�gA�DV?�H:��/"?\�J�.!�W C<˯�_�7|�T�G޵�v.ʵ�ݔ��̶S�<~$��u��+Hk�A�@�v{�ZfH����T��*��!���܂���2��!�D�,6��@7ò����;�0����?�I�Yz�r`��$[�&�����w`]?�G�6�$}Q#j����W��Qd�)��<�Zs(�0�N�U�(�A��o{�/�[7�Vgh������|Gn�/p	�1ha�<�཰)�F�G�y�L&����#z>>%?�WK����=������*q�[D�.{����b�x�v� ��Fo<h�?ʢ8��oL07{�mM��`��� �C[Zx�ͼ+�vy�F���@ދ������H�-��>r+���hK�S3���֘�ACv�y(��Y(��O�q�1#�)B�8XN����#|B�C�]{0����r���,�Rk�`�����:0��I+���n�~�!ht�IFˊ��b�o"0(�"�C&D�����q�*ZW;%��#�������I�w�6�"���w:�p�"�����'�{��mHG�I��1ظ���� 9�7v!�o13��N{�N&� �l�l�vgvz�O�����d*q(�y�3n�"3&4}5%am ��{d������(;��kQ-���9�g%��+e��?:�~VX��?�;���ȩ����/�uY������F�9� x9�����V�A�,	�K��l�&<��!�i�+� �o|Ya���G�/�������G*Em遈��������x����"��ÄqI���������z������I4&�)�I֒[�[6�Y���)0Id=B��|�����X�I�b��U*�	��C��]�:@���F�O�#Ť9���u�?@� E��r�����k�T�z�jL^��k�2�ȃ�Lr���"H�r<?ީ�e2�,�$�*���Y���!_B�5�����2�p!�4f5u�<�+%2��R͢Ɍ��5G��PX�1���$�,YZ㬣���4/0\?S����qT%o_�� 91�_�e�.�D�b����� q�-����\��l�(�#ߵ���W�:��kuZ��$WU��4�x�m�t;-�����4�L��m�A������7���/��+V�i'�BR��C��YTM��W�����{��ꬋ~�|���u|�\K�6����?�؜�L�R#�ͭ�a�7u[eF�P�۱�ܟ�/RM�1������T��e�������{.�,I^����/�����;�*�����	�&c�˳.��_��Dy~K3*܎
[��X:��X�AO���^P��`�W���ԏȇ�W
T|�?���)^������L���ǧ�9� �4��e!�mk���s'V�O��X� �K���V��u�ğ��kQ���a!6	��I�QGYEO!2�I��kL�������Vw�:�^ԡ#۶�T۶VǠ�������Z5e���6��R�� Ǆ_��ܲ��ȾO�����h',4��!Y�،�i4&��! ��7ka�$,?����S������Q:3�!|V��A� �����+���}�=@p�Z�e� ��V��I��)����z�`�5_|P�N9��p�|b���ۚ�����)<p�;ȠEb�1�+���X�x��2�~���+�e��}n��ڻo=jEօq�4ď�`A�P�ț�r�� ۻ���GA�_m�\��g'g���A��yBC����m��G��-C/�&V�&��N?�E������Ч��VgI�������l66���
f�8�ojm~����i�Zqڕo�ܔ�+�eN�}�?�7���U�8��+4�bO�<w�K��;%����ȄqgY����i����o��>�KĎ��d�X�4���u�K�g'jG6�ή-T=������׮���U�آ���xnڃ�՚;�Q��L�)�P�5���S+�W�(
	�� <�a,v>�R�:��p�&g%E�B,�vp�NS��&��PSp���{�����QC���D��Rnݡ�+�+��	{l�g'�/��eX1`����Ћ����hW2�Ҽ4��@yR��Y2t����Gd\�������m*���?�o���4���S�~�5-~ۃ��[�����2:f�"�(��ҽ>P����9���7�v�XV��mk�ɋ�+i�g_%���$gf�İ�?�H�v�����Gԁ���T5����'�FU��&�6��)S����6�@6���f��
�$��b�8���:�:�h�Rnԃ���ѵ�h��Y��th*�ܖ����4-��yʬ.���%o|�HoL���̒����*���#�3n�f��B����O���~8�i��a�x�)7��y�O�&5�^��V��5'�X�W�`����;�<���;j���b������Z�rH>+Us��!_j$�e����~;SH�ZZ�J����q���	�=�.Q5���<�Zg�"�i4ښ��1��o��r��Ųޝ	�b"�~#'��؎�]�t3CBEi�M�O#
��s�It��{y���]�m83B�zk�i�`>,�eQ� ���U�/�K�8�QmT��P�e����:
[���a�T+
���Ew�:���q@7��t�� mg�,�j``z�9w���A���X�����)�|�촾��ֆ^M��zf]{��ф��X$�B OӘ�.æj2ֺ�o=?k�;��T�#ދb���A��$�"չ;��Q�ԋ�4j�ݗ!u����׀��]l�B��Ƴ��fb��O�!����y���Fy ��u}����j8�r�Z�{؊kU}�v�sS��������j�m!'\Mգ�:���q������huu���~_  ������ո��v�e�#T��A)�S�/�]���n>ò|��<���RIX���1�g��`�.���׊*!
�h �p��x�($�C��o�ہܒ�����! �Cj8���SGB
;C�(� e��#��tڏ_0�i��
D��uz���C��[u��8��ݚ8Sp�*�G�����cs��drz�'���z���ks�w;#����+n�zi_
�u3�g����6��"kI�!�F�����i�	1�78�����Xp�B�VZ=���ɿh��Gp�7f�'<���c�Ц�OMӜ w��+����Յ?�Hx�oA�'�݌C�·�Rp��5����'��}5ެ �
A%���iH���	�zz%���&���Qxp?b>XǮh��>i�"����	&�f��|[�,�iM���16���b7s��'���i&��y��s�#�r�!`���NsZ͛Fe"�S��H�Uڰq�a^�f�,#m�hݦ�u���8��� �Q�<���%�����I8�bk�����t��	��UjMi���1�o�V2Ig=ڮU��"{W`*)�x�Ց
�<�4&#]�6�Ԅ[c�f�V��4�M���	�O�����+RYڨ�]��D�iG��G0o�uu�џr�I �[���M�ߞJ4q�<�<��1�)��uh����F�g�ez�[��b��a|���͎-ILy6g t�³�$֯Tc� yF�z����^�:d7S�'����\�ǽ�@�[-@00^. �59�֭������(V9�c�M�ȴЩ�>/rtl�F �*��E�Ʒ�(B�W��Ǳ�;�|'�W�#i� ��5�n�j�na1QC:L����7�ӻC���=�(O�7I����q<�s���#8�;�"����L(?��t�k4�e����T^-pc
�y����J5���;׾�(2\��7��>��k6i�RA�Qg��X��І��6��<��m0��*ȿ|=O���r4M�_���
�-����9��,�G��yF$p�썔DR)���6��/ ���blO���y,U��gp��.�
�[[��l:��+����n2�S��[��b\���_�m0�"T/"�ɘ��cX&0̓��Î�^���a���G�=�2�=�`��?�;^FN�o�=C{�Yފ%���@CX�H��߻���L��DL1�,h�[�0�+�k+߿��C�|�̭�rs.p炌�������I��o���;����*�VOyC�!���<����:
9:��Z=����K��ջ�iw-��WX������8J*��������IZ��nĹw�fA)�	]]���&�u����ZB��R��Eݴ�c:�?��� �,:=O��TO�����&fm�	#�w0�٬��`����㽘�!���$���I<��M�=Y�w�ՠ���.=�����H�ėpQ��,���đ�����;�r�V��'�9&3�個部��ɼ���L�I�ޟ���+�����Z��eʮ	П��./EJr1��ܠ�y�w���8?4pf��,���!j&9���h~�(�<&�jFڤ�M�͖J�x�vp?w�Z�&p=�,���M�|�ԑר�4V+�O�Ù�/��ʢ�h?�u��H�Y�a��$l��0& ����B����>���F���A�S+K�ҧu�z�OAQ,_~(+./ow�)�{𤤸��S�Dfq�GP���U��0ͼQ�ވi$8����eE&����g�AS7�r7Q��Q^g���d��Ǣ!y��p\$�.���/��
z4�����+�lӎ<�2wE���7I�А�ڽ�w
&XFB�P���S�G?��,��՟'0���S�*±���#��p�F��[����c#X�dRnق�u4�H�ml�Π�cǥd(P��i0{��-�ؔ�`{|�Ӆ#7Ȯ��s����B����[bf�G�9=Ic���+�z�[r��gn���x�i���忣m�p�B���Fh)|/U�����_��ʸ���E����)���`�`H�p�4� s�# [zYTơ�m.���q1�S&�J�у��Y���l���\�� ���uA�V"5�qIY�tT�R��I#����u��(�.G�����ϷK��S�&���Id@y#+\Z�Ƕ�@���D�������ce[�)e��1S�ok�tZ.+�X��h���ȹPO�$��i�ȷr����:�iY�����\ s|���v]���V.��iM,R鎾k��+K�"�������x-_(���&�����/5��3��࿚π���W���6Kz�x�/���X�JE)x/�2�4�*rXOȆaR��sǻ��	�]��7S���G�� u2;��P~���Ę~���9M~��]����Wb�����S�x> ��v\e�a�X����i|1��V��ȁ���㵔��8�J���d���꧋���u�6i��KI!��s &�����9�X�J��_ur�fZY�:�)��kp!
� GR�>1m�����(������ɏ�x"��:5ϒ�b��2p%�����[�*e�`RUL���e�b	�e�kfV�O�fKG��ڍzt���
��ǣ6�u=�nZ����}I���xF*k���VX���A6�����f-��Tu|R�|��_D�
�n��qU�[Y�b�3^�����`����1�?�k���X�S�_2�(\B�,Cg�h��((t�Al�pK�l�㦔53��FQʭL��Fk;��M�
�A��Y����"$���2U��(�w���M�#!��d��a8~�5"�20��jBۍ����V]��N�p�2&��~f�&��m�r��cfSBHͧ��8��w�K�Ig�*Y�ڹلBOAˌ�0uK��c4�Txth>}�ջ��۾(����l{?"����ۂУ�9A���t�s��x���T!��
\MH��:�v�#��6؝R]b�;�Bze�{����#o���^�4˱�s�@�DB(ʌ���t ��]��
�š5ʸe�1w���b9��<#���әW)j�ռ��d�qC�nr�y֧�?�~z�T��Z�h�ԛ�N�X��\��C�<e���ao���5��h�C�"�ňJh|Pǝ�:�u���t��Q
�m;��w`�j���[fM�*�<�e�~��������O|㯒�O���@㷓��<�+�4�����|W�䢺�X�L�7�]�܍�O��b�E�q��5��zÞ��)�ʂ��3��4�G��C?NM�]"��*�d�/m:���������9J/��g�8�[�"��#F�	�ޗ�. ��5d���C,/Xr��q�ְ���w7�c2R���1��1����J��� �f��L��r�7�h�ީu>� \Ť�O{lXz��Fb�7n��f"A��d�����Fφ#�����r�}���Yw����igL��#[�QK�J� B�?jU�ů���0M�7�JML�O�
._�q�&ѭ�}K9$� �һ�1�����0�"��W΋R���92:
x�Bdܛ:D#��R!�~�n��چ|�C�#�U� S�I[� 7�K�ա5�C����X���9�z6"r*=*�B��e�׺D���wf����RTU��Ҫj���B8�)��ȓh�d��?����Ƥ���9������MB�*��6H�n-C
���j6[]����������le���/s�O�u��Q�w�X���-���Dy'�j}��lǫ��6[$4�$�@j�9��L�Dt���HD�>S8E����@���A�n��C}
��eCm�A�FW3&����B���+�����&D{.>��:?qH�Cz���dp۔z���5~_�0Pc�FG�2(��E6H�)�w*���@w8K˚��mgR�Pd�͜��˓W���|\�`)|ݍͽP�ُ����S�1j88m�Z��r����*� ��e�`�\�&�]���y��L���5g�=`�N�d�����a�aHcL��0�Fn��N3��pRʇ.>�$�׉�bi˩� ��h���L�;�Rd.x�^���3�l��JKK�#Ѐ�pn7�`����+U�ͺ�t5�~���fe����(ٖb^�B����S�/���8��'��W䟊��.3�w����|�e ��U�c��_����;�n�~JI�̟jYK���~�����I��%��l�p%���F :���]``�J�����V<b%�Ē��;̬���|����R��3L7$�%k#D�m�_��WV�{�?�{Ф�<L�f�_8������Hݔ���{Y:_.�P���9*��P��W��M�����|T��+t�)v �u�C�ji:e<���P�l)�Я.�p��p�8r7o�/Y:�M����+�M+X���Z���uk�g\����RF����z�J�ʐd�oa�~R32��[��Z�j�9�ݐ�,�>�ˊ�RR��/s,�O����O�QV{_�T	�!G؀2V�ʳN!��`��~�l���|7�"�a��t\�qz�����a$`�)����fy�.��E�hw�#�'Vc%��X��*4��E�;I!�գ��Q�TC&�D+V��]��^x�T�n�nH|����u��?%��w� 9��ܦ�t��YzK��tC��k�˻��W�ʋ'#߈6�7,��uCa�)D&"�	�")u����W}�
3��<D�ݳ떞cn��	:
%�`�7?����R���A���ie�%���w�ӦPA"d@�8.�t���U�S�C��i��'�]8��-�.��5�������GjWA0v�W���V�!�u�������8Ê��pcT�R*-���t��844��0�K7�u���·N���'�,����b{�T�g��B��g���c31��>D�Q-�t���:҅��gÎ6OI%R��۽�{C�g.|������ZW��uD��6����[��~%�Vo[뢘����&���8[�~@3`�%�N�D|�	0t��|�~�GgO��8l�w�S"'�8��r�/;��=�d�ñ���6�#�o72��Q6�*���ҿR�X9�e@�����tÒ��bѥo��Dg�$�2�'�t?s�#Z�hѪ�U0���+3�)/jXi ���[����Fbr
�j�{�P#��E�����V�_`��8�]3{��C�{�f:�3��=|��Lm���6�g���vdO��'D���ch��8��o�h�j.��/x��
���b�R\�C�hwW�P�����w��/��L���Uey�&��?��PwSHteP�+֣���F$T�*��.|�_9�v~O��G�:b'ɘ_��@�:������7����M+�S�DAr��Ǒ���)�%NT��t��U�t(�z�AMh�(���p|{0H��h$L�H\��߁Җ�>��F��#�>�_�/^�	uC4��pt�ya��ay�u�16���D^�l'���������W<����@�dDt1_�{+�+̆ޥ�A�rw��"	��,Й5�6���M!�ZzL�!)�B��;a�s�Rĝ�ےC�ĝ'���HYYN��
�v�����1؅.�vX1(��ed78Z���x��<��ۋ�P>��I5��R��MW+�1�U_`0h��V��a�-�C��<f	�A����oӵ���l��W�2Q��T��-���V*l+��Z��w�N�<;���Қj���ȥ�J��&/*��+r�*���j���R�`w����b�~>q�.0�i� D�N�����Q7�O��-J�٧����>�71��4Mgge����sD�����>�݊P�Ů7�ߣ16�Ȑትt����G!��1A�ܭq7��Gvx\�}�~�Z�G�z;H���a��V��(h��ӷw:��.[��s6]]���ďZ	j�V۠���g8Y�wN�Ib\���a>#�l�a�grbdXc�L�|̀2���?���D�� �U��g_�*S,�����aa=U
miAo`Չ["F��\�EtiM����qKe��#�pT�����9����`��i	�?Zh��VU���?�AP��mB�Ax4#�H�G��6��x"�x�6dyE�S�JLS�?�"�'*��{a����x���֙��)�ih���*�=�b|԰dN����C'��� ^I�c�|Ճ(��-K�P;%+&������,>NX��x.�/<�zhP�b*�6͏֏덚g"�uFE77��2����f&Έ���6h�3���3���ե�$�߯ex���51�V��q�я`K�nz�h����"����8F ՗g��Fg(耎N_D
�T���� �ycʁ��n�́,ܭ���W���w�c"������а�g/ߋ�	��H�6t҅�{��>~�c�%��z��)�Y�aG9~ډ\�ao�/�C��ӂn�}�������w��=�k�$l��䚉򴡻�xNÔ�n��)�r^2�k:{pE�E�� �/<�`:I�U8A�5��q�ȅ9$D��0r�<�H�#�=�����^��Zf\$��M���B�����Ǜ-�A;q�u�NI�����)�=�D�_No�ֽUfH�,�x�(f�%���{	���c�˺S^�ܥ������X�&����ՄL#6�p{6|e��?�R�����0���l�w��t��F���|ud,�VU���-^��dq�tM�'��Z�d^����*Ѿo��K+9yd旀� ��gw>��a�̴%��QZ�13���	Ov+�'���s7֣�/%U�^�#�7��d�w]��h�� �lb4ڛ����.T�`����,��$21��B�������X�Ԙset^���;%߁9�оW/��-�g}��:QZ�C
��&�+)Ww�ڂ&��WA D>z�Zrv��g����޼f����������u�j��]�8��38K[�c�󘯼��9Ō���-!���C�L�}��hs^�}�2�t/�&fG�z��>}?\��`�̴�n�F_{@J�e���c\|E[��I��;�R�#w��~VW~��S!ȣ�`c�?�$�ӏ���!�X�ϻ�.���"�� �B��0b��Sd���4�����}b2hS��̌��ɧ&n�`�9��[�s7F��ܦ�6	���Zx�>B,%0���?~����;Ђ�O�'�󈹝Q��i������;f��@T&;�@��z`K�S�����a�ka#�f&>+7��˭�l�'(9�9��*sFA�3�Ǌ4�gI4�S�'�j��B����+�pZߵ�\��q�a'�']�Nf33���Dd>�c��K�r��s�رzrr���sQ���9�盟�Y�P����4�0r��)��E㰀?fE�]�Rb�PN ��\�z�Gr�&2�>��ʵ��wC8y޵oH)�?ø�q�:*�@%�Ģ�L�ŲP�G=_�#��nB⏵|��V^/f���u�?���<%�T%k�F�f��U
&&\���F�,L;�8ׂJ�����%����d@���T�Dakx�V*�������l@����&kJ��;�.w.��@h'��6��V ;����qlk�ұ�X,�s0�[  F���y����@3J�1!��$ n@U	ڎ��F�p�O�S]��.����?L5N�u� �V�03���b�D�b�P+��"oK�Z��'o
G���qw3�����q>��{�~IN�[�����P�o�)!i���dH�5�T�N�����4�>P��9��X&V/U���(���������K}���HN,�����X���(���Ma��hy��D�Kǰ���Ճ��!$T5��vW�<筏�OX����*@C�0+�)�(/Ơ������L�Euʄ�ŉ`)8:~��
��윩-oP�p�)�����nqԼ
ԟ�q*lb�ٔ^�@U��A>��{f� BPt����v(��%�#�4��Ds�@/>4�p1?t�N��X�[���]Yh� �P�d(�F��g���^��GX�f�������>)-fljF�]��1G�}��w��5�T?�y)�z_�(;c s FL��yJ���v��pZ���b�嘈���P'>�4�6g�ض)��-n��ن&�0�cg�)�5m�A|]��^���ݾ���H���TXq��<-�J($S%չ����r�@�Ik��!%B|��Y�5�F��L�
�� ���àv;!��J)�m9
;6�~�^֠�V"�4�P"|!й�̤L�.�F��2<ØtSr�ɢ�`9$<��T�`P��ñ4w"==�3�QU�K�X��y��ұw0�(�v�A���4��O�f�Ur�>N��Q���˛Lp��6���P���fD�i����%ر 4��l�<.��*%P�˫�����m)��y����>dۻ���������BV���ź��aZ�J#�=��l5�Wo���R:���Б�9$�>eL�a�W�w)F No�X�Tɾ<�r�$x���O> G��*L�wȎ�Irb��{�����T�3<���%<���{�-,���F�F$��R��eY�����b�v�(5�0����F�n>����� 趄D�#a{L;��,��ְ��dE�49��;慃��8��7z-؃tX��豢lĥ�Z�VF��Y+*f.��K&x�j��WK�ϣ���g�_�lYo</C�*^�����=��_z�X���>7�:�n�y3�c�O��8�uS���T�5Ӄ���I}N^��m%���z^��
X�l�z`p���.��j��ul�``%�0=��"8��a������]T�!�
u�)�@9~/��i�|<(>���R�5G�N8����(��l|��ptB�w�Bq���*{
~u��!ҎKGk�^2��r*7D�~��J�π1& ��*��� �0��JR��o1Ey]ʕ�����ϰ�(O�ʙ/l�͚����_R�7SeҦ�����Sa�+��N^yx¹.J#�����8`����y��3�=k�bs�囜 Y�;�ڂi&�f=�N�S\���uc�P����.#�Y�r�O���q��[Z Zۺ��;H�o�3*���zhec�h�ᵌ�I��dDhֲc#��`I:�+�JK�0�
�(�=���x�8y/���`�!�P��Ɂ��m��\�+Tp,G)��YS�-��"�T��������b
D�!�ꦴ�j�Ev$4���ωc��u`��q�!�DЁ�'"+H�(�%��w��9 C-��8�����'�r;�֦4\� N	p=E����`�FV�)Ri�i
q���O9��#�uqV%2C4h�����|X�##]K������˶߱Ԛ��3c��E��;�\�n>�I�s���������Qc�
Y�y�!�O˖�.j~)����b���Լ*N���G�I��+���IA^�U:��$�w�V��)�������w��$���M�'�/@,r�,K)~�{�x��Fh��J����y,��&o� 计>�s�5�oM4k��ɕ��ѧ�乊�n�嘷z֟M��|��gk�~U��^x�:)�,��Ճ��|=�߷�tQ�P˹sṜE�Æ5���ŵ;���!d?	:M�O�A
�a[���N��f��}�Mg�)��)� �|�Nx�hV�M�Pw���$4%���#N��CsV��\��C��(1���/"V\���fVG����qC��S��q�\�O��t�ڈw�cJ�.5�b�߰C�Kf5�/��6H����n�R���Ȟ8���k��z����$�&\ܩ�W�DYě^�co����tz�����sb�'�ቚ!���5jM�b@��ޏ
�:�h�ԞS�|HFzG�/ٴX�Sq�0
�1��������kk~�"���Dߖ�	�z[���2�+��5z�x�'�e����cgz�D0�+ݰB���te���
�[0-I�p'J)��O�Θ��HyJ�I*0�T7���W�6�;+�B+�\y-�ق�؋T��8���]��lG7!9��6~�	A���FNs洴%��u�xR���
[�L]����V�O���a|^��n�҄�R/P�mg�`���Z�0YL*�F~}�7ƥI�}`�&z�'E�8QOV�Ly�w�jx?Wa�P;&*^�Fb�$��aGt�hn鐦�X� ��ٔ�F����3���	�Y���tS��2ݰO����C0h[8�C:�/�l	Ѵ����-�>_59�'6"�����2w�-BV^M�x���}�5%\�O����V턋.��׋�юp���;�D�����y�� Z�bz��seL5�pR�A�گ��M�e����I��ie���}hNٚ�m����9�5P0c�%�_Zuj,
=d9�@�����9��$�(�Ր�Q������Q�L	alguy��_T��H;���'$�;x1�
�3�m�\MW��m��GT[h{i�0K��.R{&2����Wl�6;$�)~����Qa�z9%ƙ_vm5�jB8�+�)�A adeꃜ=~#ް�g<��`�ۋ77C,��v�;�h�R֝�N�4��J�t}���+���^�|�&�g�6���֧�=��ѓ�pһ����#뜱dS�|9b�����������g?�D�Q�Ñ~�UT��x��`�axk��9���W8X�`�ǰ|#�ɬޠ1�.��,� 2Q��Y�Ŀ`� �
�z,j�Ke���=�T.�V\��'KĶ�e��%+�&�t�����P59�(�tH��D>8���;��yi�F�'_�e�x�n��G��p|/09wM��d�0��q��W�o�6UV���5Wt|�GX|�J~ؒ��)r�m���b(�4�(>�Gb�z�}<�ɶZ#;���NZ�� ��?���CC�>U������t�y4��,G����ͮGC7�I���
��ɦ0rE�r�9+����ꢂ�Mȥ�����nD5Q���ˡ7S}�n��:'��,�����z�P}�-����0M�v;Gݢ0��4�cT�$8�� �@&���>.��i���P���'���?�ơ��ٱ���n�1I��������Iw���M,��6a�,N�Z%_8o�9��:�jp�¡2`�T��#�V�_$ߘ�&���s��d�	4�I�8G7������)2M)C��J���f��o�c*NI �07U��B�͟)��n�R��WO5@r�s�zM��[��Lٙ���f�j`E�	�-� I�z2�T��`��&��^��������Ү������szz��9��xM;��0����u]B�Z��*v�`�#J��]� ��<p1场��1c�q4�6�(��x��E�5���5R(Y%��Ot��d�%���MqPcV����4m�z����s�N�����z�5��p�s�ϖa],s}�D$�y-��f����� q?���V�)VJ�S��Ҩ6�e���U��= �9[y��0����e\,g"�U�|������C��O gi�ԢJ���%�  ȗ���75��&��L3r	�v? ��|�,��*��|����3Bp��1�X԰n�?���A	
��"S���`fYW_��MS���⦭�lv>ӫ�^	���]��.�!���� ���p�7nջZ�᳃Z쨓h/QL|��J�*Gz嫖@����:���0�n35ok�@E�x\�S��7�,�E�j����9���-/�zO25%q`xp<�Zo���b�@�����(3l�`��H0�``�5�}W�e�����=E_^䓇~}v��\�����.xe~Η��ŀ����S����T}Ș������E�	�1i`�D�e���*�ą�XGO9y�9�}��bZL�Q4���74�7� y��>��_�.)Y�W���c��R�Z�i֡���7*1Pב����(��h|�k��%!���Z�h�2��#O�ru俚�W�WgK
:��$�i��#.�o��������%"(B�A�����S�@ꪲ25���=-�X�U��VaQiT�! n���k繘s���U���x�<D�5�t��?D+���C��%�]��%�h�N�y���n3��,Z;�i� Q���=���Д�r�����5�S�%W�}�~Vu0��Mz�A�U8�,L�\(dyZ�*r9S��Y�(�h��R� �_:ʵ�6~G���")q�h���I8��a૑UU׮����txԐү��S6v����"Cs�s��ٯY�3?]�g�����}O&���,^9��9L1���0ҕbb7`�şW�>�/>���V\d�E���l�J+��`݃7���.�!��]��W���$J�`�������M��a;&i��P6;��;�"�-��	�����ս�JU��H����L!*�~�ΛV㊨�_��ţ*��N�F��)e?��O�k]��杵p6xY�=v)#�ۡ�K����~��Oo����T��'r�CNt-���b�N�"�E$�w�B�%�C�[G�=,}�W/��H=�ʏ��E"�I���zm���zi[��c���S�f�^~����q$�T���a�FxE��"s���@˯v�P�3i���N^��L�x6�T�?�_�ӺV9�|���D*�����j��D/�x�߲m�$�R��Ѣ����C�&M��;栂��m~�t�	��bܳ�3�@j��E-	8�=�!�;P����}oz�#���G@�2w*�,z �6��p���ˌ�ɯ0.i�M����!���mxizT�+�}����9*�C�^�oi�<�P�"�9��T����Jյ��q{i�aWl�1��%��V>3��a>��\�X�ʄF��S�򤩾��<n�/s�@js��t <�4�%{gxL�b�βhA �J�_b� �03�2�Kw�F��!����b��P��𰯇�}��h�!JL8�T��U�Ϫ�.b��K����,�;��Xl:���R���a�o#C��}������U/��3G��E��^o��/�mܱ��
�d�3�s/S�t~�EB�0"\�t��l�+�x�WO��ϟ����ph<�È�� ���-��q�����	�=����7= �O�����,�PU����5�����7x Ѿ�΅���	�����O
� ��ƅ��<��LZ�]bdM3(��{U���J["�z��� Y�Ρz�V�D
U	�G ���?��oP��Իz=�d��#�~����j�󹺯`���u�B��g6���gUĆbX�#��aC�-g���sʣbY����׳Pb�k�����5|H�}A3��l���r`P�n�gV<W��x��)F�OLQ}�V5�^y?4�������0HE���#Ze:-�Z�xZ�	:�Xt�ݓ�Gs���ú�H}�>R�=�2�[�ǷV�n3\�otI~�our�-c���*�J��ȗ��-5;%w�����"�{a�{�&�菾`���$��K��8����R�BZ��Wa�y!��:5��z�#�W������>>o��E�/q=��Ȓ"��� C��\A���iM���j�<QwT˜��JW �ʽ��h��uf�	x%C�L�F>!���_"���:p��F�O"f�w�7��4#V�'��5�?�����F̊3�eFu"la8��}��}�{���@Ȓo0]D�N�Χ��v���>�`��|u'A������%�C���T�5������Xv�a�G����shc� 5WN�b
�R�Mx���}����n�2�[�pQ���	D����B��T��!N�sq���ݰ��-��#�79\���8�D�NT܌=���ΟN��C��̾xގ�=�J1K�M�|�M%Ǝ�|�Z��5��s-9'�_�ʽ��P��@�z	×+��ӝ3�.�AR�AF%Psq�/d�Ju�"���	�N�s���@0�Ďb�9pj�\�H'�i�2'�!�|H�m�w�W���k������@윀�LK�3s���>��mq�Sp\�Ta��G�{���_����ˇ%'�}�{�¾�Y���Nٰ��e�H�0�(:�j�L]g?ܼ�e���Q;�)��Oƈ(
��l��%�7a�.���$x���5�,S�0[Tb�2Lo��w���%ot>`�#�,��Qtq���6Y��A�\!���[mZ��B/{�Y�������kn.�1�/�L٣E R�Sҿ�p?����-�8cI6r�8����E�7��9j�s���|8�M�Y��עn�d�2�k5�kW&4���5�Hy����2���X�}��qA�/k�3��Ќ�\k��"�h:<�Cp�w��������t<���j��fQǹ
�@�R�4��x|,_tL�@�ۘB�YߒQnC�KV�Ia�["��)��	�2l6RųP��K�{��Wiŋa�1��P�T@Y�n�)l�ǈM��p��f"ǡ�j	�U��e%�?��>��dl�A��3+Ǆ;wl��<���lv�>��l���ԝ? q�<��Z��r��^���<�Q�Z;!�4[a���MsX�-���p��d�z�?9fP�`�i>ܟ=���V�5l=D;	#�����9:�(x�C��G���DQ��S�$]���v^��V�BtqM5H�ӵ��7�Z
Y�b&ɚ�O�	�u�V ]ޑɍ�� �4F���D� �QH>��H!ܶLŖ�=�)*_��L0
���#y���Tno.Z��_v!4I��$i�~k�GP��%L1�,�Ia���ziV�ab�#	�Av�',��Ӽ�O�[���k;�݌�1��߷�F�I�~���S9`���2$^��T��*6J!"�8�S3Uh' +S���?������uM�/�hv.�oEE�M?{�u�bqA�/9�`��oV��k�˹q�f��C�;�)�~�sݚ��sEbk�����D�O`%���@p�X���!0C�6�Ą��?D�ZԌ3
ڷRF�𪀞�$I-N$~�r�&�!�n3�X��?&x�����l��Eg/�{�E�A�Q=�M�
z(KՂOZ\�؂he��j��^�bh����E٘R���85�ػjy��Ӷ�	�ڦ<�����G(��p,�k��c��պ�V���
�lr����=��ݥ�&�=�Z��[OmŲ�8������;9�Ĵi2�����n!�vֶ7$��J*��-/v0.đ��!��
��v|�=�8�/%��ME-j?'�C�;���G��ŗ�2������cB8&�*����o՜̅W�f=k	2f҈E鿰Ʊ��PZ�� }'p�͟����ۘ.Q��">bZu�� ƭ�2��7+qc���|׬o��D�w��
��|��(��։���D��I1�z-�8�/�2#�S�L�v�� ���Ǟw+���m�;3��k!v�+%Jae�*9�v?B��5*X���4��(a��-�Iw�0du{�1��7�=8�}��kg��YE���#o�+V(i,vy��ܔ��0w�&���jw"����xd��/��\�9(e��n��������>�n��@���x\�D���"�:�}K�v�:P�J��M�ˇ�!P0�dva�Όy/K˴J&�3K^��W�Yv�������D�N�,acҙ޾��[Bs�:W��;-�-� �QE�4�{\�B#4�Ù���y!C���!��1(y=�u����h>�����5a���R�:�3�s�ݨ Y2���΃B�.x��f�n��5^��&o\�[�{4g	b+M�2�\�P D!��҂�;��'ʀ[�Bx3Ǹ�a�0.��In�5��
T�s&Կ��� Up�^�z�B�3���g�f���E�����M���5Γj�dZ�VO�i��t��X�q��#�P�f�(1x�Vs�U��A�g�?�����Ձ*{cL�,�E����޸w��{��7��+���~0IT��&)hV=��e�SaADNϪ������I[^�_����G�ݢ���}ߡ8���*a$y�+���0ˊw=���onA����<a���p�C��:~V�P���Q_�n��T��A ,�H��j�eG{8��M{czrU�PY"
�T.=W �}z䅚��h�!��Q�!��%��X�K|�/��+��0&�McGB�B�>���vG�����Kҭp�ď��"E�Q41S��o�H���	`s��p�/ޖQh�]�^GLO!���Cܛ�*�� ����_ܝq5�"H��!AH�Ъ7=�3f��f��QF�i�1TKV�	�Z���ؔx��&��I� �DU���-X�[�2�\y�.��m�����<
�0���`[{UW���ƾ8���(�ߡ�o��3���+V��(���u�7�-�Tț�Q��n	H��&2���qY%�3���l3juj��8On����}3�po�I��Rq��: ��Ì1�Z|�[�]�~�0 B9����d�i���4)y�kͿ�C��)�]�p*��b�:c4��D��T>�`�b#�ɯ��.&��t\r�|�8}��	��\�X�O�JY�fX�NX���r��1v�N����AO�rY\b�dm-�%i;cg�4��Z�qR8�5�����	����l�wEB
��9X��q�K�S�ps]����k@�N)H3�l6�>1M�Er��r���U���7m��֘�Ob��\���P�N��h�l�0�L�O�
��U�� <��e�9�Ce���VqG�}Ǡz��2g�?��F��԰��FC3zA%avܮ��g!��$L\�u�?9b<LGn���/Q]��wI��U:0��+6�@Wե8hĨ�3ΜAXi�M�ä'���l�NbdՆݵ���T�Y�R�uR����Ũ��E6J���mÿM`�lbb(�4�O����%���Yh��?ͷS�}W2{�1���<�h_���m}6,m�L}�M9h"��?�;�*GG�b;T�wH䖿��Ӄ����~���F���$2�h�Cl�t+�4#�5�Gyc�=�+y\���iD):i����Al �]�!���IV��`j|䝖��1n�ּ�
�p=G"�g\؈�.��M	z,�3
#rJ�\~��%�;8$2"�﬊��� R�1��}k���bz�%WCRˎ�E\��B~���=%�Ǯi&6�"��	����5c%/�w���?J��s��C(�/{�m��"&��x�p��7av�~�B�V.^w�󤭗a���_,@;��C�i��r��P�iA'X=4�:V���o�`-~AR�J��7�3T�M	��O9P�jB-��j�ë��ھ@#�� �HG^����(�J�N��U��Ĩ�J=]�(�ȃ�7�)FO����n"�~����K���@g��?����ezG ��
5x'�����>���Tp��<�"s��t�y�5�W�y2D!mjX�P�ѦS\'C@6�[��	D�}���_��#d�K��X��|��T�1٪��b74 y��8��)�����f��B�r���N�4��`ϧxQ����h������_1�J�[�K*L3�:�o��ad|�S]�-^遢2M[���,u3���I]�ߏh	2�J�R/]�Հo��͖��Jz�V�=*D��U�*j��N��/�n��YR[�W0��9�g���tC�`���W�3�E=_q��N�I�}������G�:^�zh�@\#�s�G|m5���D+�;�b_ܮ�tz�'�Ȭ�j���-�������՜��􂂥J�)i��$����'�,(+��șڽ_���)uޭ</`)NA�l:��0m���1S=�"��7��6F�$��I9b����6*��g/,����q���{���~�����O^x��9��M�@}?��~���]��XG�Uv �8Ǳc���������n�o$>���߃�_/��i�i����J��^\��/���C'��z���1V����{�	���Ks�\��¿�,�*SS���u��
_��l���.�����ʸaܯa$R�#m�	��or-���0�����Ź���f�xU�z��)���Ȧ�U��	Uq�?mMH�59%V���Rz��c��|��GYj������գ��l���n�⮼R�nZ�u�}���}�*���� ���6۞�p���ȉ��v�%Qhr�9N=[gL"�Z�����?8���J�~+���+w���W��{������j�8j��	܇���܍��X�3�Z\4N����Ua�}����U��^7 �5���/��g���	J�/�Ez+\W}�crVם� _��@dz��|v<�u�B͹�Q3`Re+��c����||�WN��؜�!*�����1wh��"�@�AnU�";�ͷЍ�����`�N8�|�Bi�V��ʬ�VqnL-
ߜ���gT��������$���&J�3ĝ G��)� �Y$�z���íj��s/�_�6�_#�,��%mjQ���p�SY�o�Bj�v�lb�v ���MX�O|�"qyd3y�d�|���|kjX��ּShW<�S�������u������1:����Ux��.i1z����#r�E�8|�k��<nJ�-���v+���#�u��G�p:�Nz�+�@���q����5�Wʯӥ�k�\P��ve|R;>&�S�>K��蔜��)����m)�o5N°)/W�i��۫󁙹9�)9�<�H9hЂ�a�a��H����~̨`=�?
y�/L_��@wc,+TM�.N?T0��$���΢��,����ϚF���]˖�����N^�e��qS�R�AR�y^��rh����+����|� C�[�<���
)I��u�����d�qQ���M������B�*/n��Du~�cS+�U��+=5�W��-��)iy"7�E�/����]���qV�x��_%���(x���
������� VL�����:��ُ+п�Z�f�Y��>k��pW6�rP�I+�R����7֭H1�R���o�9���̒��~:�_��@Ǻ�>m�,'�ҋ.�w+�y4pjE�!��q�Tp��(��Ǽ�))�0���pL�������Y������j���;m�NjH���zniL�\�9���Ȏ�v�^�񩧐�g
y!>�������m�xRፗ�Y��"e�K���ET�u��1g	�����͏x�֛��"T/;*.��+�5��^Rk�7\���aZ�ʰ�r}cJY�C?ʵ�|"��eC4�j�D)��e�7,�"�K�=�|c1��*��!�gz��i�S�� б��@;vG2���}u���1��5�y��g	���aA2%���8ڑ�T�m,)�x=A_��s�DU�!]��X=��m��	��A`2ڵ��_���C6���0���h�V\�Lm �w�^n]7)��ʷ��$&̊PT��ְ�
� I�>�c�<�@��NC_���lBk��]��T�]�vb����CD�ֺg9yQ�^\Q*̸��.m:�tRP���b��� [oL�Y�� T�����6�����$hs$��δ��GMp͉q��Q��1�������L�I����k� ~,������7��V%.�\�)�?{'E���+��!���^o�c���q:
9��T�	]<��\�=��=:��i�K��Ö���Pt/�?�̿���ޥ�S'�ۥ8x�uM[������_��X��G�hgј��w>C��S�S��U��u ���4z�*���R��c��5BQ�J,��|ď�X@��}��O�m�ZG�D?�x.�ƾ��J>�hu�C�6%n�!�ri}7�N���Z���\��pW���D�;�)=щȻ�k�<�P�$�.����b8��3�@��KXtBc��lV�\�
�b���l�,�e:*������i�Z�U&[�Ӛ-�󇕋d#U��=��rΜ���RH�	���@�mE�.��L��b㺉@��U���E�'�O|�3O�FKQi�Tx̒�c�U2���3��ܲj3�n�I5@|W���57|� }��G/��V�*�s�G�
4g�Ӈpo��NjU*�b���>L1��D�)��(�y���"p���c��"��v�w�������b��:D�g�>�ڏ+�ȥ�Bɱ"�����×(�3���*1���O�*�s�O��q��b�[l	/�S�� �X/���c�v�d�#/W��8	Y���f�s=��T��UG�"HDk�99ցb�ȯ���
��PP2)�ZD]#-CPVW��ʀ�u����h��[��0P��*Б٣�͍ޑ�B"Tp���P[D�9
a�r�֧��l^��`��y3u>z�|4�Q0��t��C�{P�X�m���+Cd���"�!�%�ؓ�S��15Sl��d̀��f�e'��]�>(����ƅ�L=~/�Lh�8����m��yŮêc|�R�ӕ�:�3�Js��Ĕ_�֭J?)7��6U%�~���&�i A��(C��m�'%}��>��X�᷏q.%�o��V����#b.�����S�4�Oq4R �ŮsSYW%r�W:�@���1��i�V��j���D�0XG�� 筗I|EZ����.�
Զx��M�@򆵣�������^�B�B��ӹ�`��7f92�QV�X�4�|�qo>k���P�� �y{� ���jb"�Mkkz�y������$٣>E�FJ�V���^���#��#L���lT�����ҭ!�{��)�n ��)$�߳7�;G�C�!<���I���f���-	�����"Df�`��*��:��P	X�+��1ZA�Ng�4�6�&U��r)w�u��*�/\Em&�r��&�/"H�Ӎ�e<����z�e~�
SzV|
�Ș�J��&쟎(�j�؜�W:W~���Ni@L�wױ�b�ˍ\���cЬ&O����Gc-�����`QX�۸��c��9Ӟ\�)��ͪ}�21Au��ۜAP�k�>!sy܌�~�"�[�NR�1a	��6���~�.�-WK�!M8>��̶�4V�9Xb�X��.�;�P�$���5�iZ��#�}�3��q��\f��1�'SS!�o�5���_?�]r�^\|VT]ё���I��[7�&er>�ɸcsqN�ƈ��A��ǹe8i.a28
�!>��S�4��3)�ދn��韧jPb\d�9�����$
�n�R�M�9A���x��� ^$vDҭ��ЄM$:Vs\�/ 4\̲o��r�y��K��(���7z.s�(G��Js���Dm��HM���&�E�T�U5�O�:�5�܁��K�l�ْ���n<P�'��z�i� �?�t�=�)��aX��E�����S�NP=]_W}_�;X���m��o6�$0-7��7r0\.G �21��^�8y��=��E;y%�*�Y��я�.A ח������������*�#7q���>i-b ��� 8���۬mV� (4��"��4���t�f�9��P�(r�{.@�SVoEm>G#�k#�X~���Z��*>Ku��u#��s�F9Á��~��ϵ<:Z��[����1�R�����:fsE ����+t�jJ��]����;l�I�� N$|r�gx�M4�<o�>H�ꛯޢh�C�CC��C�����O�Pd��B2砋�1�bi�
�)������p�B��u��?\��һs�;z[`Y��A.��w����쓉�V#U&d�~g_���s�d�;�=
!h��$�t�����X+X�U��wuP���
��1X���Nn�j������Њ,�[m]HM����V�3)q��TpI�]�<��3���3�E��]}Y�EX0!�R�!-N�=�4*����jx |4�` `kv�����bX;�I5��]U��"��O�3W��!Un�UJ�&�#��d�a���Z��.��Չ7=�̑�-˄�%J��xm�=T'�МϷ�E�2zZ�X��'�=L	iP���mx�"���%7����@�3�Bkgbt��6���Yc�5�L�𻺄o��[`��7�{sf*���;#��y n��W#��X܀�V�f�k��J�e���U�Mc�=6�7�ɕQ^�"���,�E��O��Y���(�����VS�
U�(8�t�*�RqW��V���j����"?�%���}&9�"1Rԙ���`��k}��v �.)F��"�b��X����?rQ��ջ �h��%����,��<��}�����T ���7-H��3ϭ�U&�^�O{����"S4#y=ab�(B��%��L=	2�x�YL,=	����8���!���0X�A��;�}���N�Lگ_�0	w?�VT�3�~w�_�?�a��H�f(�2������x�{��]�]���X~L�jQ�DS��J�-�;~�LP�a��TEf�*V%�.-��ԅ-�h�w��9��.?�;��h�ӳ68~o�4�'�bJEvD�i��X8UVG�Fb �)&�zO�%�!�	���E�g�lX���J�K��e
��+,=3T���q[���>�O��:��R�@\m��c���,�yA��wh��)�3����E��p���H�������5��y1����zZ�]�W��o���A5�U{�%�H���W�e�/k�]=y1sKK��8��uIF��m�("����V�Dt[7�ݓ�j�{�ݲ�}�=L�6��&�k݌�L���1Ą��F�U�3]ܝn�j�:�O?��m��ҥ�+�Pp����t�Q��~*�,i(�B{��&��~-$BQ�UNuw3���H��<���h�d�0���}�l+�|ꫛ=�:;ԏ��D�-�J�bL��n8h_�ز�
&Ni���c�5b����@�Y�+z-�u�Y���4��Ƥ[Y��2i_���d���m�J��)BO٧zܴ5X	F3_;��!ˎl�/?����f�\��N�]�Ucx�<c"_��ͮ-q[�5!c3��KH�����%p.�fda��?c�͚��S`���� h��hH�NSn�����2���IX�h�i�~�Y%�J5&���_}�Q���W��Q�J1ݔ����<r֞�y�αf0��֊@�HU����D�{~������_�e-�iZl���ؚN@r��oF"5ð0�K�r3_A�-[�a �j�l<h�@��hI1�)�w����>�~J�YIY:�5�.�R�R�_N��{~('W4i,���:Ng�M�����%à�C����}ެ<��?�;�� g2a���tP���\��]�� �H�q�G*rh�e
��x���#�{�ݦ�ĺ�@k�����CC���ʂcH����ǁ}�4=JA{)ɂ<�l�q�bw�:ô�\2���%uP�$�\���dns_��n9�#X.{�����^������*]!�T��ց}~��(�|]bS�������q��(eL4�nP�g�7=�*�,����i�{h��b��1�	uR���/R�M��kbw
�`��$�Ɛ��~O�{$�a ��@��� :̇X��5ΰ�5+�-�mw]b>�uq������䰶.d�J��q����h?��G#�#yr�Eî�l�Z>E��ƐTeYy�4�������}��F}��Gfs@�߹��zi_������9v;�3Y�o���T��[R��z�P'� ���T�k�u�V����Aփ�V��ӓ����:�I�q�OQ��^�ƺ�Eb���c�=B ���)ז�%E3�44��b�`\&V�:��$�,Ʌ��'�{��wjD���%�VP-L�OVF��W�(�`�ܖ��=ce¨'���~�����ef���<F�k� � ��+10K�m��N��d�F�L��k��JZ�tk�g���*��U2_����D�v�e���ĳ��sU�.���v(]e�nz"�PpM��u���~�6EK_Cr2��[$f�!�skR�����N�/z$K ��)����T��d �j����1w�-������xeoY��:8ñ��*@,C��ajZ!��r�:g|r����c������s���%�^�雅�t�M���Z�a�>�!��<��=�},�H#�l�H�la�3)�[���4"����Ƽ�������
q�݉a/��Տ5]<#ݘ����}�Jز���`��/j�#�Ѓ̗�tȥ[u|��Z��Or�N�����&�� b	���̫���	Ƌy5�9�w/�Ǖ3@���]'��2|��n4��i�C&<ò��F�z"��h'B��q�oY{�fh���00'�� �7L��&�h`trKҁړIy�3��w�T;;K�whR��8#�ؘ����ϊ;A���{�bW�)(�;?��b:��������"4��O��/�Eڊ�����;a�Q�[L.���l��c7�6�G�Lo��+���+>��0�iM���'0�Qu�������\E+�[���&��n���+�uX�	�`1d/P��������k��%rh)�L�6�+~���C��=m��z�D��	��`�-��i������ʹNm}q�������q��[�[�(�-�v�"Vj?�6���rΦ��s�Z�Uc|��,�H �&��r���@fd���a�j�י����4F�mޡ/յ7���xbcK��,5��=~����F_��\%�9\]�5s�ṾG��5N� ]��c'sA[���4
��dԕF��e��&+�x��H���-&�)�1�7�u�f�=�|e��2y�lZ���~���Æ��R��*���Zzh�� -դ���j���K��͝����v����Tr����Ù��){T�I���	ZLؗ������c�۷�ܱa��طN��s���~�i����$�7���i��ڔ�	�]�]��L�&���M�����S�рm�.�`m�5Ul�(����ld��ў6�(��R5q��'���GZ�{����b���*�rJ��܏Z�reX����5B�(Zs!T�]�ػb�=����.�q1��?�n��<�`���x3�Y��&��э��`�=]8�f�+�ݬ��N�9�'����O>���AwXm�u���������j�j���b�I@�Q��7��o��Ը�Q�~ʟ�y�%?7�~&6B<��!J9��$@c��{��Y~BZ��dß���^x�S������ɼ��j-Hf�ը�k�#U3�Q�
�Q\���9�q�y3)ס	=t�ʰ�&�jL7���(�6H�w*34q�y�-c���W퇇��;6��z=!<�/�;DI
*��q�$�Q���3O%�a9#.\��s������[(���^Mb����郖I��,xt����*3�өb�5T��	���G��}�ـ�xaoxn8�w�~*��oj���D<?��������T��:���TP�'WE1�H+N1��V�q���C0�o�,���2;�"������m���y��9�g�1��}w{��Lo�}	��ඒ|�giW &�	�93�#��F3t
.��"���Dd?J�q(]Z���y�.ES�Ғ�ӁL>�H׫[����Н�.N�xL�G��V���/��5g�o�D��N�"�k��w�EX�I�;�Ak'�*}�JD#���y8T�ԑ�z����ؑ'�CzH��
��R�m��
��-ۿ���kk]`|}�v�l�i�7r�!�mR�i����@���Öz}td��`��4$����v5�-�Լ^1�eK��hr��jW?EhK��$ϊ�V����żᐈPz'�C�7���;�����V��9c0°��x�e�E�W��xw��yQ�ٿ�6�6�7�m��G�W�m��p�Or@�!җ7V�mv�!}L���Lr)5K��.r-;��\�<`�v[:����>-W$$����VE�y�<�^' ���1�>�V���	�;��E����� �KMG`}�7��<�ز2Q�����P��~ν������:��}Id�˜m��\M�ی3㎩Q��S�!���,�+�M���YD������Wh�!h����+�+��q��}b��=_ ��m�y�0�Wd�� >����<[8���e:�8WB���Uqy��~���0���r��rYG��v�Hڷuu�H���n�d�x�g��b{��;%�u�?�_գ�9:��)�S7��5�9-ѫ\��V���4�3�Z(�-#�]C�	��_���`�)TY5yD��t��` �%�k|稜,{x�r�0&� �/{���wO�����lW#[�伴��Xzw�,���a7v�pY{hO�.�uG"Ʉ�`��^qX�3��<d?�{�Ec�r\ 	�;Li-���׋9�g��P��[[����f����R�I�+w �aP���q�����a��)֐����;��˄��e�����4Cu��w��Z�p�f��|�`�)�1t@K9��# ��vu1��\��ǵXv��,a���m��?�0ؼ�p�$������HW�g���Ոk-��+ɾ������ۘ$r+U�A5l���kN�,(��SpW����*a\Q&�/s%�q�9f'�S�׷�٠���`G�������r�]��ql�=-w5>��#�P�U��`D9{��u.�W�V¾��-_l�`DT�c�_i�̗��ݳ����P�e�D�D�u�e+|;3� ��P=��f,`x�8r����vK�� ����Yy�MZa��qE�>5巑ƾ�|�*���h�2�[E ~@���3����챜�9ӋV��Z�Õ3�w]<�X΀n�����dRn�Gl����Ű��6}�Fg�7��Q�+�Y���}��v�;��l��a����(��>�E$\��ӆss.nFx.|�קN�m�X�>���,!��9�o}j>����*����������fS�њ8E���{��H�PdLIH���Go]L,v�2�|��� ������l&������c �u
�>8sZ�q�f�� ��#>@����v=�Ӓ:T�
s�,��.��U��X�ao»u����y��:wJ�潗����4(A �ZY6�xi�܎|��]�bG�苀[��#f���-�uϧ.�'d�8Q��햫�ê�#���u���ud���d�0�f|iF�-�g��p�+"�Ҋ1/�8��F���fk��ߪ>1U
�c�
�%�'|��D#e۳���
(yX�x�Rr�;z���;xb;���'�7t�lpkS�����Q2��*�CnHɜz�8�X7�ɢ��~E���������gLE�;�c[��5�CX�=�;O2�[1A�5�a�-w�|ʇa�e�=�]j��� ��"��At'�s�uY���`�(��ң_��`�pk��6��]��~m�m�C�~���bޓY%�h���2(�E���#-"
Kٞ�\�R$ޔ7������?���=g��BJ���_^�!�SO�Q_�N�UlW�����P2A�ۉ�6�걁u�c�<��!�p�I�33%�3F��6| �	�h���!��C/�hO����#�=Ʀ�`.(�U�j�CA�	Y@ �tc�"��,>�qQ�;���z�3ڕ��H��?2�
1�+��aѽ�ޗ�������ľ��QԪ���ao���G�@�����x�\�4p�6��Z�g�[�������'�ĩfn���4`$MUMi�1]�gCd�-�n��I��һgb��H::{Ԗ�_��%�;j��݁�ʵ���Y�����h������tE���8����tu��N�x�e�&쏙}U�+�1��r2������'��纊rg,\6`�B�t�M9�q�� ������j��7w���i`�i��{��3@Z��^����S³a=~0��8C�TG0)H�k� ��Ͱjá��UX��)�6	�Ӌ�ҋ��ɂF�vGIiPLhZ�����{2���!�jA�Z�U�=A�5�)���N!�n�)�RᏂJ���	��b�s&�m��������f��KJFLkƸ�s����e'7e�KRϒh	7���}�ʗ��І�����=�����kB�P�)쳚��ogL���o��hL�!w|�!��՛��⛪9���+�6t=K��b�68�m�3��\���?��K�2�,'�#��Sm�ޖ�g��滴��=� �1���|:��ܛXTA<[k����T&eu!nu����I�ů�:��Rا+����
�?&��!tãy"�u�XQ���SO��Ÿ�醘"�CDw���1������nrƂ��h��l��!���?U���7�E.��ѐ$��Y��"~8��B�����s�H�_��/>�s�$����a�"C�n�3����I<�M��2�rGHJ�e_T�f������9q�ʢ){���Ɉ�v}\X��K�����~�� ����	*<���lX$��MYf��G��{�T>�HZ����4G~�� ��K��<a(������v�	{@�i�i��h���J&
��4C ��;���T<�u,�?�M�ڪ�x����� �t��V+�|�m��t�n�1�Tj&h����%9�RzR�q�=��f��u�|���6�;E:ҹ�o�с�E�A����X����<�1#Λ�қ)�^��S(�4��s����։
����}���9t�jI$��s����C`� ��Q�q�^�YS����y@�,>�3ReU�����`�M%�����;�:V�:��`;�����#�����תl��AG�97n��đ�B�ͥ�$�̬ͥ������X�a�r��pԈ)}��q�rX�(s��2c�>��8��K	�y��k1��kZ`�b��B�n��_u�)|��+dn	,�M�Ǻ��i�@��K�3}j`���rw�q�ۗR�smlk�Pmԇ`4pC�М[�i:;���KG$}ސ�{vw���|�,%�,8
x��\��)��V׆nN�DnT�����Ok���!�RN�9��{��1`	�X�4 �9�R��QBʇ�1�E�Cti������IQ�L%\Cϳ��8�P('ʖ�V��&M�f$�ߟ�t�h�����A�!-{r]���vKz�8��i����3a�)�����O	a�3-���>fMOH�v�~�H�T�������-�I l�hO��4K�@-޼��|��С|���_��ZQ�
���!=E�����N��ɷ�w`%����At<���Jp�,���6�;����\�v�w���Eqg o�nX��{(�=�B�;N�Z�a�=2�.��D[�BC��C�i��\_R���Ҕ`��x���3A��/�8 |�<&�M� q�]�G��%F/����TԦʜ�U5m�=~�U/��L��d}��U�6Z7g['�n:t}b\s�WJ�o~�#�y�/k~Fj�Xj�T	}Κ{������BY�Z+��Lt>.��W�>L�2U��`<��0}D]�q���p&@o0�W��~]R��"���/5lS�&��"�T����Y��Ѩ���Gzb��P��4��j��Wr��r�A�}[RAu�GX�ݯ��D�I�NoY~_�eo ����qt�AF=ɡǺ�`)����'^:�L���O��H�@�:�;*<�0���!&ʚ�/qǻ����#M���&��F]d9��u�=���\��p_^Q�%�4b�*��EƦMi|�#1��Ku�`\�xr�&��~�\=���`@ Z�Y��c�8a�ѥ6RLXݯp�?�@~��k"�+�Ѧ���[&��c[S.D��w��=X�&�1�7m�źN�jXN/$1~/ѳ��~Vg����v�|2ո��V��t�sk3�Zt�ãr�S�o��ø�ۗ	+E��>X�-�"����t�A��;���T�������N�0�����-�װ�T,���1 ~����Y�\���mJ�2:EHPWb ��jr�dG"���2��"��9��gƤ�}�h�(	�ڈ�����ш�&�����@�����w�7%�_y0���7\ݧA���ы����ð�k.��%�c�Y�M���cx�
�轒?�vGM�ߙ.�I
'8RgX��#��^M��j�پ9�)�1����Ư�D_k(�u�h�B�	d�E��#��1�w�V�!����L ���!�,�y��b�9fS`��I��g
G�V�c6�\�D �<�T棩��~|�ÝO=�v'?�9��7J�,�� �{�oU@%J6b�me#K�E
�>-�k*R�{%&Q�wVkc��3�"�/�����y�T�a�o�#��S�B�ud�_$��K����i^��o��4P��nYa�m)�WjgA��c���i�|��f�X��g�Q�n	HA��Z�D�a�Y!�B#��Z��(��^z7�s��s��H�rH`�2�]m[ǞG k�C��[����f��cOiWt���?��,NQU6�Im)�8"? a��-X��ZU>����`X̴2��6� ��@���R��{L�3_=h���@3]#����KQ+�=��m�K�)H�����\Zh�DC�+nҜ�ڸ��ƸW�3&�PEѴ�&���eτw -t�Z��v�f�K&�p>>�h�d�L�-28��w$ϼ�k�?C%Y���۵	\uEeiQ��[2�F��Zd���R���uZt����x�M�+*��n{�*
�G����.�K����~�*����>��������_��O1�a��ZS�^4�WP�������Zl����ErG�g�z����b���D֔��֤ �Uc���dx$���<��=�&�iơQ}��q���k&K�����\v���|��dԣȺ��ǟ��<��rfͨΙ���4tLXy�F]��	Q�������*vS1�bv���a{K�s6���ߨ��U}�A�k��(���c�r��b/'�20��=~�����
�`RIϑQ��B⁔�%D3�`�+-Y��S1п��Z�'�}�l[���Jpoi���	�u0��Cĳc��J8�`�x��Px��l
��|ސ�Җ46����7��L���c�(�l�1���R�.D5<�%	;�(�,t�U�x#%%���F�2�h�%d�LT�L�������I���d����Gh`-=�9�_�h�JU@�&��7�R�j:��ȇ�o���
*t�������&����:�b���s�΂��~
֥�p������<aպ{��Ph	�H<��ب.�ذ�����,����>�yۧ*��IX<d�`�G�>�u��R���dX�q <��lw��g[qϖ(�c~lys(���/���A�\��+���4��O�?@��A�"!��f��ɹW?i���d�w�i̭#n0"_X�jF�����}H�v������B/#s@�\R�:��,*����P�f�������{��L Ǆo��XI���*���);_�J���Mk����9(�uּ3�x�[�LQ�C �|�R7��;�:d�P�������ڞ��E�c
�>�٧	Sg~ޑβ�|��Ih�h��> 7�Y��w`^���/"-ktv���z�\�Q��Ʋ��3��{s^<��2�u��\�֞qQ�y|S��Y^��'�e���W�C�gk���0o�bϛ�Nyj)�J�,^�-ة�G�`#�V�.t��7"����O���8x)\�o�toAR����[��}�_M?�qҽ!�����
�-���r}v}K�����?�$��F�Ǜ�����eW��-��V';+�:
,AU�d�fg�����A�1=�j��K�*�_L�BB���$o���X�{ָ���2�r�Xó��q�Vε�8�_��q �ɻ}� ,Y]�nf.g�CW�D�@����~�p�b������7���i���.�����=n�F�P�*�0ͥs
�hf�}�_�$��I�S�X-*�w�]k���n�V��(��a����ȯ��Ϲ!�t�_G�	�	�o�ŜF��P_��-ZW�C<���j��±�i�n��E:z�%������A�+���*t-h���:���uY�z�o�®v�U8��U���v3�����fH2��AQ��1\��UC!���U���!����ɂ��}`T�CM�Z L~��;��4��xAq8��i|[`�J�.��?�`�80��hBON��/U
����-b����+w�����}Љ�W�n�nC�Ed�y�{�5p;Zz��aA`Y�Ah��T�U�l��\�w�|�,�옼2�~�֝SG��W�oۛ�K'�OğmptbBÐJ�[)�֫���<�NC�Q�z�f-߲Z�3���`���S��2еs�6�u��9�W-�ݳ����*-S>���9/��om����������ڤǸ3�Ǯ����2�c����UF�o+5�2����j�Y|��|��hCg{��'� }*#?��,��610}�UR�U�"�¥�V�SL�A�k��~�%��0.���:ǡ�ia�wkio�/dH!�>�ϴų�sʁ�Ň�!n���vYRP���50�x�����ڗR�L�����+y%|��b�u�(��Ū�%������
��+Y4�����y�3�dI��bD��E�����1V��܌�p�-��v��׬_|���?�㫺��x�,��>��u�s�a�=�/)��{��Ǆ�iڌ&�A�X�}��j�F��L�2�B�R�I4e���s0��!�,	N�`}$����B[��O\�J\f���������f��I��n� �:�w&k�@L��lY}u����~��xviQ��m�@��f��J#W:�Q0�E��7���-�B~7�g����
3O���{ڜx�5��4!qydyXѡd?��cL�4��Oе|��"�)x����vN濕�t�Vy$jٷ6.^^��U��B�1�g� �z���$�0����lG�-=������-�A���9�`m��$�<��#�=�B�\T�U��,3m�̙����~����x٦y�뙯Cc$ǡ��7^~6�����5��c�}���b�u������F�>���\LT�����aD�
�.�O�eh1�.������,"��������ׇF#D�9y�}T����\�9����-�>v��0*��\> +z4��َ�(��G{�����VCS�B#����N�ra]#���)�������ݒ1�����+�SnvW��"�*�h�z�ɛ����U�qwz�0�he�&Nq���TS»�TEpǧ�8Q���h�|���I�:�UU
u�+۠n��bN97����-�>����C�}�i1�6d�Jv��H�TR���tK���:���w�N�*9Nĳ�ˏ�K�ч^�ϡO�[�
��*�"_����q5:H��w�����qZ�ƤvC�G��"�iu�4�B��#
��6�~H��t��[q9����F�P�O�_�=��;�jT���V�倹�u�c��-7�?����d`�
HKIiH%S(���Ĩ��æ��"M�_���!�!�YD��T�	�<�@zo�����i\5��������J.�0&j���
��WP�X�_�s��2.c�й�~:��6�#�g@O���~RUEt��	�h��b�,�\R��}��|���d@���}䂓`(�w�a
���1e)��� ¶���E6���wf��@	�Ñ�ZZ6�d\`�h����6�M���h�6�7((�au�i�����̣Mt�G��&@i��Ư�������1Ev��^NM<*���I>����-Y�y��Q'V���H�~|��E�M��5Q�ú"���ثӆ͚;F 2��S�*iF��Av���]�(���`Y��ꂖ{i.��V�\�$�y?��L �r��3��K��MX��!�ՠ�6^ ��(5��(�������x�ȵ>�;(.��
ͅ��"[�'��������h��常=�2S4ʾ^0�;u#�tY�2!A`�NU�V�(a��\u��F�euv�k}pŇ?qkب`D��(,!�vp%V S(|˼a�����<܅$}�5��r�%��y����h�p�\���L����oB-��-��$c��zz���ܷ}�,�ox�����a	"l����T��j$fh𮶎r�B�ufh�d�0M�������+`�":�Q��ۯk}�L�u�
�݂U�iJuUz~�u����v���lL:��E�V��rIഔ<�@�ayr��D�Ĳ�"�9�a�4q����X�p>����-X5}�ۣ\�l��C�#U���tO�bZ>V��oNד�1~jK/럡�['�e�����Fx���Kp�N��L@D"TjAt+����������'�F��F���̪�����s�O
���ʜ�$�?n�K�{����E�ÝF�?ǔR�K]�IV���V��: M[�X{��>_R����\�3*yR�2�jH�w4���a��u����ُ��F$pY�m��/� ��~��%i"���� U�o��,�i�+>c�!����]씞I®e��ա��.X4a�BS� Q$����4�z�`�]�B�������]�=*`)72s�v�|@'���0�����Dmm滙]����2<�l�����V��P��B{��Fw"�~S������0�O3~�Iwa~�~��� ���?f��~��� �s�I�}���s��@2Ɋ$�Rf����`�����ƦB���`�ts��k6�2@q�\��0S���Y�X�M(��nG���x!ǔ��t/4SÜ1�P��/5��ڃq
�����;QP�J�o	�q�>���BkbM��ԃ����� x������y����6��LZ�j��S>�O�*g��t�I�xՏ����.{�������!#w�1Z��Ġ�W����0U�����$$3�����[���;���Hz��A�b`���������v,j"Y>
���j�VFKY�Ɏ�|���6��ʮٌ���o�G&^�2h�k������^'m�������M�3�:��Й�"�6������VX�@��AXR��)(anZ6�GHR�)]�_�hKOi�Pd!oDF��	�}��P�yd�_v�/������/\7��7#�,A7����<f��n|�p^�'/�	�"ٺ��_�A�r�
���}�I��A�,��s3�j(7L�4�B8p�8���_&�� Al����C�[Y��2vh�+���ǶV2��I�b�b'7OxGajNW�`Q���� �8_T���TU+�8�3�̈��t������4�5/�@�Z�B~@<�۫!�P��V� }�D�|q�4m;nH#NYT��#��#J�c��̗�4
�=�r��
�|)��N���\����}9�G �Oa��v�wyi��I�TP	�6�Z �{���eBAj4)h�s��%�qag8�S ���55���{�5%P��� �"�NJ[���c����pÚ���;Y4�ڞ��m�97���#���cx%�>Ǫ�/DV�b�nĠ�dP'@��'e�ϊ�#�G0�������?d��0ED9��qW�ͥEQ)�}Zw��o\�<�'�b+��&�iY�:�:��E��-�GY=�0Ymo2d�n�|ji� r"��e�c����:��u6�&�s{������߱����z
͸�{	 �m�iYh���6��n���3��Pc=�\���\���Ė�O/c����p̛�1P���$>�;��+����͟���h�l��[�5Y�����Iy��9X&� ��i)�%�W�L�"���J
>}��M{����Y{*�{2��5`������+�8
cl�	Cny�i�7*�
�HL�}.+)|�T��\D�E��28�4Hr�J0��2L�G�T�+�7U�e1쁬|R�M&�/�ý�+]���$��{�g�|٢t+3o�3檳�㽋}V����×�T����Yp|FQ��PW�ӱ{=��l�T����c.�,�ٶ���=@��Y�ؘ����p���۳K�^�9ϴš�����|�hh�KD�+{�
}$V,,t��淳��?�/_��w�X�)ܞ�<�3X��l��^�-���_����j5�sB�j��҇��:���s��O��g^Zp�
�AXN��9G(��b����?l�P"���{SѦ�fV�.����p/H�rt&�f:��O	:ҫ�!)��֮z���6���i�&��N������q��c����%�����6��7�!�\�?�������Fw��η�}�0��-`)�R#t=���'rU�/xӫ��T�=�H��1��ٕR,��� Dm��-4vF:g<���Q��{�熣�p`�����Tb<O)��=H9Y6"��}�cD�p���F"T�1�90/$K���E~�3���<R��3G��Ǣ���-yN�*��%���+��,x���Wu����p6��e9��`�Yq�	�?�j=����'�=
�æ�6�ц��*$��'Cq���
wϒ�� 
��R�N����cR\�(�e.��樀�]
��Qb�y�@P"�b�.��t~A�&u	�.X�-Ȣ�r�й9N,ֆ�ɉ��}��ڒ�����B?in]��ҡgQ���c4�ݜ��`��qp�����nL�=�4��ʶ�sa�i���ay`K�&@'~�?���=�o�s�;
/����
�x��E'֡%ٟ��)��8'ӏ.5��@�V���=� "��8�ěi�қ��~c��:x��S9�	�w#���[�`5���Y�)�5!eiրl(���~֔��	ژ��T+�p�=�g����yd�`�*V�S>����to��l��/�M��h���q#�A沑���M�i���u�D��	��i�p���ȓ�F+/�4ݱy��{�%���4�V�e��Y�3�����d��9|�r���Z�{�%�gV���>�[�]�,��NQ�lx�����ڦ�9V�M���w=��I�&�p����{f�T�咉�XV�ԙ.y��� Om��i��j��,�ͬ����ܝlN�m�tmgw�E/5�M��X8i�:v��
��w�%:�\�#
{�v�/eo&�x��J��j�9�Lm�:�E�EX���Or�_	�S�)a�<�0�z�Q��uwa%S�
�%�Ƀ��߹fwg��0�@/�o���<�FЬ�槈�%ط�4���S��;?[�����Q��E���P�b!�,�<�{8���q��y�y���=��$�蹇�x���3��ʓ/�8���!"�I��/��%(�#�DMpW�91 RC޿u�����K�SL����}ZƂ����f�,1,�%��/p�s���Z�<�V&.�������d%S6g��H�]߿��e��Z֡S���X8�0ݹ��\�*0{��0��U�W����a8�j�@�av��ĩ�:6t!��JAn�D�n����j��Sblսhb����3SUUH4TAjn4,�)���ŗ�X*S���ɪ2c"�`=�p���,ߑ7��tMw+�ɍ��F5|m��Ĕ1$�%7����m���_I��˂Uw�Y爨��}Кf�
)v��嬌Y�M	-�=ղ����ݫ�x�`7��,�v��~K63�Bp����*0uQg��Qm���!�:�?Џ!U���$I{��[�HY2�\5��ns0�B!M��E�:Ԓ[XTo:�Ҿ���Sq�Н҉��ᑀ���
|��8Y�0�����ݶ.�Pw�~�ru���%���/WV����L��
� ���S@��@493�c�V.��BS�'P��缆OՐQ��y%�^�� ��p���;��4kZm����'�]
1��񉾄��\0*U���?�r�y�}yb�!O��a&yE̿|º_Xd%[ǋ�5��.O����b&j;R25m��۩Y�;�Z����;��G �ŽJ�)h���c���M�,t'�i(������"��㓿:X�U��0�O��SX�[_mz��e���9[@�kh��:�Ԟ����ġ���)�V3JXgX�-b��.���>�C(�e�Bt��'���YJ��DK>o���T;����z
�Q�<=���ѣ���y&�Q�N a�0(�C����+Mͷ`%(�gu2���#��T������ `2.�C�nw�a��+łqk�D�9�J��.O�3��2P_��4BmF�f�s�=�FD 3��L�KҘ{�5^n��o|�È�+
��o�\�c�*ߙ?t0�%�o���</c5A���uƯ����D����ǟV@I�w�^ �S�%/!��Y��&�}�h�$��72����΁����+��
7�ߏ�E�0}Os뭶&���\�?#
�c�L�cl��Ƒ����H}���lU7,�:��2Z1�����Hp<yOal�*�+�BqC�+ܦ��]>�f��f�# R���i�3(a�J��yR�����~e
�2y6�\"��H ��\>Ibz��fb�-c�W6�R�6��BI"���K͕3˻u�3c�գ�g���Pe�~0��������..�	�6��#�ϩ����O$���CR8�S!3�L�[Qn�]!)L�->(�7֎�4ܕ�ͽ\������I�^��b�.
�<��+���c���u;��1��5�2��[�YF��b��Q��7����z�"�-w���8�#Yn�w8D�3O����3�Xs���G{[�{P��CB�zq�K�ﲪ3�ܑ������\x4��ئ�k�f���k�H�2��՜���<��(�ė0mI$@
����K=P���^��(b����kD�?�c@�I�|�1r���LcN�D�H�3�i��&�ƪ��1PV D�Nnm~����W57�b�!BP�a�&�rul3*x���L �X��h�ۿ~K߷��������V�y{�c�qO/��SC%"��#�C@�I�{o����SW7�aɆ��E���wb�]vz���S���}v+�Z��Q�}!���	G�͑�7/g2��NP�	��BpU֗4Ƅ^lX��>� �|�����ۑ� Y?9�Lmg���<�dpLJ޻���t�@�n�A>�_)/���ު���km͛v����4�g��z^�!�*v6��8�� C�X�n�cA%N��Ãe(�C��g6Y��8��je�r\�D���+�y�/������cud�ǥ`�f�RFg��:؛�?�!����퓲�2�Ҽ��l��GP;@��OO���N�NO�;$�I#'�B������Ʒ������UI�P��
�]sw�v�x�i�.����)<_���XR�}"j��?dAF/#��]�Ԓ����Qt����>_������	���g����-U9�sh�~��]�`1��Vr��H�}Ӑ�����nx�_�	�Z�4ѿ���6lj�^�3��v�~Qy��>�;\;'�����]�EP��<}�u��=�@�WKN���5��S�~�|A��n�ӔgK!�/�K��u�?|
��Z����6��a��9^nĥHT�¹sw���� ��)V�/�{8�;(��}�U�Ѫ�	a �����J�r��T:r
ZU��`
F�7;Ht|��S8�Z�j�-%|����P�ST���	��j�x�n�J?@�J!�	?e�{3H�	!�ZU�����,��<���mn 5���t-���l�&�<|;�ζa�5�-mVR�~��tW�V�f��r�"�V�{��wX"�J-4���BS-f0����e�Q㥐�%�C�T����5�ZШ�����kC���c���d"��`��N@���LT����E�x�4�:`�h����g%I=��Ej�Ӊq\�&!(͔YB��o�^��izI��&E�*w!G�5�8	����-�9���|�����r�A�dX��n��W�+�'{���U�H�nE �硏U�����������3�輝KEڰM)�����XFUs��,�VN��&�Yp����*fL$j;,�2pr�X~���n�`�����L�$c��өv������>���+w���h[��W�\�����Z��p������shw�C��B�[���X,�]Y��}���F�������J��1n�3~�t�������^�Kǚu�~�bQ�1���`�02G�|�E=Mۊ�3`�杯��v��>u��7-]g�}�Jk3��\v��~��&��ED��<m���`�6G����8̽�YT)4|��~�3����#x�p������b����liy�ގ�ǭ�vHzGoN�0�:�=C��_�M��_A�1���:9P}9H���G�'ߙ�0�jY ,��Uo1ي�$5����+�ϰ4;����0�Cf�lwp(����Q}sz�Y	���l�����
�z���@��Vf���$�l���^Spl$���
�d{������P����=�YV�s��]��CS"�j_��?y�4��2�� ���D��$!y-w=*�h����$��
;��
�L�w~��x�-�[^8���->�8�����'!�5�hK^��m���Bs)��,�
��f��A��kd��mU�x;��X&���1'�`���f�	Gt��-)+�zZa��I��������"�C�]�|B[��-��������<\���L��Ig��V�~?f�v��@�J�\�h?H����O�J��g��K׮{�tK�7�}�i(��~}}����ݬu����ќt�IUn%�4f��WI�������CfI0�f��� y/|�����:=<J�tußd;��\J�.�F���݂�;Z��G�x��5�m�7 ���>����e������A$��:�Ɵ��O��"T��@��uؘ��a��#�5��[�]5�(�&a���G�|;��nR,��$�=��j]���
�a������Q�{�{|cѺS}����I��'��FX︣���߇W|b!mS)]�ɤ�����Y?	��_s��$���*��E������3�阏@����g�ܩ���ϼX�髍�k��z0��^ж �����J`i��(���"c)e���Y�4�f;�׉�>����c�_cW6�C[�Kȧ�p��̤�e6�� �*=���1��:�
*T@��_���,��tT��Fy�!y�i��g���YgQԕ���>j�^|��<ӛ��P��U.�Ӊ�Ja��މ�OPP��1�}M��g�k0��̈�K}�S�cY�ڍ�U�BN[������ �=�gR]'�E&$�B���WI���O��S�����)C�t=N�/$���0\$���|r�:�'�T}�E��"�J��z
4��x���ܲ~0"BVp�ð�+��T��2���G���<�Os=��&�C:�-ˣ\n�\!Mlv���1U{�|H�<^����t��?�@14$�C��>�2z�-�J(s�*�ﺜ�b�iR���)�<d���T�Zǿ���u�[C�c� nn@��P��_݆Ժ�C@��b5��O��u<:�t��~L6S ���j���=��d���r�����}˳�d�LŇ���B:�nj�o,��kY%��R�9g A���gJ�p,�7��.rG ��()ʖ
�Ƙ[�k�;9�h̎ۄ�����h��jrBL���A?���[(�����4/����_# ����X&#p&�d�u14bi�>f���Fy0�-��H��1�5�.�����~�JD��ۍ��c���N���e���P�J2�6�O���S�HpK��^"=�K�Q#��O��3w�X�=l���'Llꂻ�.U�}��M�D6��q��L͏�hč���S�v#�����IN�c����MKu�D:��H;u��&SHj��e���D\X��,���1(p��NPjL���a����"馾�@g�[���х����N ��sv�FMyK���x�P2�c�Js:�z�Gѯ�o�����l�EK��G�L�,qwg�-�a)%G��7��սt�q[�YN��O�D��x�#�N`��������k��
ٝ �(�z���v�a��:�p�����& Q��z ¶D�/�y�ǎ/���O�b|c�$���V��� ��ĭC��*QG_H3gP"z��;\&����NvsY�XX�yס&���1Gw	� P���s911�{7XD��Vb:��
�H8�?
W+̧�t��{ZK��o�T�v��I}T�>�^Oy�f��
(�d�T��O�3z(�{��Z)-�XB{��8^'�d���zG�2�����]h��_CV&��~=g���r�U���PҔR$%g�4f E��@�p\��C��aSv�!>�a{|dyAN��/�d�tY���rQ���Ļ�n�ڟ�@�+fv����hx��ť�������� }dy�6�4�����.,p��߭�������}.�f�s��	Jfl�)7&��9������>�9����w��)
C��,�EOiT�|�s��V>0�j6�K�cG	�����ϡ�h76b�y�d/�>|'ֆ�G��UF\�M7!����7{ߌg�!�[�.%���ȡum�7l$�>��
�F`#�����焋����;�
���fυ�W��2i�U-��_���F)�刊!G��B�X�_�@)X*@b�-�����'p*���[eN��W�o��~�f�Q�F�B� %cw��L���u`$���ܨ�$T$aؠ��,xw�>i����[�na�9��,n�3�,��V�f6SM�1J�[-�[�����MB�����ɘ� ��	�>2NB�Zex���o�Ɵ��=��G(�$��`��T����nz@��%���2s�W��OG��4�S��'�Y6���� 0)���;+L�dQ���sᶩɗ�0`�$n�zԖ�/�%�hF�9 ���Y	�E����%w�e���W�񿦋	L��Z׭֬�6RͧO��Ӎh����G��O&~f�y�����YT�8�˧[�(b~�!�������J�Q��5Pn`O-�Nl�4��Wx�d���� ��>V�k���<e��U���"���;��Lh���N;�Ґ,�n OE
�����=4���k����<�K�z���Xr]���,�GV3�Y�2.$x�)����m�1�`K��M6 qb�� Kr��{�&
��~-o�>�
��Apr\�a(�^�VS%<$�e��~{s$4���e����̶��q���;`���Lnoq�^� �=��x�4p�\S6nL��ߢ��foP�Y��^��pN�1��:��@�NGhA鱚�ea���nƖ�S9}V���2�>f-Q�&3��v�2�ك(�Z �by;��d�/�ی�9�Ь�r����L�L�����Y��C��'��e�x|B��$"~���ܜ�3�:m��6�vE��>��ɟ��t�0O7a�ʞǸKf�g2�[��K��M����,bU*m%�%0]\	�O��Bg�%�`ٱf����r"��X���?Wa,��o���.�ۅ�tam�-�˔���</��C�M"�+qԬ��u�p�/-��-��	��Uhږ�Ao-�0~��Տ��9���>1g��bP�����4q����c��`����+9[������/G�'�шg�U�t�ٷ���G2��X�����v��1:�7l"�C*r0yф��.��m�ȶ�
xH�3�>���VCW�Y�pZ����oxV)Z^�\��]��>*F;vz�;�M$v�fT_�
��G�����D�IZH�UMp>�]$/�58��b��+����n��������
r+��qm&,-��!������	�Aic������;�C�S�kc�X `�7M��J�P4���|\u��N�\����УW/�d`��P���m3NAiF�ߊu�L�1��h�ߡ��t�OK�n�ϋ��fcdo^��ȭ�7�4z�'���R{RW2<����9x�B�.R�h
����8�d�BC�p�!����B\&²�{����[��?}�塦*DGqX�4���v��"sW�2�����y���;��"����{1&s@��:o�o,�^/�q?p�s8Ů_k���	�<UL�^��s�`������/�)K��gxu�C�.�M=��q�*X�������ݮ@q��, &Ky�Wjǟ�W�ɖ�_r7,z��ۢ"��N��R��[�;D���c�VA�XD���N*ג��|�e�,�S�X�'��NֲiO;%t�
Q���7�{�t��
0���3���\@M`_^�ը�KEx�ײ+L͖�4[V-W ��r�}���=�\p��ΡY�F�qO���l�$��B�a�=ƣ^ۆ�l�9(
H��}5�ZUJ�<	+Dy�E�݅�����7�|i�.|����8AW�҆�l(��	��0c�_K��V8��.�Ը9�c=�i������/�K�lj0��e�#F7z�dq[�3�[q�`�"��1�o`�8���yz}
皆�,a�}����eN���sZ����i��r�Y�1���&;��wL��v!��Bl�w�t�G��`��/aҥ�E�G5�xTʭ�D�� W��`��2'V)ق)4��?�|���ۋ�"�bo5K���%@��<f�Ň�c1�mm�� �����3x���:+�\���Ծ8?ԟh*����AR�{� �­q��Z��
�(�O��W��O%��ءZ���6�(}Kk
���)	''�i�/dV/�{/��>=��#����G���G�1BP�B��O�	�X�xt���*Y" ���A�f&���R��r.&���?4�!?�e�(��V]�?`Gz+'���\@ S��<��@R6��D�қ�`p�y�h��M�iѣx���댺�{��[̉)�c+��Z�},�����[L����؞ɯRI;��~�2�Y�;E� �+��!�����r����ɂy<T�Fh%ĺ�w>i��d�W��d$m�7�x࡜!�g����{����U����I���s&~V;I����E�'�������6��	U�YJ���zb��I �R�E*��֚��7A#G��V<ֹyFQ�8� �"P!c%�ci��ԩ�@�]�������^fSO��T�%A���o��cX���l�`���vۖV���7��5�o�7r���C�]�w+�xz[��K�ݹ�IQ�eˋe��`����jx%c�f �p&lb���<6F�fJ:�&ǅ}a�W�lUL5��&�
k��/�-m�3�	�1;��&S��FQ5�d��D��A�焿l?�����.��c`��'k�Ń��m�d�8Ѽ��`96%IXϨEW'F&.GZ⡰n�&��PU��6a�>�^Q5�N��c8PLuR:�Pw�j2���i=#����Lb��Z��yn�Г�a ��M ��9�NX����M=�@e<FGĺA�T���Q�Y�ь��ߟy�4�c.r��S�Z���-�f�B��oǌ��O��bSb�y�e�!��pl��m9
�1�7۽c۫�������[�8������p�(�X�%�;mS*`�ݺ����3���1��p�f�ܷ,=8ƿ;g����Rl02����~iE���%������Gm�%��G5(�C�4���ނ@����Q�W��@�m�@��� ��P����n���j�����.❾�2xw��Й���6�'mjl�G���لa��6��0��/:����e�Iu��g�U�t�#�e6識�[�u�C����,姖!-ot�� ��y'`��QŖ����B���C��y`	���D�����u8X�L���-�VoO�Zl}Բ��g���U٦��βn𮟝�P��*�+Dߟ�s-k�$U8��¾on�]���丷���Y.�hۗ=0=��o��*~����~u:#! �wL�����
_��.�^�x߳V7�����f>:�����8�X�B�=bL��V����4A���s��>��1�\N�풟q�E�
vc�+(����#ĦGɢ�@b���"���Y���o=��!n��	81=�������}��>O穲ה\v�,fOg�TH�w�Z�UF�2}���OJ���t�]�u������wy�9��y��ҵL������ݴ+�jh5|�������Q������-�C��󵡛��
�Gd���5ߛ���$9�Czw���,�&���I�}������V-!rv�ג�A�6U:IS[� ����S�aΎpZ�/���֠^��k��M�P*'��T.T�����h�r�d���]3�5���rK��t�4��:ED�V�|���^Ƭ<���ไW|�2ȩ���3`�d�33����Y�7�!��YZϿ��^uf�\ƙ���H�Hq�*B�	�UJFy�Q&�<8Lke�*�|R�[�<L,ʁ�Ȋ��;�r�Pf�l�����(�ɽw-�ZR�5�%�N�")�*� Yv������j ����Ryae~p�1}8�j� ��)�8n�2U��i�&sr��$������1���؎��o�4�bvL!��]9!>��♉���2�0l�!�k��n��zt�&
�ΐ������Bls�9��(x2Ls4���q���l����45��/�5��E=/�q 0!F90b��_��|�p?�9����	/Pt3��gTGd�YF���7
X����/�ɦ�����8,
����{���
ӊID����v6����ʪE/G(�u��ɏ!gW��[,��M
5:�}E
�3nHU��Xh;t�:E�Y�I�F���o�y���o�����
b�Hv�oW��P�^w��'y"�A�B��B�q��)Θ����MH���<̋m ��Gv	۫f��e�$x�����+�S#@1l�c\z�suGkls'�yVԧDJ~�P�@3�2�Rdw_d�.��  ��Q/��Z�)u\�d�/������օ�S?�3���`2��1G�&�����cX�bðr5$#.!Q`�]�Wz
�� �I��
7��P�}���q�N�c=�����(�HR�'����8�c�lb�ɵ����r��A8 5�0qў�ɐ�zB��H%�=��(����ԗ�ו6L^��R4��ȡ�G��ʡ�k{	S+ݛ�[`���є��R���g������r�m]�X�U�c�o��g)EA��\��
U�%!1~��2���oߢ�ʩ�sV�0�1k&b>�+�vj#Ԑ�sx/ Bɫ�~�Tظ��iY8����[�A����!⾤PhƤ�K\1�\�]�Ͼ�r�)X�·kz�k������=�����uWC�3��핍�4weCP�X��2vW2d��\JZ�oe�v~_�W*<�P�v�@���m��:ȚQ�nsz��+Ԟ,��
�����c��e^6c����V�~��)����D¿�̌�!\�=BO� �ʉR2�j�~~z�~GP���r�v �&G�?03%�$��N��=;Cj�a�(K׼{�؂$yv���C��p�O����r�j�~�7ե�I(��'�.2�'p8���ul��Y�����^gt;��b�D>`�-.R"�חnJ��n8s�-��V�����Fd��u#j����[�V�np>5� a���Ǐ�!R�E� �6T�����ԓ��'��9E�]�^�5��ŝ��,�7�
WmT����-���)���x�S������X�R��y�K��*��q���4��w��˘Ʋiꬋ8@l�U5a0h�;��Z,�,�u�����Fy��<oA�a� ؑ}u��=��Wl�`���*��j�	J��J�gE7_�N�WM2�*�ʢXì6ԫ�'nGpO��o�s]5Q������9�dn�a������C���-�{�a}�-{1Om�֞7W.h�x����#��ٟ�3݊4�B�/V��|�,�]m�!�x&VK[8S��A���S���$���[�ZZ�ְ⇡�������g�LCj��	!���thQ���$� ��<�j�������|'�UrGu'tRK�͠?�<�̕�����m����Q��6�T*u��<�Ih�v[�[�2������6s�#+���[y��JD��x�9:p$%�.�#z��0J�P�)�ٱK}�����Urgc��rt,�Z9�[W�.�����9]��Q�c�q����A�֢�K{��R���NY����M��h����AȚ�:X�� �r�3�{���-�}q6r!�s�SG���*�P�2� ��'����}M����1T��i<�/x+�3HM�&ǌ=�� ��b�2*��m�3�B�L�J�u|q��ٶ�!/�JsW��_yƻ��Q���mo*G�-䓨;���BUR��P� 5�K�4����9J:�ҙ���$�gu�p{��`y�,��-n�`s�:�����"b�]�T/k�#������@�~�	0�B���1�L���Ait�ĺG�����*%��������v���^��П�)=�L������'K�*-j�	{C�`�;F�@>|��]�Q\>�Ѝ�$ęM⋾���'�%]!Q8PE�<�6�-c̊�X%������ŚienZ3u=el���e�[0?��!�v�A��(��j3�d9k�J'#AP|� �W�/�~4�=2���T@���F`�J����F�N�ߍI����kܨ��o�óM\]V�q����۶	��, 3��m��#G@����V���y�1at��D�����_JI�<���L93h���F0$��C؝��,*��	��x��I$�����%3��1���a��u:iH�
`��X1��H�����\�rU�㛖K?�=�hA���e%�#��c����R���}��E�ύb�ń����4���9��Bm*|�0�d}
�	5h���*�i\��50���I�n��Tp�/f@lόƤQ���I�ً-�N�́����ϒ`������}�T��5w,���*�K���~7�=L�^���t?�4�Pl�X�־EDeR�5�^t��pP�|�	,jĿ ����j�{��b�ٯW&�6�Oo�z�Z��+ۨ����(��l�E��:\��`ڕ��D}����ٶ_�aգ�i��D�T��N^�h�q!�	�J3�5@�e��^�Jl�̴�mf�P��F
�g?˂+L0�gI���g{���
1� �֦Z]�UY�g�N�s�QcF�=���&��������80h����؂T_z�l#t��Xȯ�%'����1R�[�i�L��.�q!U/��ΨY�7�)���Qhg��t�Yŵ��_`]�����Myb/"����=�uTf����/��aI\л@,�h�wZRI�0@�{4��8;(A�txwy����f�RnD��`���׆�!�H`5i�aU���{��>�_z����7o�j�|�T\�eHe��`�����[l�%2�ѝ��vt>���j��>0��ݢ DNJS�z����e�Ed
����9}X���$��?/��Sw%��K;���	L�~<���& �$V6'^����㈹
|���&������U�B�׹D��炐��:��p:�K]����;W|r�S9�I\~G�=�	{���9��i=N��N�Ci��\�F��s�7��ȁ�F��5rk�k�e��	�',a�'U�(�\�����m04�8�L��o�<4W�� ���*wCNZ��! �~�h�Z�#�40g��]�ț��Gӿ�8Γ��4�e-6d��<�i��"��3昨�{i]37h�?�P$[�ʍ8MT�P��i��=�:ō��JT�h�]􍬌�Mv>�����_�� =(��Y��5��L�ES���Ri��x엖')jP�� ��KG�!���M��1]d%'���B��|:l��\<���N�x*�1!zB�6:#�ҿ\��LB`!�E�) +�3w�s*��p,a���w|;j�_�*,A��^�a�Q�V ��������㓍�>y�C�}��Z�=V��[}05�J�B��;\VA�H�$\/�3�g��3��~��r�c~�)Aj��1JXe�B![�h�=�b.�m�=�e�;z����֙��EQ�ze�P����?��̓���\�u����,KGC}��u���2���D��`�ӷ�,x��:X��6������)��#s�BEԥ!Џ5��M �M��7ڼ�-�OL0*�	��_�������x�$tuJ4>������L�<9�f�C�]��n��b���s�I�I���Qk��r3��� #�7��Q�Ǉ�<;~2�}�iƅn�h�8g���b|��h���t�����|�&KoK���7tl�Trj<z_
~:
A�+��P0,V���e��;�m��G(@�2 ��E(�_��o]
�URM=�z��l�L���D�4����|u�N�ȝ�M'i��R@��a�l�>�3:s�Plh�ښzmKm�E��i.ZJ"e�\�M1.|�S�M4�ۑN�_:���10���_�ڐRLe��u���-q�{$Q/�+|�]�9���7:F}�]u*\�'�I��:
�����5�3l��\�����h�@a��}ȅt'� ��y���$A�|CҷŞY� m#��5/���:I���O�#S�L��Ao�H����NY�W���PR��+�V�r�4�<,O�dKt�C��i��L���Pw(�99�GF ��
��oL�2d���i2-یom
P���4���ح���^�"����Ċc7��Q��E����Rg��%����l�`[��| �LX4���/�S�y�|�E���@yn7�]�+�=�(���NB����KH݄~	�!7�O�![�M�L�3�F�H"�/����ճ{}�%�Fy�w��f��ӝ��)�[����,�?���va���AN-{
*�O1�| 91��G���E �K3�~��-x����G�J�jh���ߙq��<H�|��xH�c}P�u&_�)��� ;�e|3�|YP�$�&E�얖o[|)#숣)�g��N�����	]�S�,��*�4����eb��ݧJ2��iLv=�W[�⽤ωR�����&|�V�;�f��*?��f����n澪5�숊�X�rɄmZ�Lk�q������^4�٫�L{@=�6ο7�Ԣx	� �W��ȁ�
�u}٠L�o#묕r���#U��c}�)�|���+��ӿ�=C:�e��ډ��_i�du'}�=;:#u5$h��5e	Ds+���� L��T��9�~�`b��%��)|�LAl����
]�ԏz(aɌs�U���טy99�6��h�e�!75V�;��Qq�ϯ���v��*b�.2���%[a�?����8���~��u'�h�۶����+{j�N����z���۫ճ��兞�ka�ޘ�Ki�D�$C���S�c��݉/��G�(#��q��5@�=n5J��Q�Pij��:�Ժ+f�rW�&��w��M��#����#��U[���j E��$Nź]U٘�D^�"��5�M�Q'��9�]�Fp��"��fF��Z�� >���n��cI<�'�Ղ��/�?�;��*pZӝ���r��V���*�e��1��q��+8�qj�pe��s��t	yv���u�/AM�p-f�&-lQИ�����*��?������������2���q{ő]9���]�B���O�8���Ӕ��mD���n�R�5z�s�G+�v<�gj����ưf�O��a!J�O�6�'�N�ױ���U����\U���lt3}����sT���Z:RpL�u�=����K}ϸS�v��ƃ�\DzD,lz7��
+>�TK��FT�tz���Ӎ��R��d>�Xk�/!Ŭ����:-���wk��e����n+��e.:��)��� ����C(,�����Y2��BY���*�ޢ����u;D]EE��k���m�x��A�^M/�4����r1Y������	��_B�!۽�)N����P9T5C/���4�^��7�E{󶭰���c����)��%�W�3�C!Wiw݈߷��^U0dՁ�`���T�L� �ҪAP�1	[�>�T�;N���1���,�~�8h�����1p���99H��Y?��2�Dg�>��G2I&�MTtTV�`+�Kr��1��ٓ��f���L�bC��H��Oy�:tW�e�{!�퀥�x�X�uNM�ǵ�/���臏�^5�ޘ�b��$��@���Y&��ݏn�Ǚz^y�۴ͣi����P�Xb��UD�u��j`ܸ9�� ���'�~ �������6�۫w�Wo�h��L�Ŀ4�C3@Y{���%�l�,����r�M��X�s���E�+z?c�·S���D�8$�}%���[g�1_Gh^��7�b�ܱRo�P�s1�� %ej47" dt�r�� �~�7�6x��w8��PC��qI�r��m�z�`���$��:j��7��3b�W�,;���Z�C�hiL��a{�ǦUD��O�]���~	a�� X��\���\�1�0T�o�H@�S��������f"��/���#Jʑ{�����M�*�X
v��f�f��̩���h5@;�����>�O�edGՎ� ���A�\��ء����?V�O�f��/g�ȝH恣�'�B�nt3{:�O�Ԓ�0 Xd�5I$�k�Yj�:d�R8f`u��Z��&��V���sa�\$�r\�l����oz�4�[�@^<�}����{JM�Q��_����qzI�(;�f�s�TG��|�x0;L��i�b��LL��z����`�ҸF�.b�Gi��7Ut�-�/�񢋼��@|�T���ƥ�T��*���e7҃��h�=���'�V)5��ns��C�˯�O(*j����ڝ�ځ -���;�J$��+�+3���?��A
#�YF3b�mm,5�,
p�;�R���'�%稦���6�1�LZ~P>1��	��L6��D=U�ڿ��\j�Gr8���@i|"��;�R$w��t��+��lSg�ǫm�-���
d��yè~(o��V�wV������+a^��g��G� �1\�i�f�>�rv	Z��Ciw�� �ACl?���y5�	��P���;T�o�¾N�r�YQ3��i�0��KE�O "vh�52G}�P���3��p��؆!��o����^&h}�,�w�G���g��G����I�A#�,=����}`����<i�/��s���0H�W��0�&� �=^���ްO��1X�#/*ޡ�M�~����z�<l�=���8\k��]�f�YA��1Fm0�c�-�x�&��tM�����T܊�K��[R�	�3��x%\Cg��f7<���z.�+��\��>�rma�-�'S9̸S�âV���\�����*�v�_
̸C�@@�b���z�q8��%ǈ����m����D^�,2�އ�z��X��j�w���:A��ES�V��:r��k�����D����TCَ��v�Y��:����Ʉ�w�>��p���s����I�,)�p��eReF�1sƀ���/���VE�nB����o��Z�Fn3x���(���
���P8�3"j��������M�o���i��,�Ӣ�ؤ���C�����I���|�{��?K��=��6�ڊ;�W�ʊҿ�ܳA�&<#(���qfNK{E� K��u��q��v�,�Ǒ�E���j������#���6����:;�����Q��e�����Pn�T��u���r�D����`x�R�l��"Kdg��ƣ*���l�����u~��*��M*w-�o&?y�}ps� ��[k�8�K����V�K�<�&b=�ڡ�K����U	���-�(NC"2��a�_SM�_s�7[L"mE[6%�R�S��q��f�X=j���w"�R#�#	�S�4�Сp��G�ߤҬ3W����B��a�E������;�M������ZTu*��zBS�,8d:�D��YV⽐�3�t4�T|"vAD)�`#zǱ�I�;��P2L�W�۾���ma���{��L�F�&��b� �'�x���B�y��~��S*���S|2�[{x�g��׌'���O��L�i�N6ӆ|�g�1�-A�)4��M�ᠭy���]���zكyb�!P���#�����&Ah���fF�ͻX﷊d�`:��v&�?�ܐ�������=>��W���|ts�L9�YE���f/����9ض>�%T�?2C�ȃ��1�Th,ц$՚�1�T��5p��,7�Z��j)9�MI�XDK��P*�bI,��N$B��*����%![)��R��P��`C�8J+�|/�qpƇ��W�@�{��V�p䪷OA�a�ʪ�?B1۫gvݶ�#F���s#��>���3��鯖�\�����8��¥�zɦP�O���z�=&���~����!��Wp	�#�
� B��G|�B͖R��۫b���"�I��C5P�P�BM�v�W�(j�:6��ݦj�b�д0"*O(y�XS��T�v��.�ۡWs��Ŵ��v	�!9���,�7a�_�'i�^!x�y0vd��.[QҠ��>Ÿ�~�hg`P�UG[z�3[��C�D�%ͮFs
�O�lְd��4�u�B�.��/䝵�_�ܭ��M��Ut��eD���<m��v�<q�vۯ���n���}(�zG���!<X�Ϝ�\hJK	$8φ��r�;0�^dP�u� 3�+{ �@!w�+'���s�'>fGּI� M�?'�|V���7�iW�~GR���6����Ys���,�Y����I�A�Z�� ��&����T�3t@(뙶F2����AZ�[��|D !�{T�Ԯ�Q_�4dK�U����al����m�-���ZUEf�H��2S�gO8��5�}��?�A�>�N�ލ��tT nh=f��9͐|�	���!�C�~����=[ᔿ�bғ)�����7�f{?I)"��gj��{����	����2!J��>Z�(k݁��s�I��2�܂��`7�Z��k��-�����&�.G������e{og�"�2|�
��aKJ�Q/|m�&���U��V8�����2f�^����͜. ���c���I
��J7UD	_�3HC8�XP^�|�H��Ĉ\�Սg��1���4npG�bUS�:��<��Qa(D� �f��A��k6K���n���~���K��V��3�wY�<��%X��� ^�z�bQ�Y��:?��O�~���J�6�f�~g��F�4���M�6�� ��і��e�A�,�C��s�d���4^�o	G���XH���"��LE��yx~�]��V����!fR��_K���vw������O:,B�&-/���r]����	
�]���K�:�:��6���U���P��߸D!�FgMFRq��3�M��J�V
%���X@d?�� >�|�JFv��.�`��/������q�Gͪ��
���q<���Tvcژ�67�Wl�@��{1B ��	�"�pcq�طo�$�A�	�F(x�ķ�c�@(<؟�zW��0ߟ~��2��9\���9�Z,��*I��v4e�d�n���[E��Iܸ֛�'�ZA3��i��ʄ����_�����Q��A��1�F��<ED�f�tL��:譩lp1'�%/������ct���{:�8��� ����V� ���Gp��;ФS�����4L�p1z�[�����V�~�!-;��xl8��f�h���R�g8�Җ�r7��2� ~�ZE_4�>�ܤKb#i�ita�tO`MB��d���L����>��6���sit�����l�?�1C�d5�4�Ӄ�Z=}(���f�`*�_�M��N��ِ�f8��	[���!e4Z�@=~�׿y����Gy`~QzO��a_ �Z&~��x|L�Ϭ+袒s��tX�|��c����a�c�̝P�Ϯ'�A����TO�38O���<^�Y�.�pμ�8��$tD�/��D&�39���0��|n�H������BvՇ1�;}����� ~��Es��5E����hHiKSM���R�	)��ٰ֫W����d�N'G8� %zw�����*�ɔ�m	����`'�M�����BWN$F\i��I
)��"5x�E�ʓ�O ҄M�-��G�\j���5'�"��7�o��l,:u2��iK�k�n�������KW��ڔP�N�,+�)�Gjx�(V�Ǣ�zm!�+��{�'�t�ZU��(OD�7���"os:��XT��nA�9������d�'��Mz�(%��D��@:��4��ڎ��ہl4eSc�g��K����7���>�K1� �"L?�'�J�ӽ� ��%���;��Q'�p��|
��xJ���'�n��B��TL{��=�K��t��^u�C9~!����BXa��'~�x��4'��3��VY��jFN�fo���9v3@�?h�=�(G<B��G���י��>�H���-��۲�R���^�&@Y��2c�P��S�P5U	��+��w��q6w�D��~9?E�z�'`��7I{a�c�g�&��j�!����P�C>'�G���9�׭�\�on��%�]�;̶W�<�p =����;���E�*sS��~�J,j����m�XĮ�X�ED�6J)3�n�`Ŏ��S}�5GD���GD�ORA�O��@R��
�n�'(�� ~"Q�9}fr1UT��#K`2���a>s૝�b0Y�yGq���L�Y�Ҿ*ÄG��>�Ҷ>@���ں��!���(0(,]֎�+�ա��n�^x�k]cƤ�	����g3+�oԄ36ګr�<as�meU&�}ų�CI��~��U�`F[A�2��� JQ4��i���PT��=V|4��G�')��,$bm�M�vzԘ/ߢ�䩀�	m�����e�i��S��(�]%Xp��_3�T��M�~����%�w�o������Qc�辀*�@�VA��AT�\�(���2B�n�+~�nz�X��5�%��-��ۄõM����'���6����Wg�rp����J��W��cf̨3��� ��!�dI���Ρ��.x�
܈�-�����n�
�t���W�� �~ �W\c�?�w�UiT�᳻BlY�y�W�y`Δ�`���k����w	vZ&
�A�<v�#_�?���*C�������V�Od�����������I]Vnq���\ ��B,���H�F޵s�ߪ���/F��i��gt�:�K����0 ��a[�H99���kt�g�|�B�r���و-�ͳ��ǣ�?��C���T�-���\=��#߆C����
J>�=U�*C�P�4r����V���9B�����2��c@�b�@u�����O��^&��į.�sf���!��S8C�
�f�ӏ@����
�}��1����:�D���Ԣ�%�T���o(�2�q�.~�!S��������)�=*��o��W��]ৣ�К�Sb�x���Sm��!���g�m"��!�
 W��:kd���}n�3��d���/��;����81p~#�!0��Ĵ���>��L�9��!�5��5.�BV*�zxs��ؽv4�,�n�T��<�J�<���+oV�F#�B�X~�e7�b?B��� �!�w{W��6{�y��1�����ƿ�p͎�o[���*�ٕ+��E�RD`T�d�����g�u�o��VG����~���I���pX�F\��^2�ؗ|��e���߯���z�k�tKڌ��WtPӽ��ĉ�>g{F%����J������.. ��i�[ֈ�����w���/�Fx�؜��F�E/��z�G-9�hFg���iRQ�8�C-
K���IS��>�n�:d�>Rf5$ ����7\>A�|/��"Ϸ����a�O~>G2� �H�z��M��tu(S�M�ş'v4���L|W��<z�Cu��OR�P�n۱���/�h��@"�b�ئ�L?%i�$q(u e�_А��	�V�����iQ����a����a+UBa���g]9�n��GTߒ<,z�A�I�xA5y�<|����������Uai(@j�%�\���t�Y�gw��ɞ�z��I�<�7�a0J;3(�y�e9�2�S8�:�cjTʚQ���дѨN���~��Y �`��s�f��)���H������r�F��2@Q�9�Yx܄�_��e���aH۽��D�� ��I�4�q�����_�窆	Ɏ��Ioc��V������x�խ�wbVz�L&��'�{�*������G����Ԛ�͈tu���[p�L*��F�&���#��{��e�̴���*Nc09H�F3��g�����>n�|{��[䥶�B^�
�@���Q�I﷿�R෎�R->�X��2����"C���������x�d`\L�Y�#��!�9*��*�RkfeQ�w��
C����n�5j�rI��*D��N!q��K���_	E�e̍7asӽN��.�0 [���7�X���1bc��Bz.N!2s^����v���G�
��F'��o�]jMl����E�iPLnfyi�$T�XW����\�*�F@�?5��v��;ŖJ�.}��;Z�v�:�6A�>_|�7/�Q}��i��W��d��˶��XZ�!�,'�f����%��2[.�N�|柎��7�@����~�)���v[������E�G�̳����TA�8��Q�o��x<�d�v#=��8�-�A��"��vw��?�J�����}�V���׊G�;^ģ���=�+��6-�H�f}$��X<2p���gmj�Պ�w�w=��P��C�+�����F�`YY}�
��v
ϫf�����pft����^F������qRu�Ѝ���3�H!�8�ju�f vw@=H�����RR*�X �M.�E�P��Z�Pe�T��jz��蚓w�V��_-�8&F�"r�lB���*���I��5�ϽK]���[0<�tm�沒�yܛ٣{#��\��Q;s����B\��vm ��]���<[����˄d��'�*τ�q�љϯ���;����]jך�ı��8����ׂ��0P��TY�Sf�T�����8�$�A�����fN��b.��XB'��lO�l�ǵ�DXe����d��y{���k¡O�N�5����r�Q^�6�}�ܵ��Ɲ� ��𽟊�?�9T�V����j���<�?A�fJ4��wob��eVuRI��ȭ�(#3�����)��s$@���<S����m/�>>��T?+tPɒ+��]����GV�k3�9TT�IK��8n��I��?%�Bl����OII4 XU�P�WU���"p4y��o 2�-,n:����^�eRy���۔��8[�0d!\���*�{_
`�iC�5���:M����o� �ш�' z���O�?���Ѯ��+q�c}�^+t��\I���D#a+��a��GOLM+g�	Y��}Ǭ�&Āϣ�y�w,���FF1����@<Ɓ_���/���ꛀ/bz9�mβ(J@��sO��Ȣz..^;
S2iT� �v�_���n�/&���>�:�)�?����I���l���Axz{��៫x��?q*��\ G����*��:%C�T��ϔK��wF�X`�B$�u׺����YԟtJ!U=����%�|bR��hh�&t����L�z����S�t����1
�zE�ɖ�.i��^W̷�K��A�l��(+Г�Q[)�2�ޛ�4\vx�`d�x�5�V�ی��C4������Uh�_	T�#	��_�g,d�}�2�A\*Dʒ|��.�+�(g̚Ӱ< ��,�L��G���������<�_eevֈg�R�[��?��� 2:6�C����d�ƔuB�(����R�{��)m+�eZ��^�x$}㠋KoS)�lZ�)@�ق���,Xg<,�QbG-O\�O�S�G�1�>P\:�z����A�;��N*���?w=O]�|��_�N���H�{T!�V���{VM|y6U^"�k�`��RnY�V�b�ov��M0nh�hq��.�1�m0W�x�G9a���EM�D��C$N��e@��7���F>�4o�m����udv�v���BZӻ�uSR;x䍾l�Ҹ
�c�Ak��8��?a�Nz�B�ϙs�Ħ��w���8���3�F7���Q*�rq�NfqK�"������cCkN*:7���%V�� ��k�#B��4�38�.��T�v�"�i�0�����VҕSS�nJ���qHQg�maN��#F{�K��//�p�܃��!��Hx��a��P�H\��(����m�z��4q���T�˺�/�OlH�Qn�bL&��:�<^,פ��"ϒҥ���jAu0w���z��^=����;9c��z�b���^�����-j�?/��$�YΎ��K���|��L�!� �Y3���)�Wq�� r&mZ���`AlAh"��D~ �!�s�-]��� ���.4\��͹���k�N�s��a!MT��	(-F�p%�>���1�| pz���Z����3��Y�Ǿ��WP�����l��"!�NaQ@?���M� 0{��A~�x����V������A]4Y]��T]��0�lvaa4��g�_N��L�ח}�^�V0~�C�8�ܓ��.c�h�QM���8�@�}a����b�8��̪}�����G�B?P��|r���E���1v���q�>�r�"�z5�;����>���G���Э�1yPk��j�j��C,�G�pgb�ɹ�%b���[�<��hD7�ϽȰ�`f8Sί�m~43z4�d��N�A��tlRQgF���zؾ�7h�F���+rz��)\���]�;lW������&"p-��1�hC%�?7���y=eX�)^���f{�G�.Q�Al�I�Ϸ��>4�*!'X`g��� \ouD���{xf�^�^��lM��1��eu'o_�$1�ZC�`GU(��iG�'��Y���Z�:n2��d�HԌ���5֍*��"�����N]�(�`/mP���A��OAx(c���k(�lR�X��<<��鿀b<g
e���Ȗ;�,oDlo����ܴC��^�� aUY��im��Es#�)ۑ˗���M6ck N�<lX�$/�&l���=�X�/�f�<�8���'��(�K{n}�Jö.4�O�+ge�䃓��{Zbe��S��F6�Q���;�i���r_�5�����A;�a�,���P=kЗކ}@_��S���1A]!�']�c��	��������2�^�o@B��B-�9b����i��B0�L�����\U���2J��9]��k��H��f<��_􎳼621��S���a����8�~?Ʊ��ͥue�!�8&��D�C�މ�Q�E�y�q�Y-�##������JеN0N�?�EB��1�0)v[wJ��Z$W^���Fcԍ���?F�nTi	2�(�jo"F	��)Ԣ���E���p���G�V|ˉ��3���SX1��TO��xdx�[����7��7�n�i1�����,� �$����l�]Y� ���p�־�T��9�nnm����Pȉ���45��V��.,S�5%�:XPm>�5B�S]��4�uQ=@T�륢k�&��VJ��ߗ�B�]Xhs�l��$^k��Y�����F�b"���KMQV�H�]��2�X�c�]��,T�𪁥(��(<�#8i�?�<W�P��ͦZ���+=o?>�R��f��&�R�K���F�0�!M���H�N[�(�C(���!H(^gvԞ-�dUl���|�
0��[�u7����^DD�t^�BГ7lV-{�A�:��l�㳵Y��)�j��:iE~�w;-CϏ�sN��"�J��ߓN2��S/���V��F���s�&\Zڒ#5�����tZ��Xs�n���Z>����Tl��N;0���A���ު����k(Rx���
���S�.ذ�hV,���!���#f+q~穊���Uw5�/Z/�|������x�y�����J���� 5�}�P���}��H��j:]��ebw\v
h5�+F ���yw��CM���.���@*(����'�f|�;j���?�bN7`3	�q�2\ y&���l���U����>�z1W�u�u��6�^�h���֋I�T�u��|dA&��4�lCE��m���fM~M��B�c}�VE�l;��uĨ�tT��ȃ����Tl�@W>�t/���^G��	��:��WC��i�������z�1(���~��_��Ī�X�=C�ldM��{�v��.f���R��V��a�����d�?��;4����qS��vo��a�+�{;a�΢(t\���Z���DUʶ����ڃ?�Vd������>t���e~-����1�1���NS�E���*���aP���E��V������_���e�V�'u&�V!�ϥR�жu*��i� g��M�o�v���l5�N��#>X��R4��~\�i�*gx�*�X�%���]�Hr��>�"�7��X��"ꧧ\��2��O���z��_,b����!��Y=?���l@��������e�<g�� �]��sv=	 IWe�fC�*%����懹/n"�S��/#��*��&{�5���S��	�H"���k�l��\�:E(~������>0�	��t��#O�MJKOWu!5�K��x(:M��cY���>"�_�>�/E���#B��Z$���� ���?Z���ȼt�
]ߒ�k�S]�ޡ-���X�|��4'���p%V�|�.�ab�ʈPJ-c�З�Ţi�@�>&?s�Z��:h-�7�aNζ�K�?s���D.�6�5\I/�=ԧ@B�N��U��v��dń��T����2���Uʰ;�B��ٱ�Q���0)�j������40dO�uR}Lw�ow�z3���d���8��	!4�M�ඔ�L�2�$,Ί`��oĲx�ݿ��݂r��{VR�\�Hσ#vN�/!���V�;!�WI������9����`
#���\g9>LH/��u%.�G*�\� ���a���4��p�	>&T��s�%NS�N�z[��W�2��`r����Y��8�G���6���N�E9�AQ�&���c��NgtJ�}�T
yd��va5���?=ņ�Ťu�*vU�8�On��|�3�=h8qW6������AދG��QB��6^�� I"u��9� ��b��I�K�v���;��r�H~�x��H\���گ��<A
�T�8�5P��_~]\çT�f�3���4�e�7�@�Wq�i!�7ú����bʉ��"#һ�8�`��N���\�֛(j �o����u�M��y�-⃓�����>'`?]�,���:#5yݛ|xOZl:�',�Ok@)m7`�5�j�:����c����2����"�}WW���7�D~��H��R����'�|������_��Pc���9��n~�&�Rc��w󄳗�ɘ	R12u,Bή�]�w(��T�sht�J�纘M"��v���;[>U�#�{Uѕ:�W�[���8R���83�Wh����Ǌ�tS����$+2x�p�#3��[�G_ݮ�oă��3p�[m����Z�!���!��p�@�����W%C�!�ȏ�a���}w����hK9� �
k2�Z]�������$�o��EwO��~G�(�	kX�E�D��otu�վ?�ѦV��:8���G�� C!P׈[�0��{�r3β��4�R�[�P;ɂ
;�.�B9�/��z��Jr����v�2C�{��-|L �:vC~n	�gȞj9W�6s�7-�s/^�ĺ�?�,���e��c���ϢG��+tQ֊�E�uCm8^C�2�z�������qH�(�u[_�І�	[�A�	��Q����I��`���B	�/����&��i�:U,t�t}`��77f�u��=U���}�B�f:P E���4mRy���1�1d�ohuߗ/�l	/g9��2ڌ��r$��T�$d�7Lg���Zg��׋��,TK\�7ʶ�%�:�٧0U��B���`�o��	����Q�fq%��Ơ�\��2���^N#*�@_�����'�h~6oU�<s��h�z>�Lj<���%�v�^� �>�jt��Ev���`^��+��9m��=���".f�HD.XX�ޓ���4�5� �Qj��T@2z��8�?��>������Gc)�8G��-���5)}k&Ng��������S���w]��Y(9Rx³��� � X�z
ۚO�>Lu����h�0�O�H?�:^������'eWt[��nbJ+����ڃ��j�@ǆ��G׵An4'�,����U�Ή˭�䯑�|_.�+BΝ+�}x�6b��댩���T���%�����gY��
���-�J�#ݑ�ĳ�鰯3�˶c_Z�����#�AwWDL�)������;Ş�%�9J�^�%N�k"tS}�HC��w�|�R�ڸ�'���./�g6|���5Aߗ�`3|�6���I��M��)��^�4	JI�]�{�k9<}�𔶼��>�������%Ew��n��V$��w�-\���q}�Z�a ��]��/U���v�
�R��� G3�6�GH�^��*����"�ΤF+�g�����"���$A�����ӍjsGi��9�W����5�OS?�|M7]��:\��	|1�&N��-�]��,��D�`�D>��ja/�"�lMd¸ʼ6���`���L���&��
����ι�_�.]̧���"�S ��s�TvP~~_��=�ٺ��駿J��m�|���d\<H��F�n5S6`Go�r;F&���{����D�$?c��C.���%�{��X�I^���Rf�љ(9e��m�O�"7d-?]P��j���z<{>/�p�H�k��Aӗ�ǝ��^5��m��HV�i�}�@s�i.$�fk:��t�B�N���/e�Sn�0�ef@��������g}������vg�?�o�V݃���Z��p(�K���u��cɄ_oe�Ib���a�7�m����h~��E��o-�ϴ�7X�Z�e�B�C��\oWXM�H���� �_��6$��c�t��H�ɞ,���Bs��O����"_�	�	i���Jd���n��nri�d�}#��IK����wTb�qp��<+ɟ������!����	�i=��/C3)Q+���<��.i��-͔>r5�� ���]ju& E��sfH9�o�p_z7�|��qU<3���{s]��ŐkH���ٱ*��?�]3�`�s�=��7*���&zƥP\HlՐ�Q �&�˳�3�P���O~�5�nB���N!�aѴ�ݼ�p��pF:�쭈�g�K���>ij���v�ӱ�<$�6d8��E��LG9��)".�S��1�����F4��b���-��83k�����~{��Y�d�*�U	�����0!��%����^Źz�f��/"�
:�"15�O���������(�	{4���<Ew�F�D�R�@@��P�d_=q����@����keN��<n����::5���!����ւ:7�<F�Wr]��R��і�.(Q���.+źo�������}���)@�YH��]��G��h�X��r+׊g�:��q�W����C�j#E#5�jo���*�̢`A'O�tR4�������Wَu��[�W1qBE2�ڠe[��Б��$��utKoM��=XM�J~(ۚ�f8tG����v�5�1O��(�ַO��X����K�,��u�J��a\v>.#�����=W��NOgk|�O5�(��	�t�SSd慷���Z��~��!u^��&%`�-��x�6.��z����t�R����Kk
�@��=8S������[��=�z�8�tyN�.��w�-114 ���ٰ_!��To��:��A�!�2�)�n[��N�I
#��<�  ����$F��d6
d��.(*ml�?I��+	�Mu���,�׭v�*d�}O���|,��0\\(�x����3�9�u��0I�נc�5�neK�O��"��u5Yy݄�7����1=aPj�	�@��O��|i�s�n!J;Q$ʀj�_o˭7c�2E��dH�dh�G�xb����.�>r�֣g�q�����@�G�Gj��EJh�(�$l�.mɁ1��x>��/`րsK�}�8ⵕ�<�Ku��IL���{8��i�)!�k��0�}�$����9L9�K���];~m�|y���f�&X=Ѓ��o���w��_�.(���6��ys�Cf+�K�:D..mؘ����T3��ד+�qS�������uU�G�󥔥̈́�֝��A�w�f�O�$
bh���i#` �WtR��d������xA��eK��ݏ@]�^��\�xL&�v�3�� c��˟�3;9Y3�Z��� Ǎp��Ru�%�S�h0��m���R����g�~>��H�R�u�;�����h����mYvڍ��La�$�n����ʼ�c-��R��w%R�ڜ�[�2(-�5_�B<O ݲ�Kw��'���һ⤉���W�YXw��	��+������k��]|�N��F���Ѯ9�_���FL'��-2ʮKWc�Xd�?����5��0�� �E�͇��歄W�7�T���zd�b�u�$�<��]�k��k?�$���.��w�> �xw��K�F�2�R�*X1�=5k@q� �=��m����/�bIAP���<¨9ݕ;a��i��2���8��&�r?w�MѮ�*�	ҵ�����3�^��5�*�d�'��Q�|<����U�Wa��V�Q���Y�PZ���5����E&��4��h�e_���P�m@�2:M��i|JT��� ����}!�4cr[�=�㐥+vp@��uV
akO�Ŭ1
��:��odW����i���D$��6T�!��bJ�S�:���߱Zch���WBK��)�j)�OC	�d��/�E�B�\P�3x�GN�/�ВJ�����o$ݚT@��c�3���V�=�Q*���Ȏ�>,V�rD�i��}I뼽Y� ��� ]<���E���In���p[�V�~�Ӟ.��m7�ɮ���Ii���>Uk�^G ��C�*�Q��123zk*<�Z��������El��k��)�sme<;#Y����%~�4�.�E�4��B'l�>k�M̟%��;3�vNϰF7�	���s�48����_Fb_��c��?�L�=�K_�t�a��<|�F|�4b8�U�tD���N�\
��t�q�jL��瘗�Co,�˾����0�g�`|�y�Ӈ����6)⊶`�ӚWs�`�:��ܠ��]�P����K&;�(�|
�
�x�`,~WӢ�/2ҝ�Р��n�s2H�jl���}�;BFR��70].F��x�Z�>kj-}�E�-oE�K舧Jun%�@������7\���n���m�m���G���c�̳�H���"Ċ��`��Ç�w �	�e�V~�	tDw��iTM��-��	�ŅR}��HiƃNZ�:�s2�y䊞���1*}�W�@�Z����F�\M�К,����{B���%�uBu�����1ؠpf��)j��Q�������G�*Rg�jm�A�\���ov���ȍ���G&���&�X��&���.�PU7ŵ�%ҁ�;���7����H���x�n��[)U��Y����rъ��s3��71"�xUC��A(X;v*+���අCN���Z��c�?����*�����,�ҋ��e�Ւv�%X �H�ѓ�.+/�N�GHF��n���M<"7�K9�l�f�)�`[b�j���f��'�R�n������'<�0OѢ^��]�՝�U�O>�H��b��<���
"H��7-�ߢ���L�^�QA��T��n���'Q$}Z3�kD$ONT�?��'8 -��ְ�}�n��k�BI��_�![i�BV�>fz��a�Id���iG��r�8W��+��S�Ak�7�vZ���]=I��W��,Vx�����|;���>iѐ�<���Լ߂��I(��r��N!��ۨ��Ц���&���!���IM�V"d&[��PD�*^ߦ���v{��&y�xI�Fn���{l웇�ٹn'_���E����)7�C��I���)ճ�?��)�V^o*j���`n���9>�n?Շ���v����w�'o��iwP���j:J#��T�A�-���搌7b�<�+E����v�'[�Ɦ���%z�5p��������=$r�(��td<]��ٶ����#��;��1�)
���U�JB��*��[�.\�(upb�a�DhEJ�n[k���\:R���J���Ny!{����k=\���R503�*v�i��� ���xp:�+��g�&d"�*� J�ҬjY����5�g��B�`�o �QͿ�%B&BZ
MP���V`��ōǭ���4@h�K��l-��#%�)n�V��÷����y��1�P'%�!���� �f=%o�x��@��Wk�;\ˮ�u��=-�ː�]�m/��R!�U��ē��	HѢH��y�z�	k�Xx�ڤ��K������x_�T/i�X3�$��2�,�\	Y�rv�ߓ�tJ����#�D�G�}���s��wO�?�TU��Ȩ����P�i$AלP�)�TJ.��+��Tʔ �\��q�%�.��c�3K��cy�><�Y��3��`vm"B܃$m�ɌX�:d���K0Ԙg�B2&�n'�8e��(%���[I[`^�W������AI� ���+E�i����,�3��ƕ���^�ഖ
��0�ר�;�B��?K0����4
,3�
���(���%�BF��5��Q!��������}���<E�� ���na�P�3i��h>�S��V��e�~�H.!G�L>g=�D������+�PT9��4[�E���X�H��"	x�F2�^��D p>ԣ��_9h{�U�i*GL��A�h�f��dWy��pb�_ʬ�w�%.B7�+�Y@����3��U�����T|n���g�0���X��!A��v+���������0=�Q�^�)k��� �_v�oa�'ƚ�2igu��l�A���&O�$ڊ4��چ�QB�����\��ND\��ar���Kq;u:�.!��}�op�F��h(�]J��~K!Ħv����ڥ#ۉ#���=�cm�X�[f�0�@�������W��eq��ƁP6��7�wΫ�N`��,O��q�_8Sb�f/�b�V�,Ң��-�zG�!�@[�⢐",���s�{�JE�mXk�����h��F���iH��8���_��9&�����v).`ڮN^K*F�=���x�I$�WS�aPb�mC��*Q�l�P/��t�$�}����6ԏj=KӀ<ih';����c��,�:��W�{�=8�d�ݱ�j�����{�J�� L#蔙Wxv��!2=Ε셨�����!�.K�^��ڤ����*0H;��ȓ�V��S����J����o� �<����64À��W�~�:�{Q`����l�1R솿�L��<>/?j�x��
�$�'nq��
0�2�h�t�����*�x�
Ǩ��������PP��3b��
OV8� ��u�).1�(A.��5�;i�]e�e劻pk[�/#W�L���gss�����]k��ew�|M�?��/S�������:]����{�韲=B>24�aWw��x_P�b���D��T�mO
Ly��%c�(�_v�_^gt�viO���a���%}����5�o�<s�;0�	\�>i���+�w�bF���*��
I����J�ÿ&�W]!�)o=��ΏQ�L��7�_?�|�jP>Q���H���Q��Jm�Q6`�o�I(�_+��Xb�lo���X$��o೧��~ػLI|�HAfu���z��;�V��?@��/_�_]xN@�ΦN�is;Я��A�T�:������"œ�-|�����'��isEN�X�Q���9�L�8u4s�
�t��ۺ�lf@��R�,"~��%"�酦 3�`�
��U^�T.N�+Y.�Cr�'�ڇa���i0��@*E���A%\��,��SF.�!X����V�������_���E/,����q����.Xө�8�pc�i� ��@Kf��c���ګ��h�a��\�s�:7G3��D�-�yR����劐�ѿ<B���^7��͈x���~0{��~���^�;z���{t�tm�Y�Դpx��Y��Ag=�q�m½��M��RB�I�J���ٺ�V�p�۩�ֳ;dP�����3�FX#��ڰ69tB\d}�QG�U����I�.$%@�[c��}���(��ch��ևRC,<}�g"x�eSŖR�����\	70�=ʏ���=6�,OR�dB��!�l
Mǅ�J���K��%a�r$��<[2d�
C]�VQ(�|CYd�����*k��ѝO��l�4�U6������T*�f�O�6׼�SR+Zu�݉���1/Ma�76���(.S���G�2"F��'3��?��ۡ�M���)���T�!n}6��r��F���{��""��c���2�)�t�[wJ��������v��'��A7:&>�@5�<j����
�E���Jx���DAb�����Q�}�,\������;dO�.�|u|�i�*��O���h���h��켅�J1h`�X��G_<e��LL5��Oď롹�lB�#�Z�P��,J�K/��:H�2඗.�P����^ ���J����/H��?��V$�����OVG�gr?� �EUS+����<���F	p�~#Jq��q-���DJ׎���_��	�槖0��n3&�`*jݖ!d��滑��� ��R�m�&H�Y$�!�"Л��k5�[SO�%>�N�\�ۄ�;\#a$`��k��]]}�ű7��C4��ft��ChZN�&=����
�J��z~��;1�.����{�f�2~�b�x��l�R^��䧜!�~H�g=#���,��|���E��M� �h��T�k�rjk/�,)V�
fR�|u��h�[>]$�b~J�ӟn��8��j�Am��ž{�-A x	���yl����G���"j�|X�u�5
BR�^٭g���:-JK�p�*ě��J�6���F���D�	i��)�ʦ�K	l=<�����MeL����^�&�}�Ģ"6�+j��9
�g'��;��8B_�o�i�w��n�G;�1����`q�rZu�؟��.���铧Zz�2Y��	ul,��?�q�ac!7��70x�Ga�,�cj�V�'R���m�ﻪ���N@ �O�@�&�Gt��Α�n�ä������x�V�҃���//[�-d:9�d9�a6fw�	��)q0���X���{"ph\wu<�"�Ѭ%ԥ�^�����Ġ{l�D:����Cg��X��O+�E}�����V	.O���U#����x��aJ���_.*"�h��������cM�c���T�(VL�ߗ��
���� 3� n�3��n0�T���^tˀF_��nF��yS��X_W���>X||��H�4^�M�&�1 Wҽ :J�:���u���M����8M�nx\��`��Y����n���D�/��
�z�])n�"�&$I�o./iJ��D�)�c�G�0v�ׂ
�G��[F�_�8���>��']	�
�B"�R.��A/�\r��Ղ�`Q'K�^V�Z������Zk�G{�ƩO���� ��J��?�Z�(������e�}su�,
�-�؋�I�Γ�|i��I����ݮ���/��;�6�_�Wu�A��&B�B"q��3e祇vgGcԽ4��4��S����~C}"�XaG����<L}`b�|�� ����eC��894�i��P@��?�Q��4�u�E��^c:�8S@{�F�w#^���� ����*sK��x��?G�sE�Kc;fF �����`I6Z�A�ɵ�zL���K��M[�IL6nx:�=o�[�a��7l�B*��҅����*����^rv�0r3�gd�r�������O���&����B5���v����'� C�I�������q�J(�]�b�=<�V���5k����i�F�{ �E���k=
�V�
�Ы����v	F5-2?jT��=���f��S��\˯��m+o�^G�^i��3S�\��ҙj�m<�!�X�����/�iU�4�F�V8��Q�J��	`��=�cx�D�X��y�,�b���C���џ�+,� ����ւ� �9��?L �,��g�'�!����\��P;���7B���g�D��9�nVlY02�Ttc��ox�]��0�(]��ݒ��`���<n����e�W����Q��Mo�6r�b0x�k՘-k��T$/됞�_�:xɄ�����D�?���.�`R��_�y� �}c���;�4���3\�׶���q�]HM�����"�ck�R�๜[�Q&�_x�~���;�&�<�K⩈�H�D��אQq���Ѓ�nKѹ�Ƽ���"���?>�>m��N�O�
��@���Ŀi7����U�Y���S5�����Z��^�����x&ƭI��gV�tܽnt���ͷ�c)Jqy� !ͧ�;Z���߮���-��ը-��PS��e���^gɠuZ��g��\9C�B�y����>271����f �cC���6��P��������g�Q�	R; X�~2bs���܋��N�\e��r~�F7�8҅dFO��q��la��ˁ-�DN<)^����c��H�N(;}o�3�fZ&��m���w�B[0���%��|t����2 j2�v�L-F_2�����f����RF������������[����1G�b��B*�+�AS����A�[�^6���K0(�\-@ٔdK#,��Hq*��Pm��������X�̈́���9Q��^@N|�Ω�:]�i�u���ύ�qU"DH�ó�/�EUj���^sN_ǁ�����,����j?=����r��L�؀)1Z_��ф��C�˙/x|�m�/I8G�\S� ��bN1�MT�� �L�Է!��Ra��p�)�F�ڪ^�;�޺�$�d4�:�K_@XֶoQ)����n���Y�0�[M+�F?��QK���7���n�{j���.V�Τ?�hWԧ�K���G�������7_Ī��	�e�r�u�o0�>;c1�;r[İ� �2��p?{g�R�D��N�JI7��@tW,�o¼��(� ��֠J�gs@0��v�\H��z&�%n�NA��~#"낅nW�>��ݣ���HXs���m=}�J���2h��o�Op����eto��3��S4yW����Վ�^� l��w�����5X k��y\��ut'&0y�Z����ޞ:0b���s�^�)�����3��#?Z	��_��h��{���2W���S�"7�ɡ�b��b�.�D#v^!�J���B^c�O��� �j�}�&KD}�����"k<��'�叿l]�d 9䲁�����V̰t�;#���yqՎ�΂�̯��*��+�+V_6�^���hK�Q�1��e,o��o`�E�xC�� XN8�g{4����������ߍ]�O�5�e�[�n0R.U�,e��,ޒ�4���x����J�]_�;R����n�L��o�&�c��ݺ���+F&h�8+T�u@ϒJ��|����m�7��7��|ˈm���=�*sTc����s;�g$u�ppy6�swr�L�yg�
�>l)I��黉�ڦ��Z�7��V�x� ���hc8:GQcs����:ؼuz�3F��8��"�-�; Z�%�p�[��7fzh��(�8�L�*�R���tv�޺/H
s����Ĥ��!Oq�)�f~�&����\v��5+'���+1^���F)50h����|�Qrf!�\�p$���{ZC��}m ����yϮՖ%�2�$�5���x�
�%�Bԙ	-�o�Zؘ�e��(�7���õI["l�E���R{��S)3�U��&��RȃJm���|Z���ww��Ϊr{��nu�w�﫟)^=�����k� ����j|[;ԃN�>M}F�Z�C�,��w��99A:���U𾨩�Ɍ����,�"���O=�[�U�B~� 2�c����ⲗC[�sz��nċ=q$�ڵ��r��"_�*��C����҂��Y��1I�ՃJK�5���]�:E3V�܂��?�� �ufw�7Ϛ�nٳs%ޚ�'q:m�>t|k*pJ��U��>����˂�&+{/$e�Ih�!��5�?'�+� ~��
M�D"G�P	���I	���Q�0ؤ��#���h��kt�_�hQ��\�zp�r������G��!A-��A��xaTB���Leq.:Q}��;�4��~��;��-UX�ٶd����0�/�6�\$d��Ň��;�H}b%����YNχ��8Ƶ!Q�7v6�8㺖� ��;�<��/�B�j��F(�u��"����|_������x��|(�����3M)H���p/�N����W^�-�+��4��I�[���?��jגD�|�Z� �6(l�]�/eJ]$�x�I�&PQ>�#_�cIʽ��'ƈ��/�3=W��-M��7��Q/�J߈:\w�Ho���W����eQ����������ꉼ��Ͽ�=�S�ml�ӵ�X �5����,qߨ�N�>aW��]���� W2�a�+�����G���EeO�U&��ѻjأ�|!+ �;��O����ǃ��!}�z�]�K��Xb#M�Y�!|�ş �sv$����}�$)#��:� 1~ђ����{���c���^Vq�L���"���)����T�<���M���t�?����qP��B�`{�_~��3��9~�Ђ���;�E�{��t({�W@ ?z����[���\�s�p+��OZ�rf�`�W��.'@��^����Ize���}����iT�q:���hV�p����\�p�I�7w��m������}(l�/����:!�k�,�qM�CNel/�x"�R=98쏡�0��8�OV�G��>D2�!co��ǜ��d �Ψ�v!J���X��)�Uu�"���;�p���!�p6��k���`|q� b�z���b��ªc��-��B ���;L���ٽo��v6{E)q(�����p�}PE�)�}f �;�q����W�+Z
[*�)�#��1��A[}q	+�8x�k������-9���,�l�.���y��'w[&���n�8z��N*fh�Kr����̈́�g ���}�5h������o��Ŵ����;Q�(7þx���3 Kڽ:�D�y`�����]k_��NW� 
I���N�}\�ޯ��&�=�
M���[���G�hS l�5�� ��5�w��So�Ȩ$䶮���q���r���[�Ȫ�J*���L�q�D+����b��Ru��m�A�� �bW�{��5	z�C�" ��ؾ��kkG��.�i 9fa�B����4k�TPI�֌�EFɼ���1#KԍP�s���b�<��m9Vt�_��9,�$K�D�D��x��v6R,�����D�r�dO�4�ճ�D./�I�B�h��soI9�k L�*�\ήC%�FM�3�%x�9 %%����Ē�"��h��#E�b�m���Vx�@��Hn��V������#oc䘬���C_�K9	">O��91>a��{�p4�y2�މ���N�\穜�ʠ	����A�����B����N��D��
F��A���|�U�|0!&c	�7b�:�"�K�FO0��p��j&����a��sc/#m����;e	L�>���!W+h��E{ _�i	+�Tg��j�@2��f�	�����%uM���޸��ӆ�Wa3��؜�Md�<X����pϸRr}�1�ԑQ��LZb0� �\Z !��?�o��C"�ғc���r�)u(qF%
ȣ�	���z�C�U(�VN�BC�.'"c5!�|o���G�[���4���W�Y�M(?مe�"ȾH�Nx����j�"�.C��M@H~�u=�B���E�	=��[�.:7�7�*8�Z�M��`1�4,��[�c���z֛�yw����ۧ��{L�V��U#
m�o�����������ž���m�?��>w4)���Z0�[0FԿ������4'*�1Z/Ύ��~��O���,Q+�A�\w��|��P�]�e�Z�B�(b��䮚�r,K �z�e�P��O����B�_&�O��]d�C@l���@\�-��u�)�7��L�!V�,s�\~�{ǃ�*�cd/c�8忀� .n�sM`�t��./�-�P�u�����;נ����dAң|�g��&�qŰ)&�Gl�Q�-f
x#b& X箭{�%��чwޜ�{�����$�?o�w�� �
�e��*C�ȯ�ݝ�J�P>eԵ���<�c�Ug>U� >��0�i}�Ѯ�k�m}���:}�g�{�����w�:��Zܺ>8�����Р��ĺ��3��T5�s?N���ф�$��fG�98�7�K��Qu�>c�� !i�U�*	�dtK�n�n���i%Yt���~O~�j
ЩgOFC��M���m�c�5��+���X���l��y��3ipShx<�w<9�ʶ$d6��Ku�$:�w/���H$B�]����|��[��8�s���Pw���$�δd�'h�!�r}�#�p�:$�ْ��L�jPUs�ʕ����S<�ό�j�Tv�IO�WT�h�����rWnG�)�zu�C����A[��u���̢l9��äq�np'�\IkD�8J	Hr\i��P)Ѹ�:�k��O�°ђu� Tƞ�u����^�BW��~�Xr����f���Q萅	����dva�BW�W��<���2���r�t��:��c�_O%X���Y}��[��֠�%d�>B��Ll�5B/�����Ϛ�O!�C:�Cq�l{��D��+�\�>�w3�7���8����v?T]kj;)���Ot����~ɐ�i_ 1h=wӚ��r�Ty���-ֶN4J�ݍD,Мay���د?�n����_�]@�V+�Ǻ3J�b�q����)B���8]�ם;�V,K`\���J;e��$xs�Z��rFK
k��BZ��U����a�<���FA�`W�P���呰O8�|R,fS�z�yw�;���u���*���~�:ɣ5�v� ��%u�]Ƞ��8����ϝu	8�c$��74�KEo��6�^��w?Fnd�ɑ=A�ô����|yVkju#�|�XUs\�4g����� �3>��㝛#h�۬�qΡW,��ɱ�����:`ʀ��9��L<�7l��CP\����q��_��a?���\%0��������	'.��j�f�	��MӠ��%(/�UW.S���c����?W@��{��A�~$	Z�9�{8-P��(��GwE�iʆD��<��5�zX;E��is~{PX�rg@����u9�1;d-/s:?K��H��&A�.s:v,�e}�6���/ܚ8�J FG_xI ���N"���Q	��D� @l���(`뀭�4�`#cH�&g?K�7GLl�:���8�`J.��Z�z�UZCS��R�7xe�lQڸ�R���A\�_�?vƭ/�{�m(K���3}�kS���=복�D!/��3��ȹ�]e4�*�,���c#�<2�iІ2о���E�v��?n:�)X��_�]�jsIɥJ����z}��QO�3�7Q�$�߅��H��m#Ȣ� -7�S����e��L->����x�-A�*����9o���bM������"A^���l����S�n����N�����ŶmE�K_n�A���J623-����_X4�>��Q��ã���Y5�fǅX̏�*8r�hU���ďϿ����>����*��F��u	�9�[T�o�M<����N�n�s�J]���swU��\ �M�D2������ ;��4U*{Ϩ�T�bjǯ��W��h��G��
L?�g����YUDúh�,9����Ӹ'���T�ޕ�t�[�Ɨ$��0�M%I�đ�8]Y�Zӄ)�X��|ǚl���QR=��-��X#Gj��҃�L�����&�*	�Ƃ��3?�[ii��K��ZM��hR@6�����P���d��.hg�$�'���m��å`v='�T��	��Y���!b�fv0���<�1��7�$G*������ЖG�zu��R�ǯ��66�꣄+�F6b���क़SD��k�H��j<�9�p�����+�Rw���8�J0a �gc�!Kz7��k ��o��-��)t�%������2�\�އ_^��j?SY�lF	z���-X ��ݬ�y��UR��t�^L*�"�`Z��ѓ��fCh��Gȥ:Ahg��V��~B`_*تoeC$cW�������+Ux�^�g͢�@��͡C��nt��ۃ��k�z������TD� ֧?�����k�,w<�]�z�Ty�5���saz�ʪ:�L0֯����4�U��k�M��WE��f*`8BER\��KYȯ����>�H�7[Um�AMO��0��ɋ��V��;P�P��Qs�]z8����+� /��GU�
PQ�� ��T��]�ձ�?��2��h�Y^	5�.�G�C�)���oNΩH�8��D>�zo�[e�0��U�
l�"�Ngn��s�?��}-��WߨSm�\B��y���&^��.��<�ׄj�пR��/��s���@ �D!�^N�h��i�1��=+�������B����;��Z������A��%�j�`,��zq�3�A�B���K�fJ�z��gb&	x��5B'T1 NP
X�;��\|��|�����ԓs�oH�QՍ«j���rI�g��$�PI�?� _8�O���_|%�

�X��� ڷf?R��w�ȸ��P�r��C�B�v�Ӂ@�����K �B~h���ob��cO�	\Ɠ��FhUm�J��a��#�J!�SYW,}{�$I���3^���:��| �C_�6�����	��5�u.O�h��6�ph�/��ҩǢE��ۺ#�ʭ�vwc9�N˺W[r��:E�J�pZp�smp�@�-������ig�{
�IjH=5Q�$r��R���l��y�0�,(ۊ����Fϓ�i��_49����l�c$H��X���[��p���BD�u���<Az��R�˷�"X�[d�@X��fݦ��@�� L�\+W��;�j��8j��2��0`�I��&S�r��.9�����ǉ�������8�<���cm��N��v�
���-ߞY��z�s�Xh�������A�ܣ/
�������棝�N:��%� �b��јg_<���֛��������d=�ȶh#׼k��� �q����cv�;:� 9WvV(��M
���!P��� ���L�3a��%�<��le��$�(�5r��*�ݭ�<�GV��|� y���> &,k~'im~�~17/�C�^�t�IYqk�Um噘�������`��yMh5�f��@�h�wM�56�i��ṑc�W��[
S��9N�tC>��3������q2�E��Tf[On���*Oך�~T.~�~��q���g�Qɦ���=wB(�����3b��o�\���̹��!�0�0]|%r�#4_���R������O�pG<�7��h$�������ǉ|�"R����k����c�W�7E�1�h�����T�"���W��'�l�-z@Ѻ�c�hS�t����4gPĖ>Ta�RFT��Z�E��ꄗ�����9����<M4�!�P�Eq`= �x�|�{��N���$�� �aX��O�����) N��i"���T4�T�I�Q5&�˃_9�������!n/-],<4�C��?��r4QR#��R�.=3T,�MA�܋V9���R$�&#�E�|)2��P��T���Mٟ][�����e�'ʿ�θ�FР�n�7���(s�S?�r�vrvS���M� ����$���w % �	Kz_�?ZJ���}#Չ�3��B�Ԇ�m  ��O�(q�վp�h��A���T@rmy�S�ӗ�<>�l�s�}�U��� �Ni�a_,V�	o>��f^5��͒�\��J��eIH/[
߻��_>��Fh����W�FG�wI�^���b�"��c⻣�����1LEf��߰*�Ҫ�]�Ӡ"�ZGO���Mj������\LL��E�%�ygj����d�
9&�!��Q��Bv�ٮ̄I]���$��[ٚ�&�#.�5��f�#�@J�W�>(��:W9*�VFk7=�ɴ=g��v�=��t�d�:��I��\<q���[�������;�43�%� s���ב<c|�AL�JSCh>�OO���w��Z�V|��X���z.ɡ�wB)-�Y��,1�&N�4�ln�qؚ!8��sN��b�dS�ר�k���XC�#
��C���M�нz�;	�K��[���	��o�	�A0��ۑ�4����u ����]\鬠>ΩWDa��-?z�o�o�p�/qt���rm�9PL7�^Oq���/���g3�"c�)h:����Q��}�K����~~S��c�{w�KY�Xn�������?�Δ)�gb��n��z>�],�H[��"��c�p�b�&�!U�☂�@y�8\B�7�l�q���g��}���L�n����˯T�����IzŶ��q'm��>@m���lQ�1�:F�[i�B�$4��mH��k��#�gl�ǨI@Ȳ�h�{	�0/�/����Ƃ�"7I��eM��)\J���}���@/f��LҠ��I*(z�|o�#Q��K��q�'��k�o������Z��/?!\Gpa�5'b��H��0Ӻ7����Q�oɩLP7Md�Z��ЭO�>6���*v��p��6h�F�m���	��Qs�~4NIVrۓ0Ϫ9#]
7��{��ᆝ�����$�]�#~җez�@�xf��Af�ކ�(5��&�~t�wM��Za/S4�͹��R����õ���A�$��y h�n4�A�g|г��L��*%�WA[	X�OK$!�4����HHu=#�1���oP|N	��뒑Ռtp=H�ҋ�t��!8̳?NJ6ኈ���)*�q��o�I];
Kv۶�Γ�Hf�x�����
�T��#
������?�����N�^Ȝ���}4�^���a��|�v�d���rj��;ҫ�e�i� ��#AqZƿ�ٲ�w�������O�G�+'C�a|�Z:-)2f�����[�9�?���J�0�C�Std�<G�>��0m�>��ٵ�uF�{���3ve�Ax��c^h\�Ә[��H�F��樶�Vo%�E������1���`�ᨊR����kQ<L񼢉7'j6�#H���&�'��"ɣ���R+�~�+�ݾ����!�w�N�&����k��������cHG�Q|��&�*ޒ��l�y�x`B�P��k�4��L�J.IvRn�n�&�W�w�C��y��.���:g��[Ǚ@��W7.z/,+y,n腟dN��v<�8�gΩ�o�m��+$� $'|I�X	T�؜i��ӼcMQ{ ��T�+.)Jj�D8�M\���7�C��v��E�h��>X�}xٜlR�(,�[knW�/^�N=�I�
���П/�w��L6C.�UX��z���ҧ�4>��P"Qu�eK-E�6:km���� 0-uvRԀ0=������@)����| ��x�Q/6e�M���R9$!������$ �XvH�	�Ќ����0Vw�A�8i�.��C��Y�E�jO5J�cH[N�/��Lp�N+�E�x���0�K}l���b{{Է:1���_p�}��)�G�U��C/<���R4�)O�#�'�QR�4	����i7 ��f�B���K84| :w�r�r}�`ܛ��ͱ�3�����j��ܨܟA��"��1t����I�m���:0�C����?�JJ�F�t˯#��e�U�硛���,h��
F�Z�ݜ�H	�xX�ΟvT:E����&Z�l���_n�B�[�>7���S"e��L�A�8�G7$�Ap�Z>6N����1�2�-����[�N�b6��΃��3���j:�0��?.���s�m�L>%�C^��J5�<��V��H��s�ucw͐��Ҍ�o%�>�j�Tj`@ʍVi�6~���4kG�}�nKqO�:;{#<r��'?󁿣��]�����P�؃$���g�|�ԋV��f�f���Y�ۆ��|�^#���5F��jo�u�s�N�:�x�ہdk�m�u{��SbM�٠�z6����g�@�wm��E����[U����C0��F6KCq�C�gg/�O��*�"0L��ɯ &ɋ�kU�ҨG��A�7Y��U�{R+�C���s��;��B��էI$�Ms%�<9�~<�mx����6�6�Q�w�V��ҰM�p�%BwŢεN����Q�S�$8���W�w��n"S��4�VNj��dȃ��1l��� �B�<�uQ�eC�r�;�wN����8�7��ї��RT���H����N^�g�
��h�T!����M�gw��VK�=hR'�Q��"lU�-�b��ؤ���Ĕ��H�?D[w��#Z�Uk�������i�`���� �k#�R�}1�=?�\X�Fė3���^_�#e�rT�bkt���
�����Tn?"�d�ty��P���Tg���)�|�a�X��?(���5�����b��ρ��#C�螠Twr�{c��R�|m���_$l���'?_�,|2�����wv��ƥ����O"����x�X�qL%Ow������-�sf1t���z>�V%�8*cua��i��R�@�:�y�q�rM�;u���Uj�V�a������P�Hnv������fy�C^P��gB�H�c���ک�Q�xW����^j\Y�� ��4=��ZJӂ�iJ���L��Gz���J�G������� ��;qP�0X�����*9�/,����w�.3·�_���f�r�H�7���L�~s"Ts�Gh��/I�}�V��)��MIt�N�?1��r�wj��f�Rzc�y�n��'Q��A���(�9��]ܖ��X��]4_i*���Y��8☆0_�,��ӗ�/�Z�Bq�4�疳4�M����H���9�ߎ~d�M��|���T�,�'u��n��S��"�0�=R�2�*�n���}����«a�G<��u����s3w�w4�����
3�շ�n=�gfMLEf�c�
r0�8��P����g��dr�ބ t�<��C*S��Tf�|Eh�����dA��( ���v�CR�Pi�э���[plo[9��qJr� ��E�����ȧ��c��ז��q�5%*�[ >��5�Y[�@O3ƥ�˛*_i���&�,�J�S��}��1b._Rh-�3z�hEԿ��%���1au��d\8��9˯1��1��Zf��Pȝq��&w��	�fL�E�D1�k*��ECP�̖��줇�h
�٧~�
Ģsy��p|�vO�"{4��~K�)e,��ץCD+'���:|�#H�.��]��?�����⭡�b���8v�`�[��,�fwc�L�s}�y�ʞ�3�u�@��jF����q�c�ˮ�:*T�� �c�\O���43�jG�\��	`6h�r-(������p�h�+���C���Wl�B���պf�N�)I��S����Ӛ��)�V�t"����)R���m�8�x�61y�8�#�O�����D��tˎ�0O���xڥ��d��.%��(��İ��&,�N������|*2��g�(�Q��]'����2��� ��t�P'��S��mtM0�l��;�h@Z^	�F\�tZt~9��+G��|)A�J�',�ix��!�`f��24�[Q@(Yy��N�{Lʘ�䗥\/jc��	x^b���/ZLr������`q�ˎ$W�=�������C�&yj�����"A~�r\/��	%�Փ6<� �Աyo`:j�̑>z3��Ϳ��ޖ"|t���R��l��o�C]����9���D'�,�xـʛ{�n<��OV����A�_�l��gەF����C<����˃c*�X�t�A�M�64�/���h����~o?��|�K��x7*:���"���*�y�nF�n��%�΅l���o���HL:M����6!*�)�z6��S���P�G<>�w��V]�n���:ﶉe��s���&��,�5����~|�������]���O��r�~W�bG���.�f��PB���WMxa�13e��`�Ӽ�S��=dY� 0���AB���S�3׾�d�Y�g�o_�5E`?!��(����I���;��DMȮ��߷Ǣd�p4�#�q�~P'DQ2Kdp��aݾ�F��&E��hP�{2K��~�q�gF�vJӋ������W_��˒�u'rGc�Z5G�b"�J�(�;
i�Ш�t���a�Z	�m �^�����i����N͑�Y�~��˪��'�0Td&�-����R���C�7�G�#�b����u�zߒ�i$}O��b���GI[}6NY�nm#�|�G,ó�*3 �4��6{rM��Ɩc�^ ���**��h={i�W�sþ���-5��^@�F��zZ�F���5�r`oV\��p4;��5�E�����8�b`
� ��U�{J���^d�D��[¿@{�'�r~��?%���ק�]F�Gwg���$/�[�2��bvS:�l�ؿqL��Ow0�4��$��*ʳEGV4�E:!�4�tn�13 �	F�Y�� J_��P�X\r�0����@si�����D�j�n��5/&|�.�k�`���@���DD���K1�:����[�q�����#b6��,��:��bo9�`���M�r�Md���,ؓ�FQ����!y끣�9#���}s���_ݕhf�L�#�8��UΫ�6/�JD���f��*ʃ%� UUȹ�:�GJ7F�Fj��<��A��:H�s|:H�#�H��<#;	�#B5sQ�A$�Yޞ���4{�"���|V�D:�yt>"ސ���X!Q='j��8��s]�
?�8�4>^��n%�z�@uOiSUY�Go�S��0�S�U���pl@�e���Q�l5����.��<E�eZB�#��;��p~�g��"[�/Ey
a��ɨR�݌��!y":�l���T���]OI�ґZ�3��a��Z=� ���_���]��q��;7�H��
^/!������@��ro�K��>�- lTd��=�Y�#L��6z�t \�N�zFP�/�M�s��GqpW��{���'�x൓Aq�)N|�?� �@֠ý�ȼ�f@B��R������A��/�d2���K0x�s�u��� ���"=��.���2p�ŷ'wv�a֨uzS�,��~.�~��:�0W�l&$��V��n�p����8��0�p|�	�R��ӕ�'��r{��@���M�WJe
K�jh?)���@�h�k�0�\H=`�u���?�Ũ�:ˑ2qn�0�E�p��1�"�
gyY�YtK����9S{ �b�V IY<�h?��|�y�\�(��¡܀E4&��ϯ��(�'����q�� ���7<[�Ԗjɑ�I�`K�؎�ą�=�|�E�lݏ6v�g؝�6���2��fA�+��*��
���Fw�A(H �������3a\VQmu��I�uiv�af$�mVa�-*`��|u�%7�����sR�aa##�Xo[�:��Fwg���52��>~Y֚�4R4L�2(�F�[��\	[#��$evX�{=����w���G��� �u{[����� 6��_R�D�|��?�ٲ��פ}�<ygQ5�3�����n�s�1���W����	�×`C���tT�"�
`Y����G���}���Y�� ^�cl�K���&�6��'`~'M�?8���,,��*ydP�,_�3�Gj��#�]^Z<6s)�L��Æ��~?�(�r�.�OÕLW߬+ �ҹr���M���
�J�����c7m��D�0�����$|q����qb�zZ�n?'�,�S2S����%i�)�pZZ+�"�g��B�dnC��^S~�Ў�9.��k�F�`�u���V<�>�GCЪ��m~+� 9]���h��h~���#��[:/����|rq�S���$&��G��������'�QW;맢��D��fCcn���sd���K�:���?�?� 1D�K� 
"?M�T
:��kK��XBlJ#�u�^R'%�E�pW�戢���c��Oi��O�ߵ�a%r�h���o,C����̱S!A�+W�_�$E�37�<iC��M&\�{�$��	��9Iu^1v�6"�w�iHE���	��l�]1�JKT��w:�JQL>ǅh� y=��0��]ʸf}�2?�w�&��?�[���ɷR�J���O�V�ؕ�P���8���Y����C��co/�
=�2�?m�c8�����x.�NoXA��Z��o��|��YXg�O��D*���ᾝ���}VH�(|����N����1��k����ɀF�P-=A�ajx/ο�S����r�#_���n�f6�Q����i� C��U~��r�Şs���Xݞ��S�e��ALE��*��ki����sLf��Ň5^�WL��dd�s�������T$��CjW���b}
T<�p��q%>�d�o�#�z�~)"��ĝ�Tg튖:�rS�h#�~�Մ�1 A�M�(���n��rc>VG ���H�U
zfٴj�G^o��r�2\�m����|X=��Sq��� eA��:��gr,V@X
�h�4"&z�
�a��&��{[�ܛ�.\�3�)R��E��ƍ;�#b�f�L�x
�SS	�.�8���]��s�r�%�%n�1��'��i�98�ܾc ��~a}�;�L-���+��w9�yƮgM5?)���Ʊ��[��cf¬:�O$ @PC�O4<qk 6kh����#�gՅ��"�	RE�m<�/���ڀd�<�sUʗ�=�T�
���_����))�r�mj��R7�½��ڨp[�e�7h4|mpϟ����8�xKB�6�M�Lط�Vb��WDڊ��V}@ &��00��S8��b��|�g��&W��5���1�����G3K��p�1$Tj� �gu�S�$ڶ���9]�����'��Wʟ4`��ٳ�g�0����y�[r}��@���6>.��j�n�a[��J�Q��3{�w�"T~�ek���<�_5���B��B�r��.���V:	�k�=7�&�yƩ'�s���&$��=$�`֥re���ͪ-�����R���dr�x/]��\{>�s�|�V1.|�c�AH�w�ǋրZ���`�R+�[
�@�%4� �eG�vO׎����&ai��R���1~؎�Eɷ��?z���Y͛����`b�$����oQѨe�)�� ����8��~�vL"3��L�Ah�]p͙�r%�<X�S���U�g���"�!�"�o��6��Bi:��_�IP[�p�o����j
)
�?c'��H��9���N ,]�����Ζ>��qY�髭��#"E%�T�9��.`�Jz��=��b_T�	��ƪ��s1
���6m`��	eܹ�1!*el��l�p�(�_��یuPߩ�R�
W�����s�NҘ_�x�:k"D@���_s��?+�Z��y��h��ԈH�x4��(�����d������Q��ǐy �{�m;	Y��@�6�Ϝ�M�����apF�&�{wP�f�R���K�À�u���'N0�*M�Nv��)*�-�4Z�2��ھ��E����/�ݭ�SY�i���P�&TA7������R�E֫�-]K�QS��s�� (�z?�7��/=�@��&�a�`{Ssz��%�,桜��$#��Y�����ԙ�j9w_���6���{��2�}���h`-������A֏=��p [�@�T��&�M?L}��d�|�}Y�}t�A_X��lQ�|���d�0gwKT��-��8���bͤ	r�+Q\���p��M��'r}�ن6�1G� �w|�M�(���t�O��G� i���
B����1��{x�h��>�z�n�����~f9\���~�R��G Z�Ckſ�HA��BiP��ƞBj����P���e]�3�> 4'�B1h�$>!HZ���*g���E�C�^R�%�@��-� ���/��)�s���qg�d��e�32z��d�T��`��ex�5r��`l�W������$�X�٬%��1
��[��:�����T\�bƛt�[D�m�)�eAc^R1�,	��U,ڷ�a���tfv�@"���2�G�Ր�}��SW�h�T��ZCo���?�!�J�Q�^e-�Op�5D�G��פٞ ��<<�8fq�n�4���L	^˂�2z�R� �a�IF�7���]3���O?Ɣ\���>���]�k�>ԺT�P3�7)i�V��;�O����䥂1>م�B�/2�y����?�c�;#4u��\!��7�)I��)��Yb�^+#���ҳ����h�0ub��Z��g("�;��ǿ^Y1dV�Ξ::ӆ��r��Wq�u��I_$��@�(����pIDmps`᫱t�.��s�
��On��:���s���?��^f�2<��i�e��Ж/�)�f�Xn��G ���Տ��%A�bH��QVF۷�!#�y�[��f��]�uO�����_���p�t*�|�W���1 �=p�k6�e�ޥ\��%�5,�c
～92��};[����f�b��M�� W��o�u���@�3��{G�A�W��cK׶��V�ϙ�l���+�����8��0K������nQ�<�o0�i��6�Y��c��ۄ��$ɨ��7����ƷLA�r�U��u,���S� F(xJ�p&Adl�(s�:��9?�o���n�eZ�;���fL"�Ĕ�}��Ѭh��ٍ+4�	����oBg��)Qv���w5�͎p7��]d�`jn��R���M�q�v���(}�����"���Y/U���s1bw�;��29:;`>��̐����ẈwUݦH���1�{�,ݩ�.B��3�^�&����~bOIg����������T�B�S�G�i�2`�sE�&�M^:9��^SԪ��_R݌��y���j�C<F�@F�-�m�[���|B����W��Gx��fB.34���Έ�Z�K_��g&�$*J�H�]f��Y%�xGEE|UR�ZǞ��:�e�J��9�\{@�`�Ml��z�h�h�!z~��~�V�{\����>�m��s��������0,x��?�Qb�9�B5���-R2���]�y�Xc���!��:��nF���4ub��A�PܙOװh�5�Cb��,Q}�^c��3���i����Z��M��&z�%>�=Ypw���q�b8�%�8�ɔ���U�S�p��� C�Ϝ��`���[΢J�S�ږ%�l�0���|Th�[X<��=�R��7�ӻ�xj��A����P|��B���'zU�1�ї/�z�#vJ�kٲ��"�E)�9���rˇ��:^���	�8m����
%z3�p������{��g�Ћ���	}��h
�At�+s��l���r���n�eQ9����wT݈���re X$A���$s�d���!��:]7��Ԅ8�ߒ��6�I�$����$�#��V~s]6���Q8Vk�YH��þU�(�$�`o�)�ᢤ�M��z�v�c<��з�p�/[�&�'gcoqm���t�:�@��G�9�j{[N>5ۍ�_xs)����řMo\7M�2�w#/J8}$�Ek#�v��#�U	�{�!��{�]ō?#��l:q��Y�(Vdq��)*ψ;�V�E�:�>��ҾP�(��b#��+�}���w��v6|�7Y��Vu��އ���_�y㴚o��
����9�:�/��9��3-zL������H�.��x_ ���#D��$R(v^�Y%M�'Y��^-G:7���7r�)>ڠWE�iHI��D%Tg�Ɉ�c˨���Fd���26����g���3i�e�4xFt�$�'�H����a]T�A��#x?��r{m��w{n�S��I[�C,\�|�+���#ܖ��� �T�q���RMy��&y�*G���e��1|���#?�-��E�+!�uh��E�E�K�����b��=!(<�Qrn���=��|���9	=ā�s�oL�JԨ�(��l������De8�>%��v��t�l����u s�BJ#:��>L�8#@�'dtT�7��oL&p¬j�@u@l�n�9U�4E �+�!�WX3?GKu��pr�͔���r�?=P����.9�[����<�>h�-�!����*>�p�A'H�f!�U�f��mjĵ��l���|��W�O�K�.\ඍZ��p�N� n|���]K������<	��͠�6㆕	/�o�����%��.f^h)!C�s�W��K��Ͷv����-5��U�r��eWg�e�$n[�zzY��m�5q���	6=k�@�����Sd�ܠ3,mԟ'.@�Y�n�'%3x\`�P�:$� ً�L*F�E��A�ߝ^�cL��(|;Y�E��rq��\ũV��"��:FZ��w4C%29��S�&�o�my�*��Gk��°��RF��_�7�Z�zomI��2����`h�9V�P���Zr)�?�˲C��g��9�v�pCDD�� i�HO��c�I�UeL�.�<�
�Fb��t
�v�'��R1�T������zo1��p�*k���o4����'����RX��<a2�\ζ&��ՁO�>: 2����nCK�&t�������o���.���ρ��.!>	{�F˭��
�K���nF��q�� kP::E��d���2�~�w $�<�@q�i��]�7��ˍqx�͒Ԫ�'��>��(}g�8�L�s�Ì\��r�ص�n��Wgb���m&ve���.�L� �xq��{C�o��k�+�Z�!LSJXj��D�v`Af�+V���^���$EŰ��Y�<v|��g��j])]�XR�RBs��]]cpi�Qv�w;
���S'���J�y�=��O6�~H��ux�Ѣۨ|��,�v�#c`�"@��]1NU�k������Ė�d�uէ0�$�_0�)y�)�Yr�E���u�q���3�=��<��{����?�t�����;��5R�2����p�z7���c$3����H�m���	.�
;>�s���d������ �Ӊ�5T��و��J/�N;�����\�@�)�opW��Ovj��7�߬��W��[����1�n
Q9lD�� �������R%/.u ��4��x��:�&��Ű=j	�����{#��2��Db��7�ǩ��~�%w���!f�!uyq�x���I*����@'��D�� ���8��jD�?�lM)�,��T���Ԗ&z=ۨ��eǥ���͒X7:�EE3w�duY�p�J�e��%��Y�h��!{�@_:�չ3���lƒ�η���?�ˤ��+5c�vh@�1js���X��>���}t�/��s�
��z�Kd�W- �P�p���jC�E���)n/�F`P�l��*v�.ݯ�qv̿R��IF���ýӉr�(�A��`�� ��
��ǌN2��O4������$z �7h�����.iY���5U�O�����w���2C�1t��	��ycA�ov���α�hw���'������Y�'-��n�9x��c�Y\�L"��g���}�f�Z�鲁�����Ԍ��i�0?a�F����:m�iƽ;e'V�X�EiK���4���	�p���t�%S�R?NP���� D�HA�q��	6
ŜHt^���?˥��ԦYc��Q�|�ɺ��)������F�qj��gQt�c�
�g�&x�F�q��N�-5e��rA�	��މ�)���S���������H���D$���|�7
�I���e�ɦ�*\Oî��1,�y�c~������ڬxw#����V,��r<�\[�U�;�t8��cO;���h����g�^�.#�J\�`|����S׆�5�e����w��tx�@�����:�=��+R}M FV��BYTh���1�@�����E9^K��J(�㫗2/cM_{�+'�T��,��=�9���ڞI�R=��'�> ),��0֌�Ե�f��46������t�]|�3R��SR{[�[\�~�o�ۏ8T���;&��;=�IJ�ҩҸ�츤��s^�].�gFBue�oλ�b�)�I	�������!��?��Z0�4������^>JU��)D�����D?�ήWG�/o�x�$p��8��� ���]�&�b#-�"XQ�HH���� �c"ݗ�'KnI�ˬֿ ������i��GPM�5��j�;ɲ��т΀xtY)��%��ܙ)*�-��s<�&Z�z~�o�Lh�8*��x���?�i���g�;ϲ��>ɃnJsk/!d#.��ۓE@Q�?ь�TK0I�܇bG���oۏD�}Q�ݳY��l�ֵ0�� �FrjOO|4����ȷ<z����!�7�	XB�R+������� ��H�`S�K��x�bm��%��ٹ�^M�Y@�QZC�|D�WU�w�������E���C�n�5���9��(����-��k�5 }�to+����E�zQ�b�J���W׋�8�0L�F�n�*h�����[1|܆@8�0Y'�q���tz06O����L��<����討�b�Q�|�7t�Q��Q���� /���m�A�4EX#�N�ڻ]9i��"(�������ݙ�ډ���&>Q.��t�ޔ���697�{�����1����<�ڶ/
6�K�����D��>�0��B��s����$�&�����I��a����{y�k�s�9�ZR�[��J����h��jP2�ܤ!(� �>����������8^�]U:X�t�I%��D���^��l�r�j\���d�qvEx��'��Ht �I�F"B���Qli�����f�X_<G[�WUğwl�4=�s_�Ӗ��Z$55�?��$�u�U�9��	�n�/���A�]��"1#A=�y�,�s����B�n���KH7���Y5OXߌ>�G��q��Ē�R��ƓHJ��Ƥ&;[tr٨i�']��\�t�#��kL3����L���Vm�M��16�EN�y�����U(�6҉j�ak�ѵdRq�fI
�D��Ru��S�]^	�/3�:#ĕ=�������<q��ނZ�D���A��o������	���֏��I�<��#R��&g�;�Kz�1����f	�x���~���Vzy�N��':�=���}D�K�5e(a�M7�Cg���C����E^�֌y�8u�~۞���6��'-ĵ	�Rxڊ�����JG���o�&(*����s�S"$�Jp)��f��/	���D���-�s�J���$\���m["Dw�A7@MNbK���x{[���Ʋ˪]��|v����`s���Oc6��6T�)= �+J�a�yz�x����A����EP���W?�L���|!�����lz%<�n�휣��f�����)N:g#`�?�n��(��o���:/��Q#�����;����S�0�,JBt�[�~���
-+y#͒���>���(�j�p\���|�Y�!K�������Ѡ7�[� �}��Sd��xc�S��C(q�_	��@�|�x��|k���R#1�u��k����T��(}4�D����Q�����ޫt�GABx�u�]k�a�Ņ�$+kIey�%z5�A�p�Rj����$CϨ����y�݀�c�i���XrP��3���>��2H�^����k��e����ظ������Jƾ �Y�màQUƜc?m=p�a2-K� �
�:�,��
�GI�vJf���r%�Q�����Bw;�m_����(��o�^��>e�bIA�Nv�+�VO�2��Әc}�մdc�-~�	���h�PDC�ر�y�?�+:�n?�ıf\�m9-���kx1�ʹ�q?��c��C�3��D���K�������K}�g;?H�	�g�(u�fU3���{@?/���!�D�k�:�Ű��u/�Y .�[v�gU�e(���V�]p.L+�}���I%��<�wR�b	�Fdܱ��)^$��j��{���ٓ�׃��F�J!q��E���I^Q����QS^�m8]S���b� �V�	���f�����B��S �n�9�Ȣ�{u�s	\WfD,w�y�
� f*��D����� c�����;{��6 �(��~�ohl��e�M�*i������Q t���Bmi�^��lmo��Z<^p�Dο�D�r8�=���>�f�l�.w�z�Ab.��̼̩$�{D���ѝg�xџ'��=����T�ǮLL*���vp뾪�޺����TfAR���-祑���x=At����/�G�ʞ���|$SQ`ݩ)FD8�Dk<�I��≌<K�kՕ�9���
M*�� j��9(C���}zPqBh�¶^@p�ƣ��\�J�S��v�eahW �O�tB�;�ޔ<xg�b@r%��;�|�]CEU�BZ�����%�Eb~��ߨ^�|H��E���Q65s�EAa�ƶN�퍑2�M��3�w��?v��W��f��1���=�_�pp�J&ɏ�O%�Xw��������՞��~�򼨼�훻�G掸x�I���w(�����E�C!]|�_�X�5qg�z���޾j�Ug�8��:U���l�؛hѸ��5>+�kKԚ/��-R�BJ4�']kTJ^�}��8����!Ƒ�H9����a㠾C�Z��[��uJ�ll�Y�)�ؐr8v�ݟt�e�*߭T<���qNf��F\��'���Q��mr&,2�v�Ŕ�i����� Ǘ.���N>�n�wVA�Å��G���e���!5�ݮ�7;�c�2�p�&�tf�/Br6J���I��n�D�u�ܶ=�N���0���N.a�'(����f#[���۞*��+y�%�'�N��q0*$<s��[q�5���8�,����n�]{�a���A��{ۤM�N'M5{�Zs�V�Z?ap�-�'ｴ�f��7��55G��ȉ���iB16�~��	:l��-���s��*ސ 0�7a]r#��`+��	c��~�k�+X�����GN/b��-j?�T�&�Ɩ��~�����o_���OI�NF_��C|�֬0Y+����3��/xZ)'x��´��B�d0W��N���eN���9�ӌ�ht��_B�f���]۱�r��w�u^�'��`j*��.����>Jn��6^��8m�Rn
�*�
V #0�/��c�&��v��$"�!���d8p��)!?�ɟ�̙��BP)E�ȡTJ��U�é���l0�"26����?�URf�=���}S�#�	�n<x5���d��(st����L 0�N����6���n;6�"@���~8��U|*�R�{Ж��yc���s�}$`�Ҝ̧k�]�֎IQj�ܗ��V�V7�����^֙�`c;`�ͿT�5��������P,���7l�i���a̋/�N��c����D�|y܍?Ჱ��d��>���|S���r*Ō�cX��O��w�,e�c��6�ԡ�\$�o��6�F�/g;�Ζ���%|?��oBϪ��&uSIlŅ���s&����˙���BK\i���ߜ�gP�}��X{_��ܖ�5�2ޤ��Q
��+z
B��
j|.�d>ӖL����3.}��2;Y���A�7�O���M������1���
�B�ކ#�\^�����)�,���z�#�ڄ�Nh�rq]	ȥ�Ǭ���`���$x1������4�8r*hZ%�n	'���Q�)�k>@iPL
 7���)�t9kW+!��kj�|�H�Y'�{3��opH�l��>�X�3����*��V�$�6J��Z <�F��V~�~�%V�=
�NgYI����{p<L�<~���/�߃e/"�nI��K5�u)0�g�L!�ɛ�u��@,�r0��I�����AB}�@
a�]no��nr�N�^㖪݉���|���	�
4��Z�'[=̙a�l 6O�'�8�߼EQ�b=V`�L�w#��z���-TVB ��e�X*�L���#/)�T���0C��EK|"��	�ht���z[����
�N��іЊC`V��f���VQ�WZ��_����lv������#�9.\|I�!"�&����wu.��R�1̆!��b�l��k�'��6��P��|9��P����$�x���{��8�V����XӴ���&&����`OU���[äO=@�B��m#/v40y/$?�>?���<�v�9I%������y>���4H��V�4��e��z���x�AV�1�3�/`Pw�J��|��Q0��~�c�@�}U���]N���$n���2a�qڈ�3V+eqmM�M��Me�g�ʇ�X�~w����L�b[
(Qϊ�
��'���ЍS�J���e���uc�y����
c��`.Э��� `����Ƣ�g�Z�*b�i�h~TJW�(;�}�*�zu�����QC;���ŭ������ఴ)�,ؚ����{��ü����Ij����:�N5U��*�W�*�)/��6l񬪽�F�9�d�ͱ<~(H�{���.^����Ί_� ��%p�K�L�xN��?�-�W�P�.θ@ٰ��f�4��$u�ӏ�>��"4��@W
�\�^f�;��0����-?*�e�Vf���I�y%���*��m9|Gk�p'��Ő� ����̔��lhӹ���	o������{���'���A�Hv���TX[�X��X̆e����ܦ�T� ��!F���a�cuҀ6�Y���\�A!�}9>nb��2�v#��Պ���b� m�R�z��r�>zͨ�y����Sȱe�%?�ě����tj)UC:�����-������:
��D-���S��C���;��a�D����83�������_w?T=(~��]��q�%d�� `/ɓ����쉩�1"�.��S��K�Q��^(��ޝdh����zh�]�z�>�Ϣ�j���\p?=�w��tL��t�@ԭ�7�*��>s$�Eo�y���9��ՙ�M�u�_�I A�m��"�n�y@���[�0ѷ�����M$��j���͔��̶�:W[�$lPy�D�J�X jᶦ2��A�����l2+rzh*�ظ�k>U�D��Q�|��bua�N �"ug=����6}wW@��^�Ş��V�����(���1���g�\A��<ҥ~��֮|��`8���� ��kV�Z3{�����G����l�v�`�j����\r����rtTD��EAF���̀l۞����GQx%�3&͖��b!�9�g���� �
�Q��)���S����`;z"+�#K9G+TJY��Q
� �������C��/���ٹ��\����l�A�4���Ͳq:7��]Jk���}p�����1� �H}�!tTb��m��"�m��6Z䇃̹I��41�NylUq0�w����V�D�L��Y�PL�-��Ol�LZw�N_�T�l�ФB��rM�@�Q[�1y��]2��{e�ur�Ym0����t\ą廦��-�骍#1��b��2�>���A���2���^d]�r���E`%���ͫ����R�3d<�`�.7#Vf �!h�`O�E0V�9�/���O�_��d����܊��{�zй�%U�f�Ϻ	N7��2��1�B�A�؜i}����ct��Y �(6�p�%�y�6��5j�6�ߨ����<
+ි����dm�8ϰ��|�k� ,���s@�2fg��ƙS�d%�ޔ�q7PեKBG�����Qj�~�s�J,�2�>/+�3H��և�%���C��Ay{7��[F���n�*�=����I����R�v�� ǏZ�V{�L�����OL*[�hM������Dby�-��������+5�G�s$�&��|�_�ʨ��1m1ЈM�����Y�3�RV%�7I}��b���wU	/�4Vۃ���tj��Dhoϫ9?�U[ ��t���p�Pke�鰂h��Ȉ�������mi�&VΠY��CdH����(N�l�a�U��蕌��2.n�p`�8�+����c;By���_�Y�}����m�o��[�n��* X�g>9+w�%�Tp8�F5�VL��w�K�`I�Gfx08�2hP�RCCp���3��u�V=eq�Ik-~4*Y3?1��+�5���Ur8�0>�3�pl䷟���J,�����Ԧހ}�&W��uw�a�P���W� �H=:��Sw|��
*@�Wq-Д!8.���d&��
�uy�!�𹅰���f����{�9}(|p��m�ȓk-��#o��£ԇ��gxuDiS�`���¤O�@'�tB�]��#�h��,n�@��Td��K�Li��v������|�B��p�|��fs�ǅ����F_ٰЄ�S�������:�;��5|�u2=���9.��֭�o=������䰨����<�D��Wx�,��7i%�U��I�b� �,�ژ=��6J�����D8���(-��VF��Al�g���Y�����-b�ܩ���HД�;D��$�K�C>���ѣ�t����F*{��K�6�HN\����H����.�Ke��}tc��g���I��䇶z"�a��0�TT�}?�j/%�$a�[WGǵ���D�x�^L�V���%�N'����Bm {���{D� <d	��R�V&�߯�������$�53E�7`�7��<��"�>�M�%
`G����7r̝���w�I\���[m��k�&D�*~���5�׽n�QJ�/~��V� g�ø9_�4��q����_�h�w��aCv��^���u&�b�RN�<���t�=\Of��8p1�'��$���m6$��r=Qr�QY˦���U#:�y���0w�ŀMxӥЅ��]���8�gO�I|9���U��z���������q�>D��춨�Z��uXDO�U�s�^㳵�m�y����Z�'�YY�V,��ʴ��G�o�ڥ]=)�'C�k�tg��[�9x6z	�Ɲ�S��kO�J�#��S���4LKFHJ���r��f߅꟫D��\�ܗ-���/9W�f#�(<߿N!Mf���s��;�"�)������8m�O�҉�5���Ҙ\P,z����QJ�%JO7���P��R�C����	&��Va �?1m�4���]�(E���%F���5]K/3�v��P��̇q�P�̻P�ɮ+��Hm�d˲��Ԙ�-�"T>���Q���ǰ�>�q�Wg�.�׿+���cѧF@���@�Q��9�y��xD2u"���������QD�b$arVxf�Q���y��G���6�wlG�Y�^��[��		��iV5*�����Ѝ��ȏA+�F�вXT8Y�W?�ޒ�s�����^�~l}��KИ�,{�փQ�a��Fh_t+��8���Py��{���2��i˙3˲��a�0��}TpO�~�ޞ��}�]�1ն�Ϙ�`ɿ�i9�S��WJ�1,�.��#�,|f}轢��1���l��/B�3xub	?_�7��E7;q������B˝l>ť�@9�K�5>
�����ڌ�cHr+[	�M��$�P� �4�ك�a�
�bqiI��m�('7��>���lX�r�O��za|��unK�y�8�Hz�ϗ�'�_�����Vɨ;�o��K���g`~D	H��w�O��ߣ��Լws��9T��������}�j ��Nhw�����o�M�z\�È��ӊab�4(�K"SL��V;���4���Jwr�`��E�X�=�[��͏����=����=Ҳ82r�<Ң9:x�ڳ-�P���W�νԯ0JT.Ը�Msz���_8N֛��]I}vB���8`S�Ҕ Buh��HMo���#U=ޘZ$�o͑we>�ЎC����7X�苢cCw���]����]o_���ӕ���.:u�JX`�5��.��peN讠(480���9v�'�xY���v��}����	��_qVAmM��a!�8��:�	�=%��������b���fQj-W5룾ח�J������h��Ф�K$�L�=*�P�/G�b�(�3l��/�z;�C79�y�� ���UF�4�n]�V�.���,�.:��d^xdT��5�%;5�f�n�(}�8ꠀ!���1<9!C_$ho�G���U��'�*�1�� �h�+CWF0�RhF�_�"��p�
!�\���-�`#�Ԉ+ŬE�sc��J�#O���7�K�.]����&�S�KŖ�3Ey�VF��e����㨼��djZ�v9� DIN�$A{���XN#(Y�
PB
�TFg����՚qy��%)8�f�Q<�c����`�@t�iL��C{j,�1	BF =�2���x�#77��AIB��k�_*Fgz��ة��8 L}�/�L=�y��k�K|		� <"���r��K�u.��=p[�C����=3�*-g��a����G��s0��~-�{?�~?-��:*րS��Y�{�g%�N����:j�g'^��e�!����XѐK���FLF���܂(��E��(��97����
�p�؅6�l&���j��"��&�)S����.ׄ�w_\q'���>�G���L��Ͽ��c���mZY �o;[!��wA�`���0j�z3z�����=�xÉ�G�Q�n����`�#�5�K����+�~�a���4Ձr(��8�=Kg��Q���!��N�*9�I���k�C��Se�*_�l�[�����MG��>|ܥx�ֽ;��2t��y,[	9�um�%e�v|�Ks�-�R]�Sq�����<��2�
x�6_�����ɇh(��4y>��9è�i��y��!�eM9�|��&"6�C��Њ5&Ͳ���`�,�T$���t�b��,S��o������V,.�a��e���9���h��z��P�~�:��35Ҿ���P˃;I[���k[� ����U%%G<{�z*��Sߞ�T{������؍.�9��w��`�8�/��
�a9�#��f%&��oJ��\3z�F�V%���Y��g�/������h�(�$�m[$�^5,�	�kq1�|�6�4 �K�´<���<��nʂߤp�4Q�U@n��N�|��`�9.?��˵+�r�2��s��#�Q o4o���Sf���e���ޚ<�mQ�_�,�ADxT��[���jhT��W��&��$Dˑ���c����BTS
����N�F����oe1�R��a�4���������������5�l�a�i����O���)��i�-��G��u�ǔlT�Z��/��bQ��(���<^d���u4G��B�Sٷ�xah9�S���*����h�|��/�*�f�x>�
�9�$�p j��
�{冏2��<�Kjҷ�3�̊��s��+�p�[�-�Mw['�9�(N#V��WJ}Y�/�}�,nF�F-��YyS`�vtP�s58L��pmƎ0�ҭ���S�:�W:�	Dߠ�B8[�91	�Fh-�p)���-
v>���׶���8���0�n,�V��A�}O��]��/d�*���y�ݜ4&�=��I)�.�_���j�K��%��'?q�#P��F���=����������n���I?�|/��ԯ����pb#�-�):@|���#�(:���b��0����t�I
4��mSۺy��#`H(Uw�d�	9�6X����v�Nh��O�4�߇���p���2M�k
���6{b�ub�p�\uS�k����ÔJ�.`��
�Y[>�8��Kڷx�>�(���Mn������y�9�n��o�-|9\F��F���@���\�w��P�0ɻٜ
�y����B��o6��,����t�M��]|b�j���(�7J=O�?�$���u;+�l#b-0S�%ԧ�C(�
���ς�<�IW
�j��86m�-�T��++μU��Vw"M�E�p�n(��Y�|�����ǆK�~BT.;�a���'!�ֽe����ǿ�k���v�/�E���G-U���@�a�*s|��t b T��J�m"Tn}���D����H�heg:	5<k�F
��4<qpdV..M����BBD,#V�u��p�;󫰲g�V��}	���&���PI	�´����s:��ƒ��7�d/��+6���^RU��>�k����o(�g���ѯŹ�p=R\�~����I�
gӤ*�KSCPA�įB)�T�j������FH�!�=�9���vW0 p���@O�$��{�=F� {k�v�f��U9a�b�D�hޟ`/F�tD�u_��u�_ �<�ڨa$��;�4��J�D�-�0V�k&-�@DvtDE��>c-�yD��0�\��,�4w&���<�߈�c�Q���^Xn���7m�f���T�W|��f�'2��ZA�oJQ�P�k�o ��nM�_
J�>5l%�+X�P���1��]Մb�8@���:�.)�q\:_��g'�<ǭ�𤗱�㠲@����5Hm'IQ[�r�N=*1�6�o�q�+���KSR�����`_'�s^$/���'���.�\i�������V�X�Z7/v��sT	����@�u��yr���Rͪ��h�Q,C�?�<�7}�q�; �\���>9�i���9/N&E-�ALV�X�YTy0t�9��T�۽����>�v��^3��[�J�M��/�����?؍ߚ�S�s?�nd��c9m����.��-W
�o�U[Mg
��f�$N$@r�䚄����RC�<�T����:֮��3��Z�t��Uoe�^�60 3��� �����o���E+n7;/��x@��8vzT6?�����(n�;#��
�+��2��f���e"͎���BC�7-�����1�RU�p�<ٴ�+5���b1�,H��'^Cfi�5Ҩ�v�Q^�GY�.��>@`�v�J���tG��Bja� @��H��[A彝�]�V��c�$��ɚ-Di��ў�'Ǯ���ű;FD���i?=O}�h�q,�n���ӫ�4R�w�0.��EÂYtY��3Fb^�C������ÿh�,8��:I�X-bń.��Q��ߺ��x�����IE{�j�40F+��K%�N�
|t�>%������ML~���]�d��� i$%w��S֠O��Ji9�uK�0���.�����;(�HLo�R��$���$� z=� yӌ��o&���j����e��#d���8�	�D�8+� S�m���CG<zc��K��\;��㍏?i.:�#X�t<���noi&�u���i�ŞH*F"�hgH1�j�9��"yʹQ7��^G��B:�a�ĬƼ��\�L*�-�2�Q>%$e?�o<�d���i*��BnG.y`�� nv���
��e'�8�ɵW'_�C̢G�<�2b�Ņ.]npN=�f�2�i;�p��P����^x-z��f�?���0�sJ,O��Y)�O�j�d��l�,�G$.:��Z6�=��R��A[��WY��OXMV�N��S� R𕾠�x[\y�����[�����NS��Îu�2���^���IG6���ߎS��u��ԢQ��"`�s1�7�������3�s}��z����xg,8�Uܺr��W��?[�����$kD]��~N���AXU�m�0>�d�E�i��(i&��}��xٻl�w'5ٓʟ�Ӹ��T�G"©�w��]D��rB��v�g��7���Z��&��K.W�����N1��s�Q���%U��/"hg$
^<c�/z�H�%������ǇW��Vy <�*��g<�����D�oĒ�C����GƑ��;�~�	ԢQ<�� �5~�R�.�RՌ� �D�@K���%��&��"	6i�'�fT�ޡb|�d�u�k
���Ӧ���È���N�n��C��	��\�m[���4h�IQ*��	5�	)�*��uDZ�aƕJ+(����L\W���uZ��y&i��˩4����r2��"����\.lwd�����@ErN� ����o��؅�GP(�qa�ng 6˞�� =䌌��qU���1�BTz������=�u��F���\�D#�-?=�;f�a�UY@\��߻�c�&A���p�;E]2�D##y����cM�� ��
�`ծ�$���Y	��e	�� H�r"����ڟ8G<K�6xY�y��i����r��j��Z� XY�����<�I���G^���:~��Ĺ���?��$)�ת���^=��r�U��2�-��m�?#�,@D姞���.�oB�-α�Q*r�N�췎�hc�f�0P�^�B�٧���]X�܁�d��as�|sק8ڿ��D�	��BG�5Eyv)����9Vq�@�;i���F�� |��r �y!~7[���J5�'Q�]�ʵ�69�|)�2AJ���R�~���O��R�X�0��
S���z��~Te�%���7a`��J�6�[ɤ7.|�j9+jij6'��o��iD/��s�E�hc�Ȣ����(��,Uh����Uc���_�Z�q��.'��3Yg�c��Z"����-p���c�6�A�4���^��yօ���#%99>	I�`SՃ�s��&u�[ﵲ]̭*�G<���C�T��A�"n��=r��]�����`T �Z���t5.�ē�J���M1� ��b�M����������l����QI�W���}2�9_�k[i%���-�G\�M�	�S?o�Օ�_�,�8H\�R���G��J�翏��Yl�n���.
ͯ���N5	��jN.�8��ff¶Ϩ�bթGt>�pYl�ߗ�I�U��|m��C����<����}*��?�*�+2'|��c w�Z�>�+T^g���Wy��)_6�Ɨ�r�@
ef���/zB����/�m��,*�b�P -���޶ ���w;��o�,}�<Y���,�k�=�35Z�*�泛�|M&�4�x�l��@������[��Źqa7
�+�
;�'5t"߃�H��#>2�?�c������x��-�3��L�'�h�̃a�uoj���'�bW|�]7%<����5>d3&�"�V��}Ɲu)��L� ���d7	w(Gk+�š�H�#_�IR�h�Z��U��e���v�ۑ0Qp�Q�x�x�l���_GT&�?ː;%T.��������^�ɺ��劤/�
�%۔�R��Ap�H��͓�_��/��2v�J7[|�:XQ��/��+t���Û��>�D�ɏ{Z����&��|���8�r���HuL0�;���_�������!�������l��9a�oLsWlW����6-���m�Fd"�Ҕܹ]��QAȊdΏ������>m���^�qB�� y@�n8P���d5��b]�h����S�]�X�.DO����T2T��۪Nw`���`(ns��JM�DQ6�a�X�P��^�{��iPU�I�jߤ���k��u@;���%i~�q� {P?�{����"A�� �ཾ�v��e�c ��Ncr钾ҡ�9O�$�����8Y�I�k�w`�w���t=��{j.@��CW#O!�U�5�#�������j�������n�v�����Tyw�+�sXO��:y�i��̿�^��!,K��Xl6t't��~	��blV��$��&�Fw�W&�����*�;(������e���v�/d�w�h9�@��J�`Ro����$u4�Ii�Y^�t�LK�]qٮj�\���<�f�n�	�ܢlڏ��>�VF��|���~�z�7�n�MT�	j;����|��g��6Duo:��W�oӑ5�p���B����I�N�G2�.���B`����s'���b�8s���%&]:���^�G����"��'ð0�RyU�+}	� �VK�&����ע��ɯ��-�4�q?�A8^b�='���E�Ze[�9&A�49���Hט%� �&x��U�����!~@�g���|�h�A���)4r~��d(t�T��6s�?�JwE�;���՞z�G�#�f�:&��?e�m������5]p�\��T�j�k3b�X%��8 }튢�{u�c��M����5�1�P43��ԣ3�:<�	�.�q��t�i��H#-lI�־y��N�rQ��=��ے�yX�<ح�9mQx�l�S	C�J���˺����r)	�Yp���gY��r1�n�K��N��*K�(�J��$l���C�\!F�6u~�1�'8�J!ƥf�S��{>��L����/����LWh=�}�d���Q��-��T�Gr����7;�_�y_�,܀��z�f)-��9���ǽn�t7�B����ů-�E��K�R�ԣ+8ߘ�Ҙ7�#��x��[D���oT3*�ת6�!�@����VU)���4��nF/|o�dƱ�v3�S���Z�f�T��hv�4L��9��Yw8(:WR�ʓ2���Kᡀ@����=Y�_�7�,l��k���������x삌��Q�K�І��O�B'.��p[<�H�Ҫ4�2�7���'1m�CѝEV�t��Ae@���>)GPU'�0��\p�GO-gi��,���db'Km��;�}���*xpOe�:ɭ�Ew'0����'m�'��^?t�e1���������C���zm�y:$|[���E���Y�v���H�A���Ui��ܻ�ޙ�W];K�,qiR�E�M�������i���&��Z;WA�M��GN�7P}t������+`�T�1v��qR�^�/z��/L��j�k�<l�%~��͏�\���,�}�]�#_Y\(q�a�7J�P�`������,��MA�M��]��u�'�,��"��ٴ)��7�b@���m�Q4�ZS����̉q�T�8ȇ<(�ZN��e�k���5���,�
��2�j��;��
KF�h9�X'�/���;{X6d���c+�TS��yX�s]j�Q�:iU��Z�}' ":� �z��W������)�z����`��|�|�D�t��?��e�� �¥Ȳ�N7�{��fp�O�6���ߍR�{n�m�����,ѫg��n�����+�И��k��iBZ�3��<�qT� ��kDU��	���(�����a@_:j	K�I��0���ŷ 3�"��9їFk_��=MI#K�Oc�t ��Mb�r]�ݼ���T��g�[�6����K)Fy���4���"MF��;����5
�⪘H�Y�������A��[F�� */��Qꎧ�n�5����5$f��\��f�Kж`���^��x���{�t���Y��xH1^8�ԝ8�"R�d��Wx����M��fmL�A�_i�;�A������eM��(Z@������ռ��":XY��j�Ia�t=���!D!=�L�5�/|�l!�<���C��DŶ����HG����[h����k6�����n��Sh�u8����h���{�j��vm���݅���f�v��8��Rsn����o�G����G�TV.�.��!��iK:=��n�AfCd�6�ol� 崋�Q%vxOo��2n�AxBw�EЕY48�k-I���Q>�2�MT���H�Y�=�����*3�T���i=��UȒ����4��\ސb�-��[[��63_���a]\i�S���Q�Ή~�ڏd\	l�f��]�c��[��U�N����Ύ�Ѐ\b�v�_nja�e��[�.}��r��!�t[ю�$�%�����&�2�LCc:r�:���.�=�+��=�����;��|���@H+ө�|�Qɰ�i�#�����@�~턒�dC��yʯן�w�!���6�G+&,�~'<��@���SD�9?ze�t��O #8ܺ� ��Imx#�����G{E�
O�mpCaj�~��[Q��}�{��.�g��I4��{�K6i�Rn0��nXhU��XuV��x<*�*�'����A�zI�V���k�B:,LQTz��S��7��_f2Ҝ����i��UP�?yy��E�2BΘ�"U�a��k]ZЍ��4:&��"!���T�2XOS�%��K���Z����� �9�v�N��D�#�J�g�Tgh_�zz���v��g̼�e��"Q�L�-��\��1b��z�]��V���! �e'l�:H���o�ޓS?�I��0W,�B����hw��d?Ω ��	�~B
i���4|O�7�1d��d�%5������3j��:
��P��E��7����T=��V,���M!�0ʏ�U�fdЯ�?��ڰg��<�h��B�=��3��[�:|�dQ�H5JG��舊��}�|{ȋ?�ks�M?��22{�i� ��K�At���<u9�B=�:�N�����Q�����?�JE�5��y@T� �I�F�r:t���U�������I��[P�9��F��@�+������J�?4�H�]��sK�:����	�E��Ċ
�k[G��?@��aBȵH�Lϸ,� ��\�.@隻HH+�+�������׶ǟ:��Hj��>W�Z�/��Ǭ�����BZ�T��p�Vu�@��U����Y�W�o�~���G.κ��d{�Ŗ)���P$�L������������8?>`篔�ړ�g��]�Zy|���	�0��k�w�r��:�D�4=���

�ӘW��e�1$����k�9�k����ְ�1��Ѿ�]g���f�0�J娉���ރ�?0MW��X[ٮ�a �dm<P]Rv�^�[��D�P�:դ���}�����'��h�H�N�W]��X񵗡���/���<Ϫ�{�'j��eGeAm���#��/��D�|ٯ{��[�M^��v6�/1dh��4�/h-�)H�_�0^цb��25�"t�SX��yX�cT�/\�-���^��o�;C\���slw�1�r	y���L�!�?�	��#8������|�)�c@�}��Q�O�*:�xw��	q�����VM��{��J��Θ�:)��W ��cj��SI��k[�+$&�r ���/,Dj���-=�h��O*��x�t+�7_w?���x�J� ���]s�R�B�@J,1v�T�l�&�cd��H���L"S����{?U�����P[w|Fr,�4ts�M�>]��5����z�ahy)2�*d�ڮ8��4|t�H�hCӃ4����N,�
���VO�bw�{|��Rb�9	|�aJb����zm���p2�o��@�b����j���;ɶ�&(�@����Q��;�� �y?A���f~���������h�Kq��͜��[{���7�o���`��'�WE��Y�ӂ݂i!����������+�2�����R��%��I�%�vA���~1�]���n�m'@A,��Hc���r6E{׋c.R8�X�w���U��'��P�{~�A.{!
�5��6�H@�y>���h��s�@1���T �EQBb�Y�)
�]8G��,sY����0����H�X��j�&��?����հ�4��ڄZ�>��I[w(���(�wZ�^��-�Z�� �p1��_o����	��9C���#y:�9w~�ܦOZpy��������G����;�]��jP{bm�����^G?��elH ����,�Ҭ�#94sq������U�<��԰tQ���#�ɥOSD��ѷ���a}/Z��#���I�g��**aI�>�/�tu�W�`dX�0�D�.=7��sC�6�%���� kv���VsMe�Ɇ�^��}�����{�5'��T8_��4<W)zO�ru6��mK�TO�����&�uj�vX�Cm����h���jyK.晢���]����p�G�̖+O,�DU����w�D�eF�8��C�����m�ݚ�h�0��:�dn�L�m>"�7a��݈Ӛ�t��b߯����d���eO��:9�iM�x�qa|�E��Zl��V�s��<���Ջl���/��,}2)j�>r8Gf��0� a�߿j��Wf@���4i�[+\�/�E�af�>���&5�Pl�y�>����苢~?(ʛ������G��e� 8'���K�x7v��)y*�� ��s���:}���ӗF�<jv[	�A�Rj�ƾ߯�YkԨ�sŠ4k_�9秂�H�ظ^M%���6	R�(a��8Y��/U*�2Ft>�U~��2*�; �y���ܝəN^�����;�v ����Q��B�XSP;}��h}�YQ�� Y
��#Q��W��c]X��T>93�Y�h[�+5lH"��X]���F�F*��r{��<a߼T�jf�����6,�`�U� AI�
�����'�� ���-�|Rb+�U>�����X��6I�9�I"l�������h����Z2�P���9�Y���N���Ҹp�(l�fQM��� �A���\�3$9�M�fQ0J�}�J��ov�X-�Ȇ�743Q�؀V|�xu'E�W����;'�L��)2! kyD�iT���A�l�R�R:~'[:k��=<�o^0��FT2�������mS|}�@9����~�5�qt1f7��kx�:.�݌ޠT�(�Y�S�$�}��W�������d U|�epdn�i3�������,B,��}���˗�i���$�;��r�UZ�y����n��_/�*�mW�v��|8�g��v܈p&(��~���������J�
�"������/b�><e<��ߒ��D�q�V|�Y�ɬ.pz�/�?�?�����Yh�W�d��O�I6݉_;䘒==�05b�u�N�|�:�n���CNy���G�U$��ޮ�9o��|�� !����.��+�vO
[�?j�aA�n�;�9<�y�g�E�z�^����l��C?�K��_r~�Yf��y!�0�H���^�s9,aA̞���C�����b��qW���ǭewq���EمYTg�وO{����~G��6=�]�jn4]`L�=Xn��.o�i�D��~�����[�J�������qV�p
�K����z8ж�����8���^|)��[A�i ��2`���� ����.�9_�C(pཝ9k_���1i�D�K�J�ẗ́��b�/���Ӣ��RR4$���E�F��y�q�5b"���J�r�I���cV!�b}s��D?�ɘl���@e�����rJ��
��ww���v�bE"�8zbF�������.+g\"�R� F�OVZj>��B%}�LG��Ӧ%�
b�T/S���fņ�vA�Ԡ�swV5��{]$���|{�;:�f������ƇI
��!��U�w0�X��R~�!�J���:�`��47f��)�tZ�}N4Q���2�%o����يLO�`���-kf�w:)�M�}���W��Z�j���_�x�լ��k�lu3m%N��e�pi)�W;R�X7
mg�ٕ�b��bHK�Z�?���w�7^��Op�}�n%)�h�M�|�7 8����� ��]{g�)?���,T�"*Z��rы��Jo��>��y�C�7q� (]5�Tc���BI,?��ۿ���e��%�`��}�e��lL]���"��xE<6Q3(A��,�}#Q-����:�P�P��t7��q$j(�����k�0I� p�o�=�_`�J�����z!��2Qܵ~ʡ��4��l�%���� ya��V��b��[`�ڒQg�#|�X�ff��[R��kv���D�p��M��ζ^������I��y
]F�^�]�~<-K LXe
���ƍ{��v��[�,�����(�I?��b�=�<XjU��u/4V�Jc�u0�1�����k �M��Jܯi���m�>N6X�u,x��lg����U����K�g �\���<�E����Kf�����O��G����p�æ�@v�}��"�@�G|����S�+��r�����7�S����[�%2��v�y�*Y���|��>�#�Qg�@`�����^<��v�VV��ީ=�o`�������h;�������S�/���k�9sw��0�]�OrA��VL
�Ȧ▃�bV�wrA��o�~k5Rc�c���=fѰ^�TH	u��U54}0�&;߭o�F�6�a`�K@2?H6 ��}�������pN$�@��8���4������i�}���w N6�I�/���s �!�ݓM��gEΥɇ���:/j��`��p��\w^�MU�L��Ë��܇��a�%L#/�C�W� t7�ث�B�]�{N�&{�l��� 6<��E�z3�N����]Eq<�E���ʓz���
D��k��k��i�^g`�%@�-qͺFp��)Z>�y���؜q�qd�^���7x�p�>����@ғ㷑��6hW?�:��ʅ~��;�_\��yk|ڿ%_���
@��K$;���k�+��"u�JЊO�C��C�j���w@�Bʸb�Cͽ1�Jz�j�ӫ�7g?M螊̏�v��J;ȇ%G��8]�F�T��ƌ�Ќ0�K�����O�����σ�<�@��;=0=���u��6u1s �O�����pA�)��1�?ޛL�Ñ��@��H�i��'9�J��q�a:-6�y0�Lya�X���X��� �Duk�Jho˻>�P����X��ǳv8����-��[dR@@��:�W�΅?��^'���^8����+���Nk�32+�bU��Be4�%k��~�q)��޻���z��p���m����`ю5HS��l��6u�{����=�lG�y��z	�&�k��x	���ӄ�+b�
�޹���"�y��/^�a%@�H:9�&�(�bcS�(%n���ŷ\�.`s����c<F֡�{��^f�犝�|^lk�;�fD����l�N�٦b�*�h��I7��H�m�*��h�sυC�����R����T%���L��)�`j9K`�A�ǩ�=3���oX�R",�U��_�λ��P��ݙpmj����p���o��t �|vq�7Y$6��P�o���t�\t�Ȑ�S�MR����N'O~��\���e�$õ�:��	�&������Y�③jz{��5~,ۮ3l�L��D�Iz�7�O�J���MQ�n�
�+}r��l#�g�o�!��թ-�kh820���l6`��R-�~�n�͞��}�T%�0L+|(% F@���`q��������+k�, ��W$�h��ğ��x�܉����D��6es?��f\Rr�� )����t�F�/�����T)~:1��p����Ҷ��6m� ����J��i�Pf��L���j�5C��_������IP�Tz�^'tI4�f#��>gQBN8�q{�޵�Y��e@���M_�j�CŌY'j�	C�t,����,����Y\ʢX�✹��T�sf�JcŧLXV�p�nr��u�l� �_Rn4�������{�OI��b|��&o-e}��n&����Y�#�r+�ؘ�Ŗ�"��
�19S0�_ .��+��q{p-c�z�>�Զ>Di���%L�n���X7��n�/�Geס���,�F�t�~VA�P{@ ��0a�Ν��ɢ�qjm�����0JafOQ�c�0��u����4DeU,�¹��Μ�*sR�y�w�eo���*[�[���U��h���^:����y�G���rX[�XS^䴲BĂ��Ҝ�����8�%����t�T�Ι�'*e������0-��U�l�ǫpP���:_���^ش�{C����� 8v�)}�x�FHʅ�h�&+�2o�qILO�2G�׌�S]kv����aO|.����J<��%.�	�$O^�r"x�^��`�tk�kmz{������%�o,�ߔ�4�`$��H8�4e�=��D �=)%�=�O���s�-�'U�S�R&���0w���:�U;Xs1KY��U}�3����:_��E1@Sk�՝M���S�%J��i�۸��m���{��� #���O��י���.x��C�P�����7-�vk��ͬ�J��/-	H��-U��l8*ou�\ ZFOb�ժ��)s�mߺ�먗(IVV��#��|�[�r,�	�����i�,StnC��q���&f�����r��qo�-7r�Rq����'���75ڝҀ��]��5X���@&�FXv$��%2��,�n����e$��N�������s}�R��[~~@�~@$���4Pj�_O;]�շH�W}Z��}���B"����@��z;�y�	��P��Ux�@T��n˔#3w�5�S�5kg��^�/QmP�lACO�"�c8p�G�K��"Fc0�����j[����� ��]鵴���q�-���k���̿F�c,�8/�"fQ����QM�Q`��#9sk�2�0���������(����"�C�J/��<����s�T{*��MB�f��&w�r��q0��ӄ�G*N�<L;X��ıF|C8��*���"G#�5��6dS�a�B�$[b�xԚ/s���_+P�/{���ňAT��p$HB��qNa~C nO��K)��d����|~�y��ٸm�r�[$�4,nچ֑�/܍#|��%mN�?Y�G��v��mo;��ehEQrO���:���<CϹC�e�3���XU��i;~�2�I��g����R����,��3�,��H��A���lI���пԕT���J!�H=,u V����hZ����p	�� �v(�m��-o_�,�&E߾�x��Ѱ?9��E��)2Ų���rL+Z��{o�'s�ρRHN,3n���r�/2�%k�w��U[�d�R��$'�Ye<�:d��9Jd��7�ͭHy���۸`n9:����#p��m� �X�@;��8X ��@���5 �)a�OT��A�JS�yZ���r��y\͚�D�I��s=	��w��r�B�H.�`٭[��)��szV�O����w��s�8W���YB^d��
}.�wv'���,;����
�J���Nӈa���5�V�L稡7'�z��Y�F^���u;F���2��ba]�\�^r�Gt>A�i���kM^��(��ba �z��\��'g�pb�6<ʯA8�3%]*��8iA�LIɀZt(.>[�E�ZyG��S��[ھ~��U\̯i��m7��S�$&15�j�˲�8��1��j?���j)6�W	�/��jӑ�r��Mה�dA�`��t^9׀eyuQ�xg��^�|oJ]�n��{���dཊ-�fS1��EA�����鈋�+5�w���Կ�||z�(Ň�H]/���ȓ5j��D�-=��Y��\5:��*�p o��4��G"���v%�l�kt"��r��G�9���n�vΥ�>��5Ƴq�=�njk6b�Pq*g���,[��8@-v:^p<Qf��t���r�	�K�(J"bʲ"�K������~SzV��]��*��/�+W��v��e�rl��3��<�?�t�$Μ� ���y��.��x�<�H�=��ᰦ�|8� �x�S�����X` ��y/�=����Y�P��ʊ���W����l;���f3�"��F��Ƚc�C�| �&���
��v�PR�	���,[;t�)-���!��7��?�v�� ���(	�7Y^��r恡�4�BN$����SKg����)��������#�U�H$+R�����ek�LizN��'�Z���V�k��>���:��*=�^���`�]n�)L�x��8��Zca�Hn6�*�_h�F�/��f�Tf���S�&LB��i��{�Vt۳�+��"1�p�g����c�#��W��~��)��W
�Ū��^L��6%�Z�ֻ��F7���/�v���C����rS�ʰ�p:��e����g�u/�R�6Ԅ@�2Ѥ b�3o������B	��#S���%4��l;J�*N>��F]"%�
�Ȱ�C�����g?�n8BP0AE"9�[�K����&�"  ��_ŀ��/��7� ����4��/�#�y�]�)+9��M3�)���)D�O�\'��`�����;��ɺ++O�{6�[�6�r>2c���E��7揝���������q���_$�Z:��w�!a
�M�-2[T�}���
�9�oڌ�rlA�G�L6i.4�X��%���d'�f�q�fi���.�z�~�}1�t���	�����4�V� -���<fT��a�V�σ���&�"�"E��ߚX�?���:S5N�J�v	7��{��.Z`���S��pg�����bug��E���tE��>Dwf/�y�|EsSp /�-��iD�{�I�M'7�I�K1d�������Kk�CMh勢�����l�>��y����I�d؆۶P�	?k\�>�林�`���IWLsl,�+����67Y�tl4����$�մ>�<"��rr����l�}�0*�tq���O���h#�O�30����r�į�$%�r�
�Π4�����lXt�1k��
�dw�lb-�P�H`Jڒ�;%�L���,�r�Ɵ�1˦ɰ�>�����.�=��(�d�y�-t��ž�q�}N���z$��G�5N��z]Հm�X�?�;̺U�l�r�W�|�[b��y|�;� O��/��<��N��:��Q�*/�z�.'�I�_�2���C�.$~�3����1�����0�QbS����E��߶Ȑ��mr���{�g�/�?���i%����3���v�M|s����&�&G�ݘ������hM�]�|b`�E�;p�3�Q~����Q��V�s�)&�4mV�FB��86.n��1�(6���mQ'(�7Z�=����8ێ�~���U�0��5�J�=�{�:�1AJ�OZ�Qv��x�${9h�M}��"�b�]X���MQ�ǳ~��N1;�4~���Y��b~�S4.o��=jk�A�5���_NY�z@�����m�*��F��	��.�,�<_��o�}h�����5칸�-���e�g?�a�{�8��*U��q�'��c^p�8d7�z��P��"���1S�uoPAa ��"TÈ�0I��#���b�Y}�'0F�~�8Z��ۥ<m?�����>�t��o�*���
	�5�]S��X�fN.�|�Gť%(�V,w�r���'�ۅSfs�v��L�c��㎱���RN��+&ߎ�4�h�����rP� �I]��F"{=���������S���Q��#�@�_9�eo8�Ɏ��sW�<sX�`�fQ�ļ�c:� ^���bp����FG���G�4�����v���.�E�����qRc��-�-��	Y/B�di�vk2�=*C�+R*��S1rr���d>�b�� }���2���'���Q�=���_���'E{�c�1�H��U�ZZ!�4z�d��(��~!�랭(�E�@�:T��qŰ�:��\���F��#Z��7@P���1�Jj�c���X�:�RW*�{�2��U�t����,rh��D��=��x��rp�E�����^5��A�2����~6�St	؄[���_9ɼ�df�����޲��)��2�V���C�[������u��#�������nY(�!K��8#s3��F2��'���(�;J��e����]�~޻:���=���P�4>q���O�2�
8�5��Rp��)���28����	��H��A̆FAKKm���C�׏��W�6l�c�L>�%쭏��!<uT����Y�TN���d�MI�z(�O�9�h�����_N��3�%z�R�c��L�!h���x�S�y=�ӚI�k]ɿ� ����
��  .�f�w[>a��͇!��?	VbO�J����&��\��Qm�4�w��; }ʞ��i�BA�B��4V��Zl�Q9}݁hL�������~�qAm@�k�m+�0�4����3�����$���֠��!�-��J	�Y�N���%eh|�B�`��
v$�����7멹|���B[6
y�')�xA�>�k�s0�c�U���!�ûyH Q�����6z��ٽi)_��FK^%̊:f���f� �S�yLs���7a��7P ��(}��c����7,>�욜V�N���%�6�Ap������g��]L�͎��mp���O��d���W�� ��-ꠕ�����N�-�����`�� b�:�p7��C�M�n=剕��PX�P�w������\J�Nf�^�n��:�5т�	-�%�X�����OY���lE�5�d���F�;L�3GS/��N{v87�N��n���1�����b��մ!���ϸ� �tiS���*|��~����%��ʙ��
y%�;�W�h5�W����K�((��nn���?�Ԣo����"��D���,ޭ���n�M�N1X��g���r�`-[jf�~}��{`qk�Ə�`� l���_����+P�@��g�+xX ��B�&�N �w}������#M��4}ג�O��?��e�b�y}e)z��W�3�Ö[������3C˘�~�R�`��}�3i���wE���v�l��{C��� ������|X),��q=��l0��3m>yP�0�CY2���%7*�2�4^���[j�����9OЪ��zX��MQ����/����!�J�8	�VhUG�y �n�[P=�R���z�@��U��c˗ez�5ϗkT�R`���4 !�'w�Ӥ�M�W��MG.i�� �|gR�	e��s��VvF��q`"�):��٨)i�)��Je���A���/q�09
�� ���;���h��ɤ\�v��'�ު<����;�{�M�TT=[����G��X�axy2c��V+�BWkSf�z���:t�����pH֛ax��2Tw�(?4��x:�3I�i/��߁+b��%'��Z��U���G<˧F;��u�:Q&�Iw@.W�\o�N�i�g��%l�b٘k�� d�����w,�cP��$}�@�rҏ̪ݻ}z֏��Y�5gd ���.�)�����QV
mq�^t"dz���S���L����y
�ji՛���
�Բ�d"
}mV�"���ʊ��i���.�z~����P+-0w�ښmZ��ۭن\��=��M4���h���&G�#mv���@����6�Br��9ꑍpJZw�O���5B��ӱ�P���%c�yK6�`��^6���aQ�J��%�d���V��,��薾�y��4�p����e�ꙡL�aժ����nܻ`=���?P(�7!�sGt:����HNb��j�⦓�C9�E/���w��7 v����A�-nzĳ���my*�O�o,��l9�8|-�c��+A����X����v)��F�kˆ��ӗ�6F6��?�n瘦1pE�+��-���czyd�KH�d����{&+�m�EK- �#R���1�B(��|^,���K �����*��X����x��faQ��`A��-F�6�]�[�G_\����0����sR⪥�Pn���3��d��]w#�p����w��i{#.9�M1��5؀ޜ��o]e���K��^��U�eJ%��V��Z<k{���e�����f+��v]O{/�@��}��Z �M#NC&尖�Έ$��}Ia�q��q��e����v؟La��B�8�5��U�Kkjd�XZ�����f}-i��i�gmj�{�,��R�a���	W��O��W�Vah+ݶ�/$F�Sp�9�
�� d�ndhֈ|�g-٢����첯�X�8��Q#�<������.
R��=���c�9����[��7E*E	�ɚ����1�G�f�:ܤ6�9�(*�~�H a��n1�)�0")����2
0���p�:�+���j��0�c�s�h��B���h�֩K�����_xp/��La�t�� ��6a����/.��C׍QW�8]6z�,�����+�ߏ��@!�D�`5��may(�\]�B`]�xm�-���Ljq�S�a���o��
s/l;4�J"�B���xe��B��s�Н!�q1M'�`���f�u��8�%�_t�i��mE��}ͩ��[A���[����˸,?C��㔗(��XB7���N?��xǠuL��z$���{K�Qҋ���ρp�f��~_�]p�ݏ�m��8�	O�w��3���B������� �E2m�j��^(j�>��l�W�d�L��h����G��lb,*�tiTe���Pk��\N���u{������`����۝l̞�eRo����r]�Y#���q����L�r7Z8��מ�'	�����Z?��B#3�P�]	}�Q�xm�6�w	].����{��v���y�@�9�Z��|�g��m�I7�vU��Z��W$��l��,C���a&b,�E}%�I_�
�[%n�r/�%U���F� �x�W���M.��ͳk�N��4i�A�yXR�R/t?��~	�����������Wf���֪�_Сw�����S�ʋ�gI6E�w����I���˩�<RK7�zp�ʂm@'�㏬�|ǳ�>�<?�uF��l�z�πU�1�@(�&��s(�kw�s\uUڅ	�[�<]����Z�T)���!��nUILa��6��[Be���������]�����h]Μ�ȃ�2��l-șn�~��WK����+���z{�}�#\U=��r������&�5IS��0�l�h�R&�D�k���8%�`|�Bha�٥���_����?�T<�3��"�B�6
ȯŒ����Z-�-3:�w�(��G��e*�mH[?U`���Yo��i�|��K��ް� ��b����f�ڛt�
\Ԫg�
J��z��?��L@����Z����k�\z�,�s؝[�c$ =5�^ �4`��i 8vz�rP�ȃ9�,�upT�|$
ϥ�_��J�X<�?B�GK�kyޚ���!�if�����Vԭ�8�g�l��"���6^6#}v��f�����6�������WNva@�նU�V�[�I�1�M�0R�I�W�V���hߴQ�|��tdyN���+Yz������i\����U�D��Is�qX]Ȩ�]�Ф��b��!��G��`�i�	�w�a�E�v����+?%���#y�] �!L���M�u%�+ �t�~��8�n�u��X�'z��rG���g��.t�~���*�	�'P��b	��{��<��o����Y�XBM�â�?�p�	�a,��ٱ�֝���OF.�4~(I�)8M�COtd�Y҅��a��x%�S. T�$f ٛ�?�U6���A�A��ε#�j���g���")`@�j%lR�N�cZ�1�Lt��?)4�)ٍA�Mz��)G1���i����)	�u��1WT'����K���u���3�aCN�DG�-�3`�i'���K1�r���J��rU�಄^���m�j���(HD�A����������0�����ʉ��9|p�!e����E���Á�6����1�EU!v���!��̱:��U�eѝg<&w��m����c�
��c�+$�2�j�T��sڌ�ɠ䮊[5h&���wc��H�/rȄ�gX�sqf�&��ed<J�޸@"9���*���s�����J�{�.��ÞW�̻PE��9��:��ڙ��!�}u�y8�uy�V �q�@aq �J�O�{��&o<�@CART^�b�K�yE�.��L�㽱���yNL5|T��Xňg�;E��ao��d`(������[���
%�9����L������s *�I[X�����72�M8��̰{�����e��r���y�-���O\mL���Ip�:�%Y�x�Nzե�����'��H}���� O�D�XMqL-;�ⴿ]
�-2�u���7l69C4(9/���\���)�j�1�Wt�B���Չ��$���YV��D	�" ��M��^�Z7��Ԑ��!,�t���:���n�����V�X��������0�$f�:�e]D�.o#����U�����r�cN���)�`����/cdq�d��N:�!��^���D��3y���B��q�q~����~�Y�o����6W���~�sm����+��p�0Z��cxo��PT8�c(R���������Xfn��
OPPj\c�wU���3�t�5����ьm�٠���j2��zz�\n�?���,��HN��6|z�^⟫�gV��9\����[����k����z��o���Ǹ�%��dS%����s��Z�$�u�X�X�̢7�l�X��HC���
� EM՗��ߋ8ϊ�~'?b{�@?�ދ!Z�ݯ���C��"u��Ϛ�b�p]�I�-��mc+tZ�u=h:v5���ѓ��g�;`�����6��
1S1������)�;-X���lu� �i�T���[m���PR
���1��:�Ȩ��@�X�0�'��t�O�d��q�E���/���5��/ǆ� �8��	$�u�virD�`��<�ֆ�[z����lN wD��%�Q1g�'�&��4�b�X:uBF	ù��S�X�ǆ�;;3v�����OO0�+Hֹ��]i��?S[El_i��P��T�1��">O���^ o�ǈ�����ggq.a������H��K[)���?�)�?����(�OdNJs���ca��^�ܹ�7$fh.Y'􈓄1�5H�č�l�9����:q�Nn�v�Q��_{�%����(�w ��6��"LE)�+��e��k!KJ(�N�J!�*hL�a��C�0�Y�o��_���_���C=������'�{:L� ~��.,�&n� 4����ڽ�m�۳����)PJƢqW�#�̥����뽀P�|[ڗ(FFD�|�6�䖓;�+�E�ݛd;qz�T��K�����]�*_�_��(u�3I*K�����H�`����ĺJ�AjX���Qg��.]Y/�㽞��� <!��ԕ����׿\@��o��%�tL�y�㕴B#�j%F@>��wį�IE��<l���\I�T�V��:��RHV�d�4Á`3��,�^�/�xv��*�"�P��e�c*�%�me�Q�Δ����]��=l'�FM)��J������zk%�yp<Áp�ʷW�$�cH������ʉ#j��XUp�n%�]ǡӳ��jK�\|fl�RAs|%;$iY�&�*ۜޕ�S-����s�L3��g.��4 ����F�;�G�11�֦N�LH��t|Ʀ��[߭:s�������Q���%DR��~Ʉ�Ɠ�Ӎ�K9sw���o6�Ӹ=�FV74p�Ԭ����$�1�EaM���zt�ꇡt�$��&��L��ஷ�w�rcK528��%�ڊ<֒AW����eC�I{���.�֙���'��n��7Ԯ'���¸�Dr��RH��K�N�R\���v0&5lد�\ҹj`Jrgxuc�= ߚ���Z4�OUHFy�|�~�e%�;����{"��ϲ8r�4עk�tO\��vm��^��p*1��)��s���o�x����~YyA�qc�X���<��v33tEu_�}�Pï�9�$���r�����+�H[�H�ᓗWr�)��P�	�o��(3zX�Y���tY�$����9� ��k[��x<cgn	}T}��đ/!1P�u��L�4�0���ZL ְ����E�!��9Lg+}`�2�����`��i��Z�Tt4GW�⍳oM������t�ۻ���%+�v�#�:H$��\���i|86F>��������x ��Y�$��E7h4�'xaY@��2o�b���>��t�zdy�q��.�z�3���Gﶷ�3�mu��+��"o\� &���=���F�2���8�Q��P($�a��/v����h-f	.D�5�=%�da�d}����G���7�z��.�c9������N��3�9��y5�����[�F�"F��t[o����$a���S���������X!��L@�A�ؠ�Q�W� ���K���a?���x_UZEY_� �J�a��8�cQH��,)����6���	��ys�Uoؑ ��#�\x�y@�њ��*	���x���F�VM��.�7��P�,�5Ƕ�Z(>��D~��.~�tz_�%�Y�l��&��cJ�ΰ��Z	�1C@����J6.���h��զ \C���P��8*�����1���1�S�B��0
�$?<Htb�H��(3�]:F��c���_��2oY�����b[ǂTpN4�;$�:��'�}������/M� -"h[V����R��M�\�	��:I5?HL�&&N�� $�_.�����Tdٍ��FP2��4]���3��1*��H"��^�sI��,�-0JM�	�.�J��%��4D-�G\l1A0i�i$�>��+X�ͽU��2=ܖ���C���7�,��7�C�^�s�����}�e�D�WQ�K�C�ځ��(�餱��@�C�q��7�k{,�3ArI�<���f?�s��Qf��.����]��om��p}��E}�ZuPB1�U"o���a{y�^���9~j{f�?��a��61Z-(-�!��ڡ���H�r���Th�R�����>[cf��d��
��wv�_�?������:��g���%4C�p>��G��v!���b{â��@4
��]��ڍ�#�W!qb�颞0P�e�X�D^H����mϟ"�������M�&�z��O�4��W$8g��K�?#BK;\�d�����74�v7_�U����f�#�1v�i��\��e_���:R����n��b���X���ly��p�?s/���<V��8�ִU�C�O�	 C���q���ߏBE�u��n��O��`['���d­�D^�v�Ůw�vt�rA?80�U	>g�3]�҄h�j��;��D4�M�O$7"�<�c�B�"��
4]YIZ���a&��v2��<ӌ����X0��M���ﾐcI/�����M�����R=OZ��K��vq��b��*��r݉�^��&��	,.��
���W�R�$�<y�L���O�?#�q`M�a�ަ3��}2�p1�\W�XG� ��Ld��0t�w�g�F����e�u������/� ���8�qJI�U�J3��j�&��������XIOUA���e��$a@���O|a��F�6kx0dY��/	'��%&)�󿰮���������QJK����6=��A
��F���u����k%�6f��[�	��>�@J��z>8d�6>�5�-v�X=/��Α6:�v�������s��4���ʘ�
�vl,���:��My�O�I�='�ɬ���ԁb��d���H��r��P/+ѓkaEh�?��Á��h�Ħf��,$T��&�>I�g���G�3.�y/���K<���K�zm��b(�ӣ���0/�� ��<,��T2�P.|yq�G�c���#gV�-��U�,��%׏�0��G������_�(��6Eӗ�-�tȏ)^�v�A��x���)�͌�`
���l!z=B���]x�����(073)s}��
nB����8�q��-X��Pի0����܈&���:���/B� ,��������Ar�b_��*Z�7�?�WК��-Z?���Y��Ey�p��ۈ�7�ڃ����@�hj��XDE(&���G�Q�b2�q�������ʋ2����`+��	�}��N>5��oP2q��'R@�|�AT��au��GBs���:��R,Q�*�N2�o#j���03�g������Y|�b����Ov���ְń �2�}�%�����5H�DW��0�O�}�{�f��m�a�f���<��Yj��J�j��Pw���_]�X�NP���i�,q�|(Rp��$0=�[)�3/�I'��u�Q�����S�5�h�2�z���Oˊ(����g.c����k�^�ِ�:ϒ�� ���]�?<|��5� p�xX�p���HTׅR`��ԁ[ sg��4�5�aj~�U�hbo}Z�������e��L�l�8��M
�f������ʄV�F�j�\��aĖ�=���n䙋;�c�_j��m�N��_#x0yK;���f�RG3��{��q�ڶ��>�p�"�'B�Lį��'��������N�cSޕnD~5�-g��.�N�!�u�_��FÅa(�)�'�5���*ܩ'M8�YY��i�O�
��4��׋�D�a����N?���P3y��7�_�1k�yk9[s@�켖]��>��1HN4�m(�0����F��E������O�ۆ�z#���rVNW���H��P���b±䙔�(�Bx�l~g� ��r��]��3mq~��.!���-E-1��d��9~q��|��*��{�A(��ZUٰnwФ����4��ɫ��k��LX�.��
�cZ�.��c&�&����0�T4�J�٫׼���)��н.�hg/4���#�g�0;�A:�H�ߖ{Je��L����ۃW<�'��e}_����G�����ړo^^���\��$n����<�R"eM
��WxS��{0zl�,��D�i��%ŕ��y(Ҍ3���^�`������-�I֪K����� ����V~YI�Z8�L������o����j�9sk"��^��7��)Ѯ>3�����w3�D>0`�� �K�5�g�V�"�F�R\ڄ����Ӯj%��Yo�Z��'[�Y����Cs�3j�&�"^\O��Osދ�=0_�9�O��+(��k����L|%�z�}C=�ɘR*|R��.x�W�����vq������⤠�Y۠���k�a,?0=Ųf>�GP���/Ѐl��u����X��l�7�ם���Эm�����ʨS�&���dmN�>f��RLK��u�gb8Z�(й_�7��Z=�!�Aw��:�&7���>R���I��B�3���:�tKz���}OW��'�m�0��ˎ���yK��-R_��ܗI�p4]-+�=��,����c���\���w�t�S'��72S��b�]�"���N����9���u֯fp�k���#P��ep��0V��IK]�g�* ��`"���ӕ-�ǟ�K���#ۥ�Ke�fqk
��ze`5U#��0uZLa��J��������RձP��ܯ���j�<����R�!�%ql�X돞qvDJjwI�r�t��~ ��p?8��'+�])������@'1�")=����KH�j�ߍ��t֤����&��d��~�j�*Vb/�����/�3SY�S>�fp��3���~:��c����R*�*8�Z�.�h�&�b��:�
�_I�}b��>�A�_
�F]K�$��le_�S_�@��:k�`�+��̬T��+��߆pJC���jv�7v����"�^{F��y�Va̝;1+�a���?cv4�K�,�J&<�[+�J(.�� K�T/�����K
^�"Z1w���wɪda��G5�iT����fՉǠ�O�CCYB\�]�t��j[ ����u4w���>~KZtv��A��V٥X��u����nah�����a�Xs��ڽ՜C1?J�O[��u|�YY'o�(4�3�.~�(% k��Dn6��m��"`�<�
)�*���~�B��=$��X'����Apb�x:�J�;x�5{�O�p8�VE����IaD&��Z��'���V�\���?���c���Q��l��ҝ��+kwXfי��c_��]cw��8�ӾA�؊��ֶ�`^Ƅ�VEy�qn�f)��;o��]N l?_|�Yx��-(O��Kן��y��5�N��*GL�ޏ�Y�Ig����W��-���Ӕ��_�[�U�2�"%�7	6�/?jD� y��m�7DO͵���"2'z����.��4�س��D�u�&���/y�����H�OI[Q-oV�u�:R]�k�>�{*����8�%�=�;)�ƹ����2*�U�!���e��]��J�;Bʌ��o윆��m�D�H���m�x���Es���B�8��A4��A��&���A$��H� vG�̂���tA�e=������]��̹P�����M�`��6�C�
�{�h݌,����oG�2Cv�a�B���$���+#Z)���B�ÎYז?qE��p�B�Z�4х��8S�y^�(Jk�ת^X�l�g��}c�����؍��2�I�{��'�i~k���$+^��
�!��{J��jZ_`���a���vr�N�^m�r)��3/z\�E�b�Sh2%͆*�PA�T���r�Z��$f���am#ঽ��'��3>�H��'�f�����]�����ra��#��]kV��԰.����j���L�-xj$)s�U�}�0Gǝ��K��Y�\�o��{���+U�բ��C;Ǐ��H ����0�PСu6�����J�f�>�������q���`7	�rJ����R}_�W{G�&�'�\�w�q�����m	I���-��/����Gm >0�s<����݇��;H�싢�J 7�cc���xl)�1l�Cb�P�]W��4 kw(��<5u�xsN|m����Z�b��9ե�;*���&}�H�z�ߨh5�;����Q6;a=�c��f�n�����@|�c
�O�G"��.��d:aDQݨ�O֣���B��pu�@/\�,dY�Qꬪ�3� ⳯j0��p�-������4���T��A��éjw�-\d&A���vW�y��G37�8��8ZdR�n���D���f��Nx�N�;'����!ZbUr"��C������WB�o��+Y�C�ؙ�]����#���:��[��mk���ަ�\]:��K����~�����ēB�N\�F?V��&p����tX`�'c;��Z@n���"��E�!2����&��q�(��d��[ �&�&.�͒����=��x��n��c-3`	�C�"O���$�"꛸�5a��j�?�BqR��_���%��5��j&�c�(\P0��C���%�B^�<o;OlS�,�g�0#����ǳ��Ø����!$��߶�b5�g�֊���Ҟ�>`��A)gb�S��/��?�_I���^R�h7��:�m�j׸A4s�rXש+�eJ����ʲ2&E)ٔ�퍝�ߌ�	���S~�� �.kU����бB�c��n��,�\	Ju0�Tm��2�&�-a�9Nc�u:�]���W�[�h'@Fh�}z`Dr�r��v��n@���Eq�sP�Q?��[�������%컌���yh�PD��������ND�{���57�D�ik#�X� ѓ`��S=}p��j��W��A������OX��;�MWJ\h
�U����UE�E�Ң�ت^��~�#�p!�q�p�iWK�{"�
 �j�0 ���D>�Ґ����K�e����Ѐ�EӐw|s�?a� P�]�p1��x��,��Vc�u=�E:D�)�4Ї?OH7��E����8Z�����`�����ޒ�QZǭ��ÜQ">��H!a ;���/57�๬�l��ޕ�f��)�9t��,EL���U{�����K|���e.�3���S!:�nb�tqa�M�M|��;Sw��&[Q�R9]���a���%n]!\�r
1$�|ߒ��s�]a������9Xy��ͳ��ظnT}��J����R'�<+	Z�
��v�ꘗ�������+��/DxE<��tp�`�k�㻦���v�SAe��'F"1j���`�����>8f~�痄ݛ���l�Zra�������d�(y~5jR��;3Gg�,�
Ji�Ѐ	��uo\��ep��ξ�,�f�T����ɰƊ��[���^�ڙ81�@���6�K�}�l�����YP�%2�#�h����O��<t����,i �o����F���k����).*�����3F�u��lx�<B5J<�7*M��Mn/�$oEP�Z]�v����G�	2�e�3H7Z0�Z^�"��YK�������k�Pom+�����
��ԅ���ү�`]p�����\�6O,��:HT�����G^����$��/�H�Kbn��`j��67��ëKZNeQ
Rt[;k䐿]뛫yu���[� !��Q���#��(#xX�pe5��b4nS��9B��J�?�җ�E�F\��]����ʺ��/7��Y\��a9�6��iQ��d�Q��.d�����,�4�\�+,���Mٰ�6p�WU�7�yk;]r^:zf~g/ E�	v��I�Ge*Â�:ސ���u��f�Y
\'�ީ1u��W�s]@�Z��e:z��J�>s\����%�@��1�B��-�s�(m�IE`����ܮ=��?t>SڊM�*�eSԕ��s�"ηYvI��Ht�\��8�ˢ3~+�Gm(1�u�'^�g��]��B��p�w����N)�A�2-o6K*�cɺ����v�>x`�c���RE�<���$�4�X��{	_e����kf0��6fBC4L���l{e�v77h# �F����y̔<����Kaڭ��B0�t7n/�k�Kyn�U�7�Ʊ�����b����ߡ�~:g���8���ʅ[�{���P��0rlu�����G`U�iYs�SCɆ�O@�s?͒�=F.���%ocZ��n�풒��,�x�����u5_ѕ���K��v]�/�| }%|=�Y��0�����8��+-8Nƍ"�ʀ�T��U3��v�\��?Uik(n%�\3Ce�aNFle��׀�(�{�L��fw�0w�Vq��{�8�L{δ��xh�e\3�lv�w�O���a�PsBx�	��װE�|�7$>�k�1�|w~N'��a�t�����.de[**��C��t*��u�#��B/�s�	[O�-�e����Q��[�
(�����9����+�b[t�٩;B�+�ُgR����a��d��dCi�].�/-6.�C�3n�]�N4'�	+_h�>�����a��.���(�@.�-�yO�f�&���Wj��J�l�Ce=�\ ב�F�r�-�uK�-0M��g��8[4b���im9�@�[Ȕ#���N�`Nf�S+����^]�?4*+�7s��[���h~�+S����Hd�i�$�.*���C�,�xd�`_? �6E�L�h�nyQ�6y��81� �߹D�
���L�K���'�7
Ն;y(y��?�r�~x�2	�ap�
�l�����p7%u��T@�l)�Rl��t�(
���7I!H��U�
c�xPs��p�i����Z�{^`Q��#��:�#���kNZ*��-h`��G��<]���䡅�4˖�~w�V��VƐd�����ɷ�]r,\
�]� ��A��kf�c'����=n1=4b��۵���|�M�� �v�hb�H,���
�5��mg�1�l���Bf�\|ϰ��sԭ���*��[�8�J@:B���#�Mɋ����'��0p>r?�e.x2��3�3>�~�Me�ě8��\T�����M���ؽN�x���c����.�K��r܈��+������Sè��g=Vm�+�+qyɸ��G�}�OT/�qhEz��tZ23�Ά�Ձ_�A.銋F4��6 m!&N����e��69b+�s|��Sܲ����Ɗ·����1��M]��Y҄��+�7��o��edRE}?sh|G�xpk� p{4L��cf�^�D�7h�"ÏO��X�%�	�a�O��no����1ǆĎ�8�MF�-/�;�ss}�����ٓ�����&4�'cT!�l^&�4ʉ�6���l�A�H��P����K"��B�q
�逳,�^D8Q���t�ֶ��n�	�z�4��ꕟZ3�n ��ӄ��bS�<��8T<����k9�f����U�u�91��[�Ǡ�� R�$���a�2����
t��O�������d�1)�0���5Ej��-1UF�H�28,a$fM�����:�	VZJwW�t>���~x�E���׍��&r{��$�ݒ8ʏ(O9� ��l���G���;E�#��%��Z���Zi(��_:f�7���h�Ĩ�ELh�JG��Q9l�_:�vT��/��y�aCȋ�3	�N�t�?_я\*��@�1�jM�0��е�_^���H�!���4�.���P�q��$�XTBL��XzdP�ϕk�K^3.*Ke�P6UÿG��7�ԇ1��Cd�?�?YX ?͑D�c�U´��H]� �F�6�뵋䝩S��'%��D-'��8�(���YJW�Z�umB��!�����(����#��%_�j�˚y�M<6R�G�|�ȓ^v�`�q.
�ˆ��v��_&�Q���m��:k����?�P�Gm�؛�iؿ��fP}K/��H�Yn��vel�Cj;m�2F��6�)�v,4*	���-��l�e���c��1Z/��� j�Tn�6���(|G�q/^M��oz�5�����g�0��t��h����K�i�R�(9MZ���k7�=z�my�h�b�{��yl�+<1mN$��u���!==����>
��(�1_�IY�<�&t䙒��Kd��@о��o`Zr:�#?2�):�d��QvW�@���^�m󩽚�a%sNw�2�珺ְ�(�*�B�ft (r��c<g�2���U�|��q���aU+mX��h��l1$�](*Y<M��^dF�r�J��N��xO}��/�^ݮ�"��	�a��OjR7B0z�v�A�0a�e$��7iؚO�p�j����.8'v@0{�����%7k.�fl�����x�X�fb���t�f8xj�5�(�W��������2KŠ*�|���.�qG�n�.���o�T��r�Lt�=��\J��/�:dsΤ�v�����p�1W�	|�Μ�s�H~��K��ف��]�t�4���� �:�Ѓu����6�]�;b��������P�W�ʿď�ƬI�33�8���a��}�J|��x�� ���xpۣ����&��	�s��5[�:����u^�K(���`�@�F��?VyW�����͓|#o7�p�q��*�7Nn�?�
��o�{��� C�oN�@��Sl��,�i�7Ǐ=�5?	��9�͈7M�B(��,WN�T��{�[�k����Cc�-�jI���҄��u��
�9R� �~i��%��cv�k�:�P -�`�I*�����y�H����WFvV<1s{K��uAC�ShF�y���<�!aC����rK7���W�X���x��n��4I�C�K�x�=� ���	����3�=���ώ�����ü��G����,�����o��'�X�8���>�S�+n���b�� ���%�HYj,89�1ک4��;e��Cv��lZ��#��K 9vW�9���bm0�,�!z��^�R����bZ��$]0$<ͦД!+��L'+�-�жT<!��Vg��U��`�M����6�����d�-��7	��6ݦ��443�;r3I��M������ꛑ�E�	ܔ��{Ó��u���b�*����.�$h��~
$����;?\�'�")���Bە��py͉iz�rr��g?��cK*'���b��;Y`��.#,C���3[������(�Š�;��q�܍mw�y};�D�Ng�b9�^V�7,�MW0��N:b�����y��� �����U:�i���\��uZ	lE��j7"	e�»��h1|dv�m���Q��L����*xc,�|�"��|��:�l�,X�����4�OC֫8Y�����d&lX��pHٱ�}Q/O�H�㷴��C���� ێ&��J�}�5�k�J�T��K~��FF�5X�=K����\FM�<�'�+����ڷ�=z���io��Uqi����_i��}���p��s��	О�K��t�ţ��P�J���
�r3J�Eߑ�p���3�.��(��GE%�r}󏐠?��-4ú!4�Ե7:��4a��Q�F���R.�ir�����@`������.vL%].���<��9����6nެ�u qDl�����m��l�P���|.���4�ՏYeHh����n����OX~,���l��J����5�f]Q��F��[<�W��H�nU{����b�⺮�0@����o�'V Z8�т��;ж��c&T��I�f�K�	LK��:�x&��ɬ����P����Q�V�Ͱ��ʍZ�QEsVš0f��T���}U�� �eP�񦂺L��6"� ��I�>ǫ��|�BY,�ONߥ�69ݒ����	���%*aǋ��ȍ�_u{MK��ؿ������!��	M4,�����b#�\�f��;�b̳K#Q�1-&鰞 a]��ð4�7�_��s�kp�k5�c��N��x�㝮����T8�z�fuR�y�s4p	���JN��m)ǥ�N*�!�� ���t�	��n8 ˲Ɂ����	(|������3_K|�՝*�� ��Y:q�ca��鵆7��}˳{�^��]0�`g'u��A&�\&�cʋ��W�R�ri;�k9۫~H���DG�<��8-�(]I՗/>��P����W��{� �{p���l2S��M^�zLK&>�1�D!�~�֑&���.�6�����ኔ���w�N��� �r���HE�M���:��90e�߃��p��������k��o3J�e��P�2Qܳ)x:��[EWA�r$�/���W+{�ktp�1}���w�6O5�"����4=ΈD�1��Ѫ�Z�5�V�IZN���`���GHR��	�VJ�� 13#/H�2M�H�74����i�	T�Ł���F�gl�=��;��Q�y8.�z��>�W���^�����7^�I��e�mqL.|�+RǨ�k��,a�w�J:�.��*
��	�R�\�iV�-�4x�8g<���)�!7���-AU�!��R��m������֐4�r�;b���m���"̻��x�)|�n���ʭO�El��HV(���%�V���q�h(8˽-������Qk!��������I3w�MO���4�!
5I�4��Pc�t��"�5�<��S&����K���r�W��SK�����10�8��pڄg�R��������`@�T������P�}RZ!c�US�?p�{�KVM����8�)__t��4�fn#���Sq�-�{�2�o�?#�� SM6�f#��{!j���G�;�Ң��F�
��|���o�>�!Po�ɗ�Hu|_�����\8;d�]j���)b������x�o���=[̪�,[i���#�2ܢ ��d��N"�C�|����1'H�P�s_`n���(D�U�RVw������Bg��鑙ԝy��Q�1~'j�{z��A�J�uå�9_��6�����a�3�QǥA���x^�(��˭���T�]Ö�P�Ѹ�����jF�Pؙ#��.}�_LX8_|D��ӹ<
C�1�i�W
��.����D|�b������QQ�ݸ�*k�ҫ �`d}�~�4�X��셜���G����W��r�K��9���܋�o qOt����$0�������8"�D���"LtH⢡�O�f?�dV�G`�O�� ��TNuoR�%�*��r��(D�{�	I@��]LX��ΏT��A�aݐ���W��Xa�g����Pz=}��ۖ�]j���G16��BW<�mUQt�K�ӓF���~��_P�2?�_�K������󡗲�Z_±���A[$�~`&�N�v��G�X��j(������G�U�]�h�y2E�M�PA���L�L_��6s�@ LS2&t�z�k���ק\D�kue�.��y��Że�kv�ށo=��Ej� �cC\}K"{�(��	��U������`�F�-�2��ح՞�÷�;�jC����0�Q9�k(�&,�@h�������=V��������,,'�$5�W��+j����&��a�M�a�<��F����V%�#1AHX~Sz@���_������iZ�������'��=D�&gb�u	9&��<p�[Tb�&^�.��D
|�3�Ϭ��cҠi�@�꿍�vVY��bD������|���CΫy`��n�[��9oI����(���9�f��5ʚ"�IY�}�"p�j09��,�+��i������ȗ���H?^K ��gg�3��H8�����S�M��R�'�%�"��������ׂ�����o�d�_R��'0>E�_�T�0���C�D�!�i<&���Y���=��~�ŕ ��ґ���'r5�a�G � �QS�#+A5閔a�Y��*�q�Dq�0���N�P%�c\�1t�R;XJ8�m�S���T�}h\����٠�C6\v��53W*���îuΟ�~��}�/�:'Q ;z��e`f�s���g���� (\�Țg"�)�x͕�B$��5��,��F`h��4�g�G$�1]��~��
�W�_9�ƴe�"4��[E_�{���b=z�Ԓ1"[���s����
P7�h��WӘg���7p������y-�8�3��wvq�KDM�R<S����]nv�w9#��C@�E�����f�2��>c_+f4�lK�~���(���FG���7YJ��V�a���^�-����1�%�$�ɣ�s�Ї�JӇīwB|���(�_M�\\U'[a&ߠ�x:�4w��"���lG^�[z˓�<B�d!���x�L�˸!���|Ah&�)�6�򋧄M��:�H:˜���*���`L�-�5$�gd���U���q�tiTNe�Sa|]�pI��[W�|��`�����-�*��_w,�5��`���XV/�D4�x��B�&�w���}� �5�����ͣ�Z_�I������<�b�BR���}�z4���­��[P=�P����k���Q ̀V,��#Dh���w�~$��D�?+kJ�&��k��M^�
v���v{&9�9���/�D|Q=�����;ҧ ��w��e7qo���L[�3	}�4�*g�rcR+�t�2����R'��|���` {�aXi�G�Ǝ�"؊jH�mTѱ���&F��B���� �p�=���H��������!>ƋjvS*=*������bQ�v��m!���^�~܏��w�����t/�����)�8ԳXѰ�'ys�}��1MG�;�����p6�2���r^G�A���[�tz/�k���U�U���Dt��	=ӿ.�;d��3��I`�㴥M+��.,"���Xΰ{�����n�ޞ�υ�p����P[� =��B��j�;ְ��������gdqJ�1;gс"�O����f��I�'E�
�\�iջ�=N��橳����a,ax!~l��ma4���"�����6���
�G/�D$��eE{��ڟ<��t���Nlb�Q�� ���D�E<��d>/6n���d�VL|�ID�(VI�$�n󭈐���%�q�Z��jR�0���@T8��^���=Y�!,iʥ�?b��U� �1m���ϼ�I�E��W��@�tS���"��]W�&���>���꨼ C�hub�9H|P�����=5��-�t�գ>����B_ @�,E8X���
菉�Z��	Q�ϡ�g�$X5?��%���k^��Q�᱔�OB�G�zN�R�Lw��*�c.�`����ykYd����S�����m��\9�q`1���|S������c/�έ�KR�W�ԏ��LW��.r#��ޣ��8�b-�:������c�1؀iµsL�������-$�]��h��R���ɉb�t> ΂������m��Uڣ ���M0�RMc�|�2����5`�d[�N2рB��*���n3�P��y���m,9����^����s��M�@�(�CԥQ�f�6F��H9e��3R���޷����k!�%�.)�߻X�"J�P������y;j�B��h����hOjf!��@��͠{�tٶy� c�R�Ӑ[������.�6�cY������l	&��u��l�Tْ��ނ��U�q'b�>��t�Ђu�x<R�,%���lT����SH� �!���#�E�ez��\��d�x7u 7S\���ZC��e�⾌ѰS��F~���y� ��\���X@���b��U�����a���I�m��\�5
�I1�(���/Ə^��y�;�� ^�ow]����Q?��	^_>���$u���u�4�ZO3y�Q����=q�B��x�sdF��:�~��[�2��>��`��@��{lLe7����2_g&5k��d�c��c�`L�1��E�&��r�5�Du`���S��c��E�/��⯋��`>�1��� �n�,��5r{�.7yÿZ�܉<ή엄�܈]B1�a�Y]#(��	
Z}^z�G�8f�e�_�� ?g�XI���Ё�^�q ����k��-��;>e��\�1���T
b��y⫲lQv�s�G0s#�-�9VH���q���I��I{�'T�\T6����.q��V8(=��������bQ}k�cX��(Q�d��������E�
g��21��J�V
I�j�M!P�U������\��ʜ9#0���l��s�ܴ���Y�!c\�p_�@I�Ђ@q@���n��t#-�#쀒�[��ߺy�F�~�A"�V4�� ��"��m��W��A��ȋ���x�Dz�wG�F��-9���*�
sD����R����y��(�Q�l�
}U�ʏ.g�1@yQLs7$��:��R���h?�)0GB�h}c<r�Q`k,D=�Q��1)����mDb��HO���L��N$~_��&�O%ѱ�s�����N`�mSeXX~Z#���'�F�F�ҩt�-����"C�X;2u�T���ߧ��eI��υ��渷Ӗ�(�,�s?�_�ܾ�Jba���ţ'*:L��v��H�W�V1��Z0F;k��� tW�m[�交��so�)�JP<-!=U,.�ygKM�N;�wa~�\��Dmﭫ�*��`��K�Ҥ��F�%4���C.�����o�{5��}��#���x���cQe��l�l�L4p�t�d~�=5n��SS�4���p3��c0P 慄1vh��q	Y������=h���/�|�'Q���-N6�\��=3vk�]_*~
�c�3"ek�~�K���s���n�x����W9��@�w�8(�Z-��W� 5�)H�j��0����!�JE�����,k��k����.�� ���9�r�0UKrw�bʫU��]ݻp̵�KxH�Aڎhx�f3ۄd<���/Ȧ�0�����~]��(���jz�����\ː�Ȓ��.�t��?Ć�ޗ2��v_��ƮOt����
UwR����%�$ʿ�߰ �h�Z�:W*��X�P�Ɔ[�%��Ǝ��'u�P��,�a{o�m7E6ś�^�QNfe}|�m��<��`Ⱦ�k엛�!\r�}U2�?�S����_�W�A��ud\�{�F��.J�9�!�?�ǉ�^�rss<iyN���&>%q?��嶀�u����Ґ��_B��]Dʑ�R��38^T)2�e[����%���Kݭ�"��S4���Kg3L5��3�`���0��t5��s��#��y6B�z�g���Bo��u��$o�ʜ���2�1L{�|���A��Sj���=t��?�^&�е4��/f;��n��u�j>(U�{�����dČ�Xx�������p|�60�Y��R��'%�{~e��\iT�j���LՙX�n�Z�w$<��D�����_���ެe"i�2YS �S����m7|��2�閫�7��ꢜ��ɻ���2#�t�:�3'�ꉟ~
��7�7k�� �ƶXWSj�����H��Ѕ����˝Y7����cl^w���Ų����{J\8մ����gl��lZW�v�z�{m6�2�M��@`Ȕ��:�6~^4�$`$�a�̝��B G��:�.v��ј�tR���ef6P]�=�Cb�Nv_����˄?� ��hƠ���I�����c�j�ru� �/H�9���:� �BVD�b��y� �%u"=�+,u����&J�����y�eJS�;���~��E�i���&6�2��f�E���gE�;�S�|�	�;o�1�p�ީa�'�b��
RV$�{cvW�L���� ���/�ٝ�O���*n�n��5�����󚺊k��5��pI�ri�ŗ���a���Ĉ���"6p4�	�lS����0�6dP�0��6.���R.�H{ʽ��mOJ�U{ҽ������Z�n�/�~ǜ6�V�@���nD�\㘤Ԋ��u�$f����Q9�(V�k�]e��"�C12Y�e���D����o��k���Bt�"�&�==1H�y�iKjF��??f=��g�[���ꆚ���͚h �}���K�A�M�d&��	�:p&%6��d�X;e:ҙ�K��.��	�����Bcx걯�;E��(�����"$�qՌH�����FJ� t�z�������r�emm�[&�ϖ��uΟ?i�:O4Fգ8��]H �3��ʆ����[b���B*P�igU�F������G�XBZ�Y����4҃�9݊�e�붲)V5��ݒ�k&�+��^�}��WcJ?�C�3�n	:3���~1����|�馍z��>+���K��῰V��S��?@@�c�]�ֶ�R�a��)۷oTc�N-V��%W��*d/���gR�3>Ğ�qfG%��#[�ӝA��:��e*�ǰ�s���Fꨟa����_���P�"|5�Pz�dB�ߜ�LZ�Dq�]Y�x0;�?5�V��E�+;mw"�`��ƕ-��P:�A�X>��~פ	�A3��쪤h�[��hQ
�+�2��3���t�Fx��������j�	�=���#Os Ѥ�1,9D 4H�אT�����W�����Ǘz">��
�wH�g���OJg���2]b:?f����u����"J~�׭欪��_]I�����}Ѕ4նa�M�-�
�b/��O�B|7$�fM��Ŗң;�t��*����5r����Er��y��͆���Y�,���)G����|�X/E
}J��;�}G�#��W����eUȺg������&�����&k�+�54|KG��`^���e<�s`�r�V@���)����A��O���\w��j3ӻ��5R��S�y��&ǡ?�>(�@2�شԕ�U�j�ڡ�<��&��t\�	�{� 
�8��Y�z3�����d��D�l��.���\2�"���Z�A���Þ�|-
�۵@9m���E2�t��~��W����]�ģ�l���]�{4��E�7�$~�_�{im.fFp@GE�T����P[;sk{@���0]^y�9�?�d���Y^`6�爞�$� ���|������bD�dA��+��<�@��nH��_�����)_jp���-kWh��%`}	�������c��Z1�҄���X%{o/��Hh�R�9�F�z�����N�#?i9��[;�KX�I߹I�El���"�T����~�3HGdS�Y&������XX	� }�1/'��OM���S�VX[�xŸ���M;� 3��*��a�`7�T�88g�U��ٓ8�W�����p�2h�Ћ��*�
Ke_辖V��H����\�@�<���>����%��v�S���e�`;�4�褧�k�;��j:i<n��h��V�|\��3[,А�ثAK���r�؏���*�6O6�o��Yr�1�����`f��u�s�kE�ޅ�R;��Wͳ4	��� g������ԏ~cQ�*�A�Ĉ;3�T����۲n��Q0���j@�|ǹ�x��տ�W2켵��,� ��zr��'Yu������H�).��jR�80�x(]d��d�+�I������s+�I�T�b��Y�w��j8�N���`�&7��I3~�bI�={p�9v�h��-�kn<^[kO3ӑ�0R0r��s�-�V�)�L�0I�5�����w�:�i����h$�Q�GUw�"!�1���z�������ܙ��&h&�t����E��r��L��������p4WK��4o"}�~v�qR�A�ݑ�G���lp�z�
���:��Q{{G�˒�˥��0tU�H�u56��aa��:JiQg%��	��n�k�_t̞_��&ƽ_>&yG��+��3�}��3�ʣ�! ����o���4�x��܈3�;�$�?A��+,�)
5V��sU��%�IPF�w���j@Ȏ4s?CYH�7��ܿ!DO���#��M���z�+S�~R���x�<�(n-�g�I����6�T�3��Aӭ>1 ��ɱ�u�W���Y�u���O�|�;��A~��z�/�ω��W2��^7P��KP�/��:P��5���v߶ ����Ŷ��Î���8c@�b��y�+���h"t��sq�.�����!��V��<8�o�,����M~k�0ҁ��|�.,^��b6<���OU�`,�_:W�4�+^�1?j~Җoi'��~���7fw�E}�tQaWcT�t-���3��S�OF�w$�!Z�,�h�]`=�|M��@.�J�Dʄ0(�������k���xj��	޾
���lT(Rc[	����h)�9��P�#4�����e�Ѥei?0�q�����j61�q"�n��6�b7�����hm!GYj�P�݋�̏^B8�z+����0�p�!`��$�`�p����}��i�lw��c�k��+�_���U��|����kԠHD�1�}~�z��U?P�.���p��0'����qY�P��&N�S���G�=m1{y�~�L LoA^���;��`�u1?�Sd��>V��6A|gP�
5daܹД����7z��I��7��߿�s�������& s��dE��i�T��|�l��{��J�L|S8�*��K�&�h#=��x����B'��K���]n���~��Eo��lN�Q�PC\X4�ƹ|�H�	�Q�v>�j�%�U�^M���:�a#���8"����6H�|�fJ�R�s���5�b�Ι��>q���z4�[�E�k�h�♪_7�k$����o���<N���0O��"yf�	�6ۘ�Y��Cm{�d������ �|�-p���O�ΠS1C�Ӗ3v^�ܱ��&��9���U��^�8?�ۡ�!Q-��^�WW���{�@�ۃ��~G`9n����qp���O7ۘ�"� VM^U�d��WyZ�W�Ru�������w��Za��loɲ;Hb��2�4D�DҐr�^dlG���Ĭ��Ǵ_ѡOd�]N���ĿN	�{&�����x��3��!D�;����9:�m��}Tq�<��~���(#�~�-N����K�	��uՏ=� �[��'lk-�d�f����Ј�+��B'�Fr�_�{��#���1�E�1�h�E��-�)����1 �Uu�d ��k���NFd�WH��o��Y��ٛ������BP�(��h�Z-y���ľ[4G$�I�u}��T>���犣��N��	����D(�JA8���S\J�9�ý�-�4���z��v]b�z�u.�@�./�aTC����s\��v��q<����L+��攑J�Dc�����W�A�^�"�4�лr(l<��>�U�?q�'j9���ս�`�'ۖ�5K��L�1L� ��*���H��-�E��@�.<L�Z�$d��YP�cl���{��K;�`�5G��>H;�$U|�f�J�o����߸��������.�op�_�4�-i���0�4G��~��>C�)x��:i��JO�`n�����e�D�FY�]�/8��c4$���רd�Ǯ�d�OV�~k�%�5��.x�2Q9PQU�_=�]�ǧfC��fr�&��82�ؙ$_�����O�h�Ȥ��H����M��*���uO~�WՂ辉Il�t�J�}��Xŋ%n>T��]N����Q�qTN#T���h��r��_�H�H�ҟ�3��	/�O|���΃Q:2ē���D:5aF}$0!l_���R�HM��$���a�G��d�nY�29>Q-��l�	�sM����'G�P{�4�U�C5�I��S�{��z���wH-�����	�(&#�硐t7<0T\�K������=�����B A��� �W)�7w���� ����zN@�S��	���B�h�_,ʀ�
W�/�:ŐJ_�11R�j#ւ�ޫ�W��0���Nw�"ZI%-�g���q�COp�^��:�$�h��l��J{a��|����|�Z�3F�?��զ6m�qӢ�/o��1:�N)_�NĹ]lT���l���1�6�"�4Ӟ(���z��;�"��v�H�Gj��j���'.�W7�&z;ծ4,���/�
���05��7�,�3�X��V)�b�*�g����~=���.��BUMb�ev��R����)u4�ěr͠19�z��o��
�"�	��I��As���S� RB���u�q�q<e�Nsl�
Bo+�~��,��u���z���J�N�Vm�`�o@�m���D&O؎�n*��U'Y��2��P��K�ў�>D]o��Tv���]�]sD�>w�=YE���-C��h�U<^��b�p���I�Ö鑴���I%N�/K^b�Vgp3t�pL ��๿8j�7�S�dN��e�F�y�Ȍ-��[+Y6�
#�iP5 W�LE����c,៑b��w5蔇6�Y�,�p)��8u~cq�%��o��
�z��W�E؜pal�rt0�[<���q�/��d��{&J���ΡmI�P'��~�<D#�0D�5]��!@x��C�Ǆ��Hwz��ʩӁÅ������+�J�7 i1�/t(,�0���{S0��'*�C���n]�@��NO"�:	r	�{B�s��(��:�uB��W��GL9��x8O]l4-���>��=b���.��{Oߓ�04J܄;F�0q�["vc����l=΄��a8J�&�m)������>��R���RM���6������,�x����`킒�/
�D|\j/f��L�~Jy��P�*������=����*�NѦ���BI3~�$b\��TR��e�!�b3'�~+wB�.N^Ws�4�0���2G�C��FjnʗfHf���N��lwMY�f����r�xG8rH����^͸��C�CZbOI��n�m�����PA�MM���U�<rOI����g���h�7$Mu��	x
X�v�����FkԘ��~�ӳ@��H�N����ݓ�z����V$����Xn������0�[T�X�ٻ��F#U���F���tg''��_��)�{���s�V�D�wHV#["�U��.`{D/�_@X�=�EUn��SW�Óq�>�3,�޳A)��à�ܦm5������MMSB�gZ�A��_ڑ����빸���xล� P�e�ײ̳�Ԥ;��)[����m�>��J�cK����u��I#R�qWmgڻm�.,_�N��M��t/��a��)��?[�|z���c{�R����*�g�2��uE0�[]�[^1fv9�NQ���Sʣ�w���0�tT�pWx��4��ҁ��M���5�<��{Ia��x��ѽms��+����m��i"��)́��5u5uL=���~m���kk�/� �PR;��H�wygoIr� �CiѼ�'��[��+�E��d݃ru	>����h�Q�%Pe�4��T��֑
��e���=����{���th7�E�m��r쑜�a	iq��H*�h�۷p]��$j��w���390�F��m4	��H�$�
��m1s�r�����ͫn�d��Y�$�%} I��7c�Ze3��;z5|bȝ���ƿ ���XοB���=�[��"+���mv�~�c���#�)�ra8G�2yّ3�H�S[͓mko�9ha�v�#q�'[��E����ޞ՝�Iͱ���X�"�Y��D!�q)�@Z��`N��c�9s�qcc���b�B�.3`�K-�b�`����HH6u�^���m=�/�@������y''v��k�w�|������Ma��Q��-5��ʶ�8��
��됢�r��Y�͚~��R�Ǳ;�����C�@W&��Z���`���%];��z֒7x�˕�!�
Kj}����2�M����C�:��~��`�&(^���l�`o;����p�,0������q�mފ]��D�Rp=x�'�{cE^�DOL'��b�Oė8E��#�<�ݒ<%�V�A�}�ޫ
�'���3���?�{ʰ��jF�Jp��L��7���Zg�A�Y��v��v`��5u��nx��I��P7R�%�<H�"J��0�; [	3�����4�۝���@��?yӝ�-誊c_��<��j��Ki������&�����\���Fa���G����"�!qz��̓b+G}=��)�� �zvq����u�m�f��$4N^Y�r��e!�Z��`,�NIe�����=�� ���)��,@m��j)>�|���p������?�y�1j�2�y���I�X�x
hgL�19��`}�M�+�l���k�%8�	��������ώ��9
i#|�Fy�%78�Gg`e�
�T�x����/R�f'��]P��7?�u��կa�炊QWN�����܎H���ڐ* 		�:4�'�E?�{�y�����V-'�p=�N��u?=���X��O�Kze��P��v�o�p�����W��=�=F��*�\������l�H�}��s��3�hJ 0��K3!ſ`��NB5��⒮�3�1���kŲ��X��h/^�{Ӌ���(���pzL�a�{�wx\;ic�S�j�~�9�z��u��ɖ����~�U���S�7,�J�����xm�jf���5C~X����f�D#E����,;P�$��z�"ӭe�׉d������}W���(r��2�=	�5��g$;��oM�ZAr��d_$��	d����4<�rYnk-l��Ч�;L�@F�c��:�tc�'d�pj�L5���]�h�$�ǀ3;�����|��S�JL�.��9/�*��)��Ə�e�b �$�sg� �@�@h�_	����:#��?�<f���9�2��
�G��y�I�1"oPV�)A�?̜����y����P4AC�?l�Mc�h�?���)�+�͠�FqP��V{�����L
����#XD�]V�OY���lwF��R�GK]��3�2�)lB>�����,F ��Eݥ�@`�oL��e�q3��v����� �8(q�h����|�= ��S��!'�fH� U��)���������Έ�Z����ڜT墍��).���m������r�����Ht�K��O�닣��ZUH��_��xе,̐�/b�����/N���_�����yҦ A=0�$�3�n�ԖIDi4y��l�v���-*L5�*?s�q���~jwZ��d�E�X�-غ��lJC�gvz��V;)�lӂ�Fha���K6ا����=Nf�=��4n_@�\�Du
�!�}�p,Q���ɫ��J{�>4������O˭}^ɽ���B�I�Ot����F,��C�F�̵�������3Buw�=���m���K� �����Ό ĆVhfL7��4鳭��7՟�k'�n�<�d�e\�9o&f�|P����8��k'����K2�f�B1�6�$w������)����h������n��i����$�-X� �� Bo	%�6Ė8��:Gn�vT�k���Pn:^��%���}�_vޤ��h���U�jd�Y�S�,����P(H�������ƍ7<,����>N��O%�Ţ�Ze�QR�$����n����pC�(u$̽F�N�g�Hj�/�(���&ѝfMn6B�p�;T+�?|܍�4tly��p2�o�<R�z�2�l�Q��9��ͱb4����q�d#(\�<=k�Z3[�����и�NŒ�)0�Yp�rOV�Й�*.I�U]����]�eSx�a�1,GK6)&��F�LJx�xa��ȭ���
qĭ~)�-��aq�#'|�'�:�
#n���у���4}s�]K�ލ��0u���Y���c:�$�Ƿ�@;p>p���A7�.�i�e3͐ZܑjH�W[wVGM9�@�ER>�.~���Ǖ@�)��;"��A��6��v��"茊���#�m��Kv�:����na�9�)���C������v�4������Y"�|�_�����7t�z��"m�47�f�����f�����#�S"�t�� �1U�.8ێuq�	�(��&k$�0n��i�58aߏ9..��V^�:x�5D�O������;��/1��������%U��qZ!��pN�T�9QJV�����QX�"��g
f��81��E�ߕޭ	�f�~�Ue���t��]�� 5� ��쵤�ߦܳ;�xX�aQf��$6�zj`N|�E�Zi3m��ْ����X]�%j��~�f��� !4Xw��,�)%���;�+��:T�����#뷗*"̀lu!��ֈ�v��)��9-��2��oMg�<�'*<�}|`-��pw��S��n/w(x�`.�H	��含�n< �
\��S��g���ے��@��9���_Jd�<�nv�L�d�	�j�և��v"A�B����U�
�Ha��0d�q���58�����|��?H����0���S7`�՚K��ib��<�p�E����Lp�l'�X"��ĸ��ӗ����"�)gb����OnΨ1��@��b�,�g��^	>}(�b�X@L8f�d�̹;a���,�/�ޥ, z�Q�Q�.�`Q�dYO��L�D���mr��#+h�Kq��:��Z�����&��=m�K�y�̉�}��l@�Er&��8�V��!�����^P ׌L>��O^�p�G(�Ml�A	��Rb���$�[������ͼz�ib�[V"�7Q
P)E3̡��#��P9�_u#��XV��h<�
R��=R���������/���*_5��_�Fs�o��aFs9�F�èH�n-����� �d��T�Zu��	\\�*y��@����e-����٫�V�]d��%DQB햧�0�}u��l7~%��r�%��F²[f!0�;�7��_*���Tޝȋ��\���a�`p�����q��(�=t0({Z^k����	�J�|s�x8���h��G�˴l�*��y+�H��ʯn%W�+q/�I�o����I��+%�Ȝڅ���$*����8�2,5���U{q	?�g0\Q���	�A�:9(��ؓ\���[Qf���I+�a�]bb�_N�CSŪOp�R#�HI�=�����fOl4��%!���a�^����j�26�v�>:����#\`q}W��EM�tޜ�Xj�q�Rh��Qq��*1������3� +>����+<)U�5�hޟ�(�3�?�ܝ�vΠ��5Z��bo���s ���j�	H�����c��NV<oKe�pс-�I�u���H��M6L����I��t�[_Z�J$�f�牕\���j5��X�Q���񔫨��:��P65�.�\���Q'��#��;r`���x*q�2P��\�z��#�!��c����6�6����`Dx���@:F�_L�ȝO; Ȅ���FmN�W���^%�nv�`h3.����H�F����s�z2���O�$���e�k�E�'��,T�	;'4�䘚h��Χg^;�k˵\X���w�L�xvM���z������=a�68bS�A�br�����
B�K�*���~rXn	w��W5��Uf��\D�ӦH�h�b5�d2��აA~Β>��Bѡ�Q0K�Gs�-���&c
�/p̔M��6�h;s���Ta�A�j�ڀE�>�_Lsa��'xGZa�ӧЃ8���c����rMb%-��O�muz6��A~�Is���=����A�H�W;Y��M�b�ac{���8�U�U�.n��O	z�����.`=��C�d'���A�i�'{��I�朙�՛����*��!Q���zi��Ú@���ہ<sngH��^�
ڡ`�<uܹE��(���-6���'�**R�)(9���79�jޒ'vx���`�)�:�6�9ATÍW�ŀ��u<}�o�������E�D���<��*�e��RK$�8�y�a�x�e�\���pVK4����E��O�u��Ɋp�m*�%0�ewr���4z��U ���{R-JѤ�#O�^Zs���f�{��4>2�D�_Ա;���&�}YX�]�����`���ַI��8n��b�'�z��l��**��#	��rqɖ(�hk���5h�h4��ϟ_JJ;�Q�,�����C����qe$�ei��-FS��lL\xIj��*�{ݑ��I���\8Ҡ+�� G�m����hǇ�M��38�t��<
E��D�-��B�L�Uڝ�
9�Qw����ԉ��ƭ�?�n�X��O��m������/��}�:��o������l��=�jᝁ���k<Š�eJ��}h�f��,�ؗ3��)((�\�t��5ۼ��8?f��*`��`K��*�=���f��ݼ�kː���	�B�G�Pp*$)t��⳦�ٌ��8$�!�ͧU�(>����Y�E�l][�)4󳓦�#���#<[67�'�V	�B�j�w��=AzP�cN�g��K|֠4�ſ�6;��Q�s+��$ u�3��,CȎg)H��'�)-�P���-Lh��%�FH������,<�Ч�r&%�5w��������G����4 ���z?ϮVD���"V&��}mԁU\���Qh�å�ʊY��il��9Go��L��+�u����0����)�4TC뜜 IqZ��l5�0+J���]\z���`��GaR(�9.�7�]F�%2�:�e�v>}�*�7
���8���Ӗ���U�(:���#
W�åB��_F4[�.*3ڪ�IJ��fHM~T��C\Ĩ��8�=��:�dp(�H��8cO������}����W���u�&XW�c_�k��ƭ�Hʉ�@y�7̣y���o�Q�IM��Ԥ�n�R��Q�����2�L�G����Bع�*z�c ���\f`a&�n���/��O�O�PrZ/�6��V�#~B^��\�#��`�Hݱi��*�@����?	d����\��'T�Rߩ���Ɯ���Hf`W�+r=4L�NU'��Q�&{9p�:�]����;�ӆ�[���/�|�.[Z9Tʭ�~e�Md=ȿFϵE���Z�W7= l[BE�D��i�w��"?�y%T���vB���W(|�}u�T�5�M��u�"N@Gp��a�'8.��1���� ���_�s�R� �����i?���׫�O�,�9��E�2�кD�4 ��\�G@:�I�A�5KFؖ�s׌��R�ϲx�x�F��jo���%yes�5`�	���:�U�cgL7�h��%	�I��.'��a3A|��hy�6��K����=Iw��y�c�.��#�y�bf��I!�덚g��iR(���?����`�{�fY�5�@}��L������ՆT�f��7�-yR���ԁ\�O��}[{��a��ZaK�Md�^R��Ծ�X�:P���CW�����[extl	���U�K���$T�um�	&p��B�ˠ�j?�Pt~��O"�6�g�=�xD�0�]��&��x��ǬkX�{�g�{c�d��ߨ\����> �q#M�	���#���,�Z. �_���2
��(��r�U��`�X)׉y�?|�9�K ��	�9	닞�t|�S�����_���� �.LG��q$�|;�E^4��nX�� q4p0�@1-}�����a�U�����!�o�8�\��	ujGy�$��_��������PsW̪+����E�iG�rx|�S��n	eL��)����})��=k�\/�T���3��r���o������,?O8n� =��7��w��B�o!�[��J�:n����i ���O@�ْ;�^�0}F��Q�w�b?��4��
�m
+0�g���J��<T
�˓�g�f~cu�V:]"a=�ʪ�*q��kR-�d��H�흌�v�����h>�zG��?��D���]���|�l����:X	�xV�*�M�n&e������\���k� �BNp�E��G�"!9º3�s!p�h{�����6v�EБ��ʚX���������O�t�M�kn��
�}a&�*��D�ؼd��o�v%29rp���RP��	>ۻ(�=�b�.ܤ��n�C���ݴi���nwm���6944g�pp�J ;����T"駤���_�Q���Z�|ـM����
JvM��ź�Zvn�DA��4��H����IW�|�o~�M�;�4���u���eyn�
R�pO�q��'�jNw�,�H`Q�6n�m�c�^
�-@]?��\���p@�G�b�[��C�q�+�T����Y�+[� "����%��>A
,	��8i�~�T��!��l�)E�H}����΋��P@��߰�G:�i�����#�A�2s���}". �y݁a,[Q �q��",J��."w��0�xL�k����n�����JN�}Y)>�"�:R�����VM�e[�gjO^(�4Hۑ@������ر8D4j����6�U�M�� ��ZoG�'�g�ī��P^|��K�Vm��E��T`�>%_z���w�Nb�n$˙1(�
t���~�Υ��03W��X��miW3}%��!�����t�*��e(\T�"�� �K^��\5.���2��6`�Y� Z�ŴI'��R�̟�E�>Ҥ%%q6�A����[�{M�nW&}]��e�I]�~��DRԮ��T:M�l�.V8i[�´��ס0�<�豘�f���; K�_�2�O���

`����a�!�������3XJ o2K_�i1�HGm�<0�y�ٰbU���n3�Ul��u���eWx�<&���jR!t��K���e�ş��t5V?,�Hu�HXD���q��7�	S\q�j}EB�ᡋw:%ZO�=c�ƒ-��9ĚF�3�.m���\6�?v��Cq�Љv��B���dp,Z��qላ�{z��Q?gtWNp�h'���U�x�ƙ�e5��ñ��#U�3G�۱��������j�|�&��? Hw�Ú���T)*/����v�
��V����G�h�+���)-�Vi����%�_0m'�[6c*w�ɢ�)��iz�*D����w�O����T��������z��"`�>]1P��"�\���=�PIo�ۊ���X�^>�F��T����ﹷ�g|X�PE:��]�UY�jӸv����W����Q���>x���fн:�U�{$��9�U��?G�3w��x�T����~iZ@<��n}���4D��W���0U߾�
	�,��gmP?�ްj��(G��cۓ��*�����!�5��X�ea�e
�OۖJ��q���� �h�)U����g���������`2F��ۉ����-���[���'�4jB�{t��r�Ze�/P�:���Ā��|H�8Q������b�j7P� L��&br1G�j,���;Y@��s��;��c�(�?t���.<���8'�7�(��=u�g�ǰ�\4ڞ�%�X(�bO�v����⪎��~pD�ap�2 �tl�ψ2Uf!�(D���փ˲"z^�Y6�QW�\x��{���@�[�����u�B�D.��}�|����5[�j]��4��L�v�V/`F����%����4��!'�I��sh���y�����3w���U��qH��R[5�g.����Ʌ���n��W��>�g���F�^�k@5���s�t���c.�Pu\K$��b�>��)��"��X��ĳ��XWFL��}�I������!G!Q���H{a�<Ki4���֎N��s�X���'�1��N��4�9���G�(��y��K�7F~(�������pf|�����6A�R���0�2����s�6W�AE����AM��04��  '�×��^v�^S&��}���� �n��$�s���W ��$��.�hǧ��������tk��X�zQ��T���|?�U�����2�kvk`q� �(�k��"13��b��!Q}�Z.���� G�c�\V���&�TOGh'gPQ�5�GOΓݙۏߟ�u@��4���tȊ��I��W��Ӳ��l��ݠ#l��A
����P8j<s�3U�Rc�$_ӟӢرͫ�����K[vg�"�?8�ho��I�H���wuFJ����#o�ڱ�U@��Զ]d�4�A4�AbY��\w)Df;����w�w*o's��މ0u��5^�س�&Z7y���W�^�@i�i��`��5��sZ�}ɽinG��>vTˋa�r���'Ta��ը3�_b��Y��y���i�%j��˓"�8*�|����#�U�"���"*ø�LRU������?�F�
@W7/Sn_��ݔ]�g��[ʌt��b����b�-D��[_ҳ��	�������5)��bVW䐓��A3ؚq��֤�y�ʱ�=�Q/�-����F�!gq�G�!I9�D<0�����TB��I��02��t���e
����f����"��b�}�>1�@�8QS�qY4?���ٖLG������*M��1��KI�H�E"wA�ϖ[�bO���h	�)�1S #/ɞ�� AĐ>`�6��o�SbP^�N�|�U��!��(|��"��n����Ɨ�xp��RD7����`���r�K5��_����M�^��6��H���0����m	B�u�,���Α�z)a����Dn\ ��-Z���WR���1��T�W:HA�eB,��S�黍�o�FK6�c3�%*�F���2�3��a��}G��9�z��������P�d�9N�>V.�E�0���.S]�����m����p`t	�@��f3uns��2V��}Rn�Qh����)����Խ1f�0�&�xMϲ̃J�2��i=�5������tu#]	��b�2�7!�pv;�Z掄�O��颓�rU4�Q0�z���S�d�c6.1��]����O�ؚ�z��2�ڐ�@�#��v�J;ȋD�a��uN:5��w�z�S>��-
sk�)4�<dN���vQ���_��UN�˦+7@�s��XB�C
�a{�����V���EŞqL)n2���sa�:67!2��9.���[6��C))mįT�VB�bt�nl��
n�ϯ���YѢT=&nXHʆ��p��l�{��O-�#�O![��mi�+j;���J|Ĭ�&wQ
`H�ؼ�wx� ��%	��u+"�8�]5�3i<�\A���)_5-��LCH��>+��|�C��K�˒��>��� �H\����Q��i����W��ʀʊܛ�m�;�%�a�P�NM����A^2���-B6]U���RY�7��N�R���ћ���X�,�	'F4T&��@_�5��jf�F�\8��rSh��馣��3M���o��ѻo��*��t���r����tu�i}
f2NQs���R=��y��C.bi.H��#�cC/:8��O3f���"	��]Ȕ'ʊ��'ɥ�#R%�D��xޅP\�0o\or<a����P�S�ư$���h[1E��s��������R"S�}%8��ލ��4���	�f�2)_�o\���,n�:�9s��M3/��"ߥ5 �m8����v��1���pN��eh��6�W�
���;������D��M��0-���*�B
�<\��ǻ2o�����*���g�|�J��K>�4IeN�	#I��Յ�[�Mu��	N*J��D�Adg�Q���ն�'����l���%"H`t|sB���6T�	��T8=��=��j�r.�0�<�@����>��PUȠA;�t>Bh�mF���9�ada2cy�fj�e3^�?�eM��hAߓ����R�0��x��k)>�}��(�֐'91C���/*��t��: ��s9�+�N>�O���Uv��,�#?f��e�JlB�K��*>x3d �>f�η]��7�Ư[��ʀ���}m�聆@��+kJV�WGma����`�u���L"��3�h�V�|'���	���c�, �����%�L�ԩ����}�����k�2c)!�c${���u�݋�MK}*��fW8plL�*#\D�ݳI��h-��s���_�v ޟ�pnkQ��\��A:#&�4�iZ|V8��{�
E3���[V���Y�;(�I2�u�Е�s]�72Н�6u�梫��-~$���'ӎnr16 ��'"��8��њQ�s��&��f�$!���!]q
lM,���V�'���5U�c�CVk��y���[ňx�۬ҧ��J_���э�ǈ�qk��ցM�� ��'F�=߬�<7%:�ʝ��#V��z*MP��~\���̴Vl���9t.�W|��' ��B�O��������&�zmE���=T8��ҒȔJ����G�[��t��*gP&X�,5����=��jd$Y(�q�L:!,�ޥ�H�]_��W	�*� �ȏ�.���2s�9�LY-Abj�v��֋CeR��mpk�Q���)_�A��@J�9zt�;R�ο҉2gI̷�1��Zҷx����wdI���]sz�>}���/d���)���c�'л�V���Z�Lzė��OY�n���JVc�N��3�$���?�,���t��V�g%>5�3j1)+����6�]" ,���.=&���Djm�> ӻx[�Y��F �C�N+c�P�(��&��'FJ�ܜ]C+x0!�PT�ޏ�eri�3
%=;��*��4�4���6rt�F��T8E�����q�Km���%���Yr?�zP�7�c\9КH $�rS���%c�@��9��ʙ&�7jl��>���H�m�����LH�\I��W>ֆ�5�!6g+��/F�}p"��,	Vg�w���טEX�n�b�Bx*¨Y��V4��!��ȮxD����l��櫌���U��Zq��-�-��3D�����ʸM*�Fm���'���k��I��䉖�e�4�QN�}?;0�����Fe'��ҭ���3k]"��k��S��W#���[�~��c���{�Hu:���Ig�U��Jܜ!@0�7�,;���!������\x+6��Oi��یu���q'!�b�E���ه�ԓ�O\�:��YqiQ�S�ʇ��7��
+��_�lQ1� �	���#��j�������ds�#J$5Y(�b���s�uw�Kˣ
Z�nZ8x~�Op��]��?SKUK�'Hѳb�g{~��� &�wd���DOAl��=�s��0*m�6U�֟�J�n�0�������.۱Wܪ�M�$PD���o�Us�`+�(M9�k=6@�:��p���YT��i�+�S�Icdrq��ѕ.'l^��I�R�� ���I��W/���Q'��ƒ�v2/�ɫ�Y�Z/Դ�R �7�$�ŋ����ɾZY%����!�~-��D~
/w�&�D�P0x��6��g���_=�!%��5;��㕣k��KG��VkE� Ư���d���=x��#��JSz���w��j�$4vF�H�����*�
�0�Jb(�h��|��>tE��غ�|����;��8i���}V�r��Z.�c�ƀ���9�T����@Q�3x	���T�]Q$��8�[ŀ`*bfKȜ�SJ���U\�q �}�择�I���;�ޱK'��VEs�L�S�2�ҕ'���6Ͻ�y�b-�P�$�o���P��6���Y*#e �O8:��ХU�#�:�Ƭ����f�w�����V��^s��v5�C��wdF5z��.._���kڒ�������ķ~�l�?��@C7�2!�ʊ��}Wɏ��������a؊�ְ�|� ]7�$�vc��E���IQ���!FUȻCֿ�� ��#7�0�F>+���֘�A�[e��#�\��cҔ�:�������}S:��+�0#�h�{c�.��m&17c��$�Gƃ_A��^�Klh8=�]���w~��HQ�E��6���X��Q�-hJ���qiI9�r�~⸶^��e��|�5�������F �e���c�擳]8!��ޛrW�6�N��-�����gD7F��Ӽ�ǭ�m@����Q�H���:Е��=CJ���8��&�eD3l�ݽ�~0�;B4��8��J�
`��d��r�'�9;���ے�#�wZ>�����^/Ш�Z��PBL�,���XR�^���Z?��}�����z�⍸_ٕN�Y�6M �ƺ����'�
S"�HǨ��f�.
��hW�<
�w�8����[is��o��w	(��w�3U'<E�@;��c�T�1x�>��$��=|��X��$�ŧ��Ė=��o�S&���n�LR�rJF��8h����� �Q2���E�Ȯ������9���̫Y��8������?N��_�v��J�="T��oא��b��&]4�J�6��P�bp�^p8k�lڸbg�r$�qi�<�;b�7���Q���`&�r��b> ټ���M�!sl���z�ԜɎ�պ��z�1YpQ���.,�:�/Q{��
	f3�3�GKa�A$3���qs�9�5��|�f�)�{�̡*�(#��#h��im�HC�X�3x)� ��v$�WJ'Q��Ы=k���x�v�7�3bq��QI@��5�Z6R˃�����̰ʲ��sw��r�Ga�׎
��#muyR�]0W��a�������;�h�����U��[�6|��穒���qF�j3�&8-�G�,r�*h�/�;��X�>�2���ЭF@n<_ީ5�`�=*0?���!����A8�����rz?�T�c�s��Q���_ �/C���+�n�S�3t������)���e���MÍ���rq;�K w��$ˤ��^����=+p�&��\KZ_�Dc��bw�K�:|��Ǝ�jS�-���r	i'H�ԋN�րoAs�����ɳ:��G�'�U��X� ����������iC�4�T�쟗9Z��ȓ��Dg���z�"�y,��Z�p/�*��c���ObQΐ(7� L��ZP~84dz<k@�M�=����w�»G*�P<<'�E�ˈ����2���j�Ϧ�*{�S�ecȨ/��J:Sv��B�M@�s%��s�:�%���5��q�U�P�g3I���lȑڸ�I{��L$���٤-v����wt���U�#�S�S/�E�K��>#�u�Zi�D׭��AG�P��B	i�X2�����1��E6��Ԍr�[���L�2��+�qy/�s/�<��g YH����B3cYQd>��.m�L�C�X,�$�t+�1��"L��M�+[[j�a�qB?V��Lȝ�� A��P��
�=ط�8S+��$(��ߺ�DmEx>������]�Z��jg':�m�my
��Fa9ȕ�C�7!]6��D��H� ��ǡ��!�SŐ^̔�΂�NX�kN/u5�BY���x��g��L�C;�9�Rsx��<���������o�\��k�O��I�q�^J��h��.����bV��m	Y��2������5:�T�{+'�AR�Zϟ�ٵ7F��N��Vڕv��ɇ�rw�*>����+�"�>��rJ�Q�RPaK�?�O�F�5���pyM������^���b/�}X_ShI��G,�^��k�[�|F<Ά`.ܽ�hqq`������A)�!�>#mK�vĂ��[b��z��_0	�.�ӕr��������B�UJ�{��}p`3;���O�e�j@���������Y���lT%��ũP9rv��;�	�����ya���&�U������Ʊ����n�d3�e��j���?܎n�VZ�Vb���zSԧ�+�<��L�e���+6��_'��l|�5:��WV}���=�]�Q�<�y�4&h�>����	��m�Q
s��}���V`ywC�����2F��R�S҈~�d|0*��V�勊6s>WF`�0���_562�B�@�}��۽�V���9��])j��"�Q��Y��$=.X9:$_b%{]�t��@�>^\؇�|����'�g/��n��e�_�|x�a!�A��'�ҸJ8	ǽ̉�y�H��3�p�`����)BJ�^'�l�8h��?G���8I�W�X��Y����f�6������<W�\9B�n5�o�8*N�rW���`���m�gCH��t=GS�o�R
L�S|zn���y����]��3
 |�ﺎͤ|o�Hy��b�.����Ǿ��Ҙ�f���"ӛ�/��%�����ب'Q?f���Ib�'�ZG�V��hp�ۓU�K�&/SH�Z[&�?�а�5�����fy�Ah�͡{/�ߥQ�`�BcsQ�����㽁��bԃ_/>)#K���&.oR͵�v�yN�(O{_�r%�X=�z��[��w'��L2K���*��ыnw$�Jh���_^�B����_�ӌ1}`��j������_m?�V+��g��sr���<�qsf�k�7_�B�jF�[��C��e7]��4�����Y�kV��c�bW.哦��h5���:�*��i�L9���/�S���9����"�5�M�o4=D]�'��k9��ɹ�{�r�iżsR1�
?�)C78��Nuؾ��Ք~(� �/3��#�b\�Hc�N�R9VE���C6E��N8��i����668�헍�U+����W�c
M�s�\��`VQU�Y���~8Iy������U�A(3������x3 �Y}��:�2V���M��T~��w��x��ruF�>)5��W�M����:")Qs�i��D"�Φm\w咟�H���6�v��U,*�,�#�q��sXj� ��e��ݯ���u�:j"��e��#���@��}��OA���ߥ��į>�T
R�����8��D�,��y3��'ȯz��q>A�B�H@a�kh>�Pz@��ϝ��iuё�;%"G���Us��iL����JA�3g	�',���h����n�ę^�B�\5K�YAT5���A�����8�1zf=u�&���jޣsKd�j�W]<��h0�$͌�^b��qD��n�r����J!4ުaB
2]C�ы�D��$(vM6|J@���2�g.�Jb<���R�V�К`�kZ��!�g3[��5k�u�+p��{��6��'N�h�� ������^ƣ� �|�e�w�A3�y�K�����Y��q=U����*T_&,�a-*B5p�Vތ�b	�RT�oU!���w�7?�Y�?d]s��r�47����(2*�wH��IB9KI���O���"��gh��=�n�G�?��}����u��8MO�u��!�K��$�a�h�q��Sy���l����k.�/�����
�4���yh;y�B�GֻP����!�@�JMע��U���ے�	u(�ְ�,����W��h��@_)N����h�a��4��9��D�=E�7���;S�H����D�s���^!��>!�g}i�2j��o=�c#0#8���T ���͐�Ǩ� �t��9��S^�>�]���sxXW�,����_����F���)��"�ű��G�.s'��rv�1�xiӞ��t�=��>�qY+�5��@�y>��C% �6��.k;��/.�%������/'m1�Y�9���>ۧ�'��F�s���ׂ�z,l6&,0V�ǖ����[�����t��<q	�t�8��g�������O��5N���6���5\�!T�,V���l�9䉔�#�r�HP��H9�ׯ6�$�Q$V#�{9�R�\�������6� ����<<L|��n_���H�t�3�������Ұ�#�k����!(���(>�2+�#������F��z��k֏��nG�0�gN� &5�hL��d7цv���+AD̼)���a:. .^�2��v���G��ǹ��t��tm����<�a��
@/���	#��㿡Ϫ$N7>���6O��k�M_2�Mz�tU�j,����qj:��5�EHu����Wka��UU��y����X��҅r�śt��Q��ΰۢ%)�Ǚ�y��r���F�g��ʳEy=�n��N�Yb7���!W�u9�/���Y��-�u��� O)߸s�=gP����N'q���Qb����[�+��JT ��2qhc`���6��KB��Z���|9�5��a�l���-t�u�ע��tOO�{��e'��\�jw�6��0Po�D�����1�[%��n��m�h�-���Y\%�ϲ9.�&��o�k�X�������"d=:{=_@��՝U�`T���/__�쎗X^��u'v�<�٦؆�]�A���ԡ�h3�t%��S)�cq������Fz^@�N�#'E�zw���|��{��)��#��D@=ƛ*����C���2�sn��@����s���-�KҖ�7�e1��]	�wڸ1*3Ieps��G��tX���Zv��(ilھ(�cz1���C�[aF򨞬�~�bq�l�S�B�NCS`���V)c���AB�Wa�Z-�����:IP�O��Hr�0���a���ż��+Юza��R��ax_��m�Rk(��N2*�%��z\+�������`\�xy
�e���#w�7�g��gL'�(Oݗ��^{��7!:����;[m6i�D*6�������P��f.�R=�l�`�se�'<�u��L&#NV���W�r���ܝ��yo&#[I��;��īɬ�AQ�)V��K�/;�2�����#�?�#�<T�}$�"S �`|ԭ��7��e��V�6]��^.�]�#��8ZIgr. �0�-�0�"�C ���+�a6�����@\��f^4Ǐ���uT� �������+j-�u4�D�q���'�)�Kw���p��%���$�/Z��K��M]��U+�:`iSg��^`�H|����{)z�f��Y���ҫ8SQ�yQLA����a&��;����x~�9qE��ⶼ�{�!0� �J��б���Y��⋭���N;+�0�o��:�����B���:��ڥbS��h��ۉ�^���c�H�Y�����n"R`�� @�:A��Ҫ��X{��e�?1��*�s�7�@�f��(�������X�_Tv:0@��ɗ��cǞU\*J��Umm��;�X�p��ф��R�v&V8_��ٖ��
����$"0 � �}���zBr�Ot�^PU��X�������A��mt�w�x7p�ZJ��&��{������5����m%�߂2�o�o�z��JV)ԟe ������� @���������Q���=�z0��oׅz�J>E��-���1;�bU1W���Y�����e3���CӭO�S�tY@�@��B�F*R�HC�.��N�2zZw��n�F+3ۘ��2�i ��(n��c�+��6#t%�rR��Dܘ�U(�~V�{��/@�G��a�Gd��Q��L}�j��\�x�m��}�'O���[#V�5A(�I�5��h�Ck�l�EӶ�I��DDIv�F<�@�]�O�0V�C�tn������$��dQ���h~���8����#�~�T|�e>~p%8/�mh�$r���"<I��A9WD��.��A��aMa#$�O��2�d!����D��_���W�4A�v`&���,3�1�B��ў*��RG5A��V�y�e������6}�u�%D("����Z�7px^��F@��z��<����R1�h�[5$Dif��+I$���0=�D,x$@͝�6ҷ��wrc��ZRÖ��te����jn�����'�{�D6���_���s��2�Q�z
�H"a[�|�����2kۧ��r�Y���K��R,/��֣����LFr0��W�9���)3�C�^�3�!&`����[��A���q�p�G�~�'<���$��b�^�� -z�D��1�I�?�.i�8����5��3hߍ���f٠O�����C]>cjL����.i������σ$z�l�I�oL����+o�d�C��g=�כk�E���I�=�Z��W�V�0��)��+0�O��9@���T�Z����o@�z��\�r�MX"j#_�%�A�I���A���t�@-���8��'l/�~?�c��Bi*�8�,�V3j����o��m�c�T,��H�*~R���0W���-_֊��d�Ņ�AyL&L!��q�%�����.W7ElG�b�/Ϣ���ѥ���-k�y��0���W����[��3��&&C,>\,�g�>7����sz��RBZ$�B�c8���k��d]�Q��˦tǹ�|�!<:�,��`Y�+�o�,BW;�{���#���_q�4�U9v�����@A��%,^Ȯ�x*m�nr�-!�8��Ď���,e����ժ+(����r�|㴏��l�)Bn&-�9��w����p
eZP����C���90۸)�^g��TqK��9TM�s�]+�P/�����y!�l���mUX��֌q��XH��![�}� ���|;J@<v�vm2��X��NwC��*�����?���F��-^��j�A}q<wq��d9�-�j�j�(G��Y*�2g`�J2�YҼk�8`��l7�<ijj@���50`�Ț�p:��R������"�B"�U�/I>�{��r��7�Ż8/�}�|8lW\�j@�8�p��ΓU����jR���ڌ���{m<���ґ[�R	�SH�2�Q���(��S2x\���Sg��O��O?|���{u��:�<�(�Y*�Q��b���S�s�S����Fa���Vr��BHOE��-��W�S���o��>�.�n+.�}Ua��}:ǡu3�ݲX:����h��x�w:jģ�:ȔQ9鯆X�5��v�n��RK�d��y)C���N"����i<���xy�D\�"�!VB੺�ǎ��
@#��N����Dt[�W��X�����P��Ǻ���o�p4��%���92��V�n�|���ղi[iMq��2�<�s��(�-OmԙY%`�EnV�[��̍*�'���c`�	0�F����jp����T;��5?k���i��Sa'ӟ�;\9I6���!�#�q�7�u�qӣ�=}���g��Ƀ臟a����~z�O����u�����%��& ���hN�k��9� i0Pd<ń�T�#�'���&�i�S!"3O���" �BAu[�Z��1a�?����%��eߣ����k�e4^Ɨ.f(2%/?�Ο�!k�C:�c���$w����1&��V"^)Om
�7y]9r�w�r��(�3�$C��� �!�~�h��{����mZ�B�Dl-э��G���ΓOt�.%C���^�rZ2#b�b�t��Eͽ���tO���{�~��v����"&S����&?�*�#_���<�g��Xz"��O�Q9@��\�0 3	��We���v��_A�)��.Dx�?SRp�l���Dbf&�5�L+>�-I���1)'z��t��n���a�"-˰k<J#��\7�������s�f�zR�saA����TO�k'mF�IC+������oY}_��K>w?�r✓ƩU�!-�k�P�<7,�ּ)�G��*����[� ��b�"L�U�s�.T�8�^���F��Q�k�I�+w$.~h(�rÃWO��:O�>���Z�^vv�SH(�r�B�BЃfT�p��O(�3Zp�ܞ�]�+�2��R��A���G�2�͐�3j��f�'�nC�+�%��D�}�د%\퟿�N��p�q�wL��41p�}���s g�{Cݶ��SJ	�X���L���b.P��;�i��˔r�#ԃ��NM�׋|(S\��Y�"SKҶb^�E�^������nZ��_vo�_��A��+S��6FE�o|����?^"a�j�	v1��2͸�/XMi3�8�P�G��\k�-�
��r���d�>�Ic�z04���������5�J�ڠ��#��n]�?�c*<0�7F����[��9-�F�� �\�|��9����w��B��kS2��X[�{ae����ʅ�J���JE��1x>�*C�N`�	��.l�v��L�2�l_�����Ե��Muаl/+��3�6�9<���[�]٭s �'4I�}AS+Lm�X�>N�J��$+�Kn�Ԏ���߂���m���0B�?�=��ٔix2|������xT������}�yᢝ(9l����28�V���li����y0��]�>9��gQ�+�D�({K7)��t�kJ#"��v���t�s#j��[�X�`i��C��lY���q�ݡ8]�j�]aܦ��j$g0��A�<�Ν���ޞ V+���.:�(����r�t^�U�՛jx���Cs�'��7��Y�������9��7�V9��prJ�Z�nϐb�u����>3�8�����øqm�A��D�u}�����:'3��/#!�i[��]� 76p?)�Hjz�a3o�N����]���ժ��}����G�\�I~'7�c	 �fo��=@����?sMq�؇)1;Sso���vV������Yk}*z�Q�l;]���w��JAT�۩����;����-
 5�,m��ΰV��м,�&�%��H�7�\\�l]	M�]�++�'wj"�a
�Vp;�a��P4CAX\`�1��!�h�cAG�G��!hF�M��N��!�.�lQ@dFmg��E5�a�).v�W���D�:p7�S�9���w9�I.���g�Y2�jh��WaK��Q�n�£��U�}	�.�5Ւ.����Y�g��
��g�r�8���C��P�%����[�������S\�4���_(|�.����/[�x*6�a^�'�u4����^��ȭ
Үg���la�b(���g�|��x�y���/��`�'+�p�1a��w�?����K=W�G�JU����h�D�40��[5��[�Z8���
 �|'��`����j���P�2�XC~1�>�o~�[>�&m�a��=`�$"��O%+/����R�<���KY�7��Z@�Ӄjҹ`��,j���oF�ķ_e���AYB����&F�H�Pv6��@�Y�on��R㋴�bZ�8wpm���D�cj�9!�����ڝ:���t�� ��n.Zsh[$�R_H��,-���ut>����t��n�%ɝ���W��e_������^�,ݭNu)�t�����ݲ�%q0?����|��TO{���m/z+AU4�x�z;�t(O�9I7܇�F�q��<tLkD���Y&�U��J�q��1�T�vG��-�:���?G+H��3_��y4:�^���z�Gk1'0D���Kaww�!�"7�o<��O��>�~"t� ӣ ,d>�4���P 1�O�,Ga�/�!���P�*ik辶�N֑�3��_"���ذ��Yr��cQ9���x�� # ����T�&��d[s�H�at �Q0���+(Ip�[�=�7&�^Z�� �g��W������B7]���b?��&c#@�/�w�����]%zZ]Y=29�c������oL'�G��ٕ��j�!��6��/��O9�a%k��6����r���V���k0�]��%Dh9��(�$[���������~����-2�Gjn�q߃3#3?�P펞J��$ ���4y���+\�#���I���q�InDHyW8~���魉��1'���/�x�7�`�l˯=��5��wvg���D�ؔ�� ^���dЊ~}%���c�=HѦ��~�F��8�X���0��s-Ƽ*�$˶둴��~���Zj��� |�"�J���85�v����H�N5Py�4��K�n�n�H�����'=x�w�6Qwd;,u�.���܂:��<U8�.?
����
[1|MOP>�D^�/��v{x� ���_�E�袠&C�<43�D�d= :#�1^ۉ�"�AO�J.��+-^��G.�2�Tl\��Y�cu���fG�d�>*�Т��z�Y�!Ղ��(!��(���[��|���g�\+����4LRM�EӬ>ůdN�#�8��d�wz�G5�Lg+����FO�s��/��@�-'�����6�t[��:���NpZ����&s��B��:Y���bc|�����^���k_�}��	��02�p�	����$��lt���'9X��Y(-��� <5EC�47���\�qL�,η��?Bd�BΈf��1%���p%��}0����i��l��W~���${���/�?U��qM^�\� ����J��C_�p��ǭ�%��1I^sa|���x\Ҵ纻��KBa"��y}Y,�w��5E�ד����rT�S�SWW/��x�ˋ4ʲ�:�f��)����MxwC�LbX�O�~$�8����A�Ȼ-���:� \;��w�����6�ſUY�M�t7^6T�?�𶒔lWy�7��;��ӆ�z�����I� n������?�{�0詫y������s���;�14^TW]���
k3��@I�s�sz��d�z���qw{K�F[(>���Fri� ��V��;n{㿔��بX b�� Ry�ȉ��2ΆKi�#�o���B#*�ٻ�Ӕ��"���p<'�b+�4C�ٺ{�w�������k	j��� <Om;���tK
��q����BNz�i� 䍾
	͝�(�9j����@i��۴ZD�b.22k�.2�>s_�3zk��ua.����	z��$�*�7�/�{��A����bO���n[�H�^�xldE���{w;>�o��0>f�]�4bݫè�V�;�ţ$��h��]��
ǹs���tj��/ޛ��_�Ln���X�*�g��*��;n��b��B��1�*�CaFl�c�i�5�����*3���N2��5�X�W���_��.�S+9a� =J-����K��dh\�R՞@�� ~a@�$j�S���#�ت��?q�?��X�?��𯰹�=�ŏK6c���.~��j�����^)����@F�.���JR�Yr�A�^fʽ����(5ˉ��9��ҷP���8���+h%)M��� lx�E��˖f?�ې�Џ���J5����B�9�kÒ�vS �8@��&��L{���S#y�\1�u�c��
2=���U�����2��s�R������{z���R&m;+ ^9����.�	�k����PL�פW˳�A��)��D0fiY]��+s�۰$�ɯ�\[n�nDT�a��)F����е���� [7ü8E�lR%!'v`Bf`F�{eAF��.����0��x�49u,OEn�L1�̕���}2U&��S��� ����8��1�B�'��J�b���,���!aU���o�Ye�%,����⯈�t���4�-��?���U��?gf�T-�F��O�F��sՄ>���Y|d�;��Z�LI?���\p�T�4��\���7��HAx����Sc"#�s	�
�\�޲]�o�����0��ˣ"�ĂS?X?�.y�y��(�^
s�!��;�̮��^�C�ؓ����z=�9׈�5�ۯ)����[\̀����ب5^�XQmgƾ�ʜ�K�7����{u7��#\���,c�H�Wk)\[,�y D�Z��G%r�X[�f�0�,H�vƝ��j��Xc%he4�6��ԹmA��:@L��K47g�A�7^�}뽓�FR��GcU��y�᧛
B�oЏ����+��nU�6~qlw�u��/k�u�ɴ�ʣ�^��.�b��/�]6Ibm�kW�qدso$$j�Tu�	�4u�l�4Ɉ��%�Z��XW&��F�B�`ܺ$ROՔ�z���It%�hd!}9H[���A�pIE�FxœZdC���ak<�7�_
��ҁ=�����^�{e^���|�z�=��o�a��z.��L} �9�w��}��n{�����0�T'N�#oɽ��GE�{��"c[���+��w��.�w�#r����R�����3k8@�@E��x��ԕ��LG�'P�<�&����Lt>��W��*B=�x2>�v�#?�$,�i�t����2P���MC�UԼ���X���?`|ӂ���8��
���1�~o�$���O�a�����-�߀�q�_Z�Ԇqɾo�}���
�Cy�B{��L-;fTUk�vJӅ	^T�k�h��J��7Ӈ����^�2�����~A�]���, �rx(rN�Q���U�@4'�wX��r��c�����/�\�J,yߖ0f���w'�/����A���m�U��D�������AU/RZ�b9�ʓ?{6c�7�B�`��G��R���唆^���\�`�Ra�=d#O*�@q\I��YX|�M�~�Q�mlRy�D7��S7����ml\wF�|�[�)B۲����K�Y��Υ'
���o���?�%`��:-��37Xt���E�̖��\�B(��b�~�ēE&8�w����ӱ����\�N����G
�:�_�ܯ�}�e&Fg�<�;=p�\ƊI���Q���d�9���S�&w�h�岨J��z���l_�#���evdn�~��ѤX��m����}�.+d0������T�f=��ۘ����-�Q�J��㚈�U�˂/&�7sԡ�{��	;rZ�e�^���n`�:��.����C��, �!��W|u��K�~$���.���(�T�b���ڻ?SR�	J%tkLB�V��8�N��ߌu�Xs�$M�G�h��i�ϩ�i�q�/8�����g�X0���g���f5r��?iEK�+U�>��U#ףƲ��I����t���j�f���WrR�j��q9H��+�Xvw�\����*M0 WZ2�l����b�S������_��8�-f�~��l-�"�#�$;u-�f����8�	k#ʊ��-�g����h3�������YqԘ���V�ߑLV=�pk�$��E`��Ĥ�O���r"��?IU���
���̆x8�&���3���H.Ұ��ۯmz�y��D����*|ӓ���$���b�Q3�!�$J.	p{@h|~; l-n�8e�y�\^�F~uq,�P,�@r��W���`��p`��DȄfc�T6ZVS���36����C�i��R=�ָ/�O��P�����|�7Б �ƄB��o����o��]7�4iՑZ#1�"u���	xk�*�Z�yy�i�� v	��V/���Ƅ\�;��ףMc�ʨ<;�"v�՘����G�0�k&�8��zT����E�c�_q��y�Ɇ=!�ۤ1��"��Wc�ʚ܏�eS9�����9��Q�Io��fv�{�$7K�sLY�.������DZZ�Y*�Q����źM��GX���j�C$ba�l=�aZ�W7�H�{�������Q������{w��s,rԭ7�Pg�(��y��$����.������9n�	�|Yc�<H�򉹨
א��
%mi��`I�z�6�P�!�`gI	GvA�܅���5C�Sӻ&9�j7��3���/#kw!����-4��s&�����SY�������_a�s70i��Y|<�h��u��D�fOZV�7A�B�����/.�P�ڼ
�9��d�3��s�gӫoMU��#�Dq۷uĥ�[Rm�l���9M��A�Л���f:�.�z��#V4�Ƥ��gİ�e��"ux��Q�<���4����e*�	��.0�b�R$H��Ơ�cSx�G񦌼a��Z�6Yn����3{;�u�g�	������Zpw���T<�g��7�3���_Ư�<��W�ak+�CQ��b�X�N]+��xx��2i����\�lh��M��.�̭���-����߭~Y�)F�� yo�eq;t>�e��M��UN�w���ӗ[�}w�H�H:��VLYޓ��w��¹��34�֔s)@���dT���Ɣ�z�QMVtN�*���
����[�(w^�s�^-�{_�lߵ�Y>m��T����b'#�F���t�W���v���
Q�����S��kq�%����zxB"1d��������<d�*tcw���}�����-\��J,:�"Iҁ8�´A�aBV_�P4�?'�57������ꑢ�\ۘ����RSa�Ƙv}rl�S����H.=�S�kV����*�����vx�	zNBN~��/SR��6��0~�Lh u�(к��=T��	)��O������%��m{�O.�K�'��V�d$,����aX���	�ٷ��^%	�;�
>&�K�+&L 
�C���T��i 5���+�\\���"⩐��֧�]��,�}�haB�>��;���E1�Z��j�?�-S�"�fe��|%#)>�H����~%��� ��"Z_�
ɠ�ػKa��g��=-�-h���LYh��%�J�Tb�.'h�"�ʧ�P%ͤ�r���n'�����gF!�:��P�U�֞C�5�G�gZ�I-��DI�pV�&ɕ{3��u��]���B��2&nm�ԙɠ;Ni]4�i+�2"!�D7��JQ�y&��Q�UƄC!*[b_UE�o8HC�C�5�zQ֖ܒ�T���� L̮ʽ �t�u�I��L{ie֯x.u5��>���#j����)~3z?�O� ��cX�ԛ�?�  �7�h���^��R��-q�¤��aQ��bA�O�Wt�����v������Y���v���vq��/r
�!f>z�7i�FYk�o8��g���:}�@/�9ј���gG.Ȟ��d��!k+6�Q��t��,Q�.&�� ��&��S�P��8�Y�����1���N$�څ5�@O;;u�>�r������7_�ݥ��L��?��-�kz[T�9Z�wv���W���B�����jV4��_��R芷Q\<u���*"���f]�[E�����<B��(�׶'��;�g�fEN׿e�lڧ���E��A�ޥ��p��T���d�5��A��^N����˲����el����/BG��4� �`\�Af�.Ķ���`NR@�æZ\���Z�R�HL�Y$
$}5pI�5ɏ��@� H��D}*#6��)!n���K6!xތ[�ϱ�̡�5��@o���X�!'��s �/�H�Ff�����Ϊw��B
�:ҏQ��(	u�6X�h���\!��3j!b�wQ�	} 
�I�e3i.��Uw>�����M��6�Y֚,����
�����g�z�������n�7�����/{!����N�%�~ױ�
S���V4u������5�
�2��\h 0���d�z��R=�����%!5�gԭ��U�U?S��&��1�|D&��w��α@�rVi��e�M��P/ʂ	��v����� ��~D�����Eux��?��?����7{�O,e�Wm������?o���aB�0��u�A�p�5=���P"sk\\Mgw��g}P���D�Q��D���B �&P�.�������ۃ	��QaQ2>a@�W|�vl�e8'�/�L�ai�{W|���	]��H�V��DBۗU��d�|��&����l9Wk����O(]4�����`ѓ�$�4��������bh��Ae�y�\Ľ2�N�+h�)EZ�JV���pE�|�j�U�12��}��؞u
$H�SY���)סxJ����fH�AX>�ߏ���=�P{"��$���.�O9���Of���	<u��>� ?oѐ��j�	ȃ�'�K`O5��w�u{�g*��a}�����?��*��U�`��Jl���ί��� �G`Zt�����]�{Zy �W`/Πp�	���]{'�D���K�e1fyQ3���	��9x)/Ӵԥ�S
�]�|�f��ݖ��;b���)��>�3�H{�M��'���C�"����S�S�sHG��{�걌��:憒5M�s�˵�Z�}TB�M�HB�F����g�DL��ew�ӽ�˳��!����t�ь�8N���eS�]��y�x8<���`�?l�N������;�D�x�6��4�p�=��.B�s��W�ª�X����y�h"�
�U/��Y7O�TJ_7�i� "Cc�x�l��n ��~�T I��Ձ<�P&LE�!%���9�J������s�����=aTb1<��z�tz��^LT�aػ���:�]�.��g�Ŷʽ���}���-�ө_�V��eu�!1�Y�q���g7GմL�	�^�E����=��)�-ͺB%YʋbT}hD����&{s�CX�u�#�Խ�Am�����z��I�Zi�%n�G��^γi~f7�/�B{O;g�|7��Q�\�N�9?`����D��w�2e�& �w���zڷ�X�f(�S�P����'\���H�A��D�U� w]��ے�9��N�*w��SE��e���A��N�Zt9[־��Q�����¬�٭\��7�m�(P����ȏ˃aB�ZFId�$�7R)	A�"<D�<k(��s���E65,c�������ݛ���VqU�7���5wcA�Kn�ؼx����v��s��/�1�%���w��na4����p�6	���Fǻ����~[Ku�3aO������x������y@���D�M1$������.�Ņ\�U�I��M�c��c�2�Z1��������AI���K
�E��<+yu�k�t���C<D�=.G��H&R��IOQ[�ڻ��k2P��%��P�m5G����<˕�?i�>�P3�w�,A�I3�YK���&o4(� �	�_�
�pyE���Y ����A���%Ԫ���6��@�5c�-��I/�K��I�e��NvsW�E��a
sO���|up9�m*��Rk�P�h�Uul�ڗ��fY�A��j>����=
t�s�O�D-r����R�'3�{&��.)�����U纃�v�5t'���ݽT�;-Td�5gq�@Z�t�ߗ�x�@O��DB>�d-�%=2$4����#P#���R*�'WXV�!�%:��J P��ʂ@�|^M&�A}�P��2|�,epF5��)Z�f{#�N@&����{E�c4��G��w �T�����/q���MQ]�6���@3U
��7��|P��N�&LO��������%����Ɠ���g��\+�it�O(���Ne7̇#mZꆐ�na�z��z���<z|:_���MT}^RUY����5Y�S�m���~?o)j,.y	���,�K�a������|��y�w��B������)A���<� �:�����9�m�V�oJ��IB���׮���ƭ�h�����r��+�R�3x�� fb����X��_x<&��p��߫�7b5S�Zx�(�\<M���]")��\�^'�K�t�
�>d'��[���<1ۍ�
_��՟i򰌬wA�#b���[���6n?_�J��J���?]��m,���/d�i0\�Ʊ]{{�B��@
�~D��/����LHl_Q�)��eg!f��`>�+��َ�"4�n򧈴���7k��Ϟ��Țs��Բ�ΡK'ܰ�����K����w��+K<��A�ow�7��; +�Ģ�@��/�F�ՂB�l��w{h�,F���"�u8G�l�j�f�c����Y3��FAA����@�sG�Ѡk�Ug�"�3����94ֽW@��7c�e�Ù��Ό�y�i�����~��[UH��2�u��aϡ�h>���i�<Wl2�,~�o��+��U��*�ݟ�>��z6����t�]�����cs3�j�A������a��F��9i�p��k���{1v�0�W�L�\�<���_��=�'F&��u���I��yW*;�C^:�ULʬRJ�k!@ߖ��Dy���]�<2���[��EG���K�D��x��w��n?���A�����3�������&���A�^C�5Aw��$�`�b~O�	���J�k���ά�q�¢������`%'��RK�=X�����4����w��,�h�P�s�V�W"�!�)�������)�����`zͶ�g(v��6
28�'h���N���95�L�x�M�Ʀ��o���'��7��f�@�O��.����Ȃ~���W��^'���B~����V�%߷�[�Y+���2��T�$�]�>���u|�1{��I�<�)�ؑ�&5腱����0�7ʄ{���au.g�����ܲ���F�+���p�D���毱���c����K����&eHh�5��aS����%��5xΤ���ҧD�����9�?�L�uh�U�1P��idzu&�P8k%�Bi��i$�"K�l����!�6�ᵣ�ŃZ�M���A�=�|m��ӷ]�.w�7�*/=�-/�OC�@*ᅞ-ױ���:%V�h�ތJ����u��oZ�+��x�a�z�2��S
�ǽPX!y�Ъ�9Fd���l�͟��. o߮�0 k�_L\�Rؒ%=���$eD�(=����w�+$��֩�a����(dc�Hm��5������&��i�;`��2� ��������i�xW:rdZ�{*6�^k���o9��Ex���(�&YĉǮ��\	V˓$܈�'�g�rvv
���h���\Qe�l�,�t
{�(�*:�"�$,�n@V�UŤ��`��;��0���G��]�3��/+�<Q{�
"l<�[�;���"�>���Ta��l!U��Un,1{l��h���_Y��d��O����$��p�]������G�W�!���v�3���O�"�
����B5?§-��c9y��O�k��� ��M�p<�-����Zh9���[����y%q뜎����������iqw�ʌ~E��ڛ�y��uI���"���n�@�û��O$��9C��<Q`��F��!t~X�M�m`_׈�5o�X|Gp#�=�*��{��tJV�����)�W|Ȥ4���ǟ��+�g��:�kX$a��{ښ:d;/��ɧZyoF�H��hc�4�O'���[K���it�I�Ň?�e�����BX;u���B?��<���u��G�:�# ���h��n��D�g�{\��ً7�<>�)�ϗ�3O��S�0l�\�
�e�+�/�g�9ޱe���(_���j�D��rd����Df'tR�4[��K�|JV�f��d�3��%���L��_���Y���ߐ�J��M�fM�Gu8�S��-��+6�j׷�Q�D�5D���(��$ s�CO'�/��R������W���u��P�_��SQp�F�M��"�nA#��,2Ql&R-�|���e�r ���ê,U�4�_	��O�'f�T��𓃤�E����I�(=V)��+�<�=
���������$E�Ϧe�X�=J��}Tǫ�#��D��T:��^ַ�	Y#h�G���csDm��P��;������5�H���6�L��p�j�ڪ���L&{Z{�Rs��Pa��r۫}�#nJO	!7Ӣ����n�`T�+���mT��@~o��O~�԰���5�U�b���j���~�ys&���*���s�qd[
�Ƶ4�z�� z	�H�U��m�Wa��v���/��i�9u���V5�U�2��0�Ělj���T�@��#B.�j4��(��������!{��GF.Ɖ��#�&���#1L�CF�4�-M*��I��1L�m�E��R�����M�$~��x�/�f��+#��01�us�mtx�8����t�9���n��O�2��)��&,�_��>j��^�,v�;he��Y��4ͪ8�^���)��g�i�|i����^�#'JA�t����s�W~H?5��9��}`mvv�*�r��W�e�wD���?��ȓb����zI�Kh�Y�J�:&�$�p����̤˙Wmi��⼥Vs8���Oc��	uaJmR�\��A틘�y}Qk���M��qo�X@\���ƍ�6����ns'̫g�|�dK=�&zr�(�ڂ�n.�k���AM�~�*U�v}M����w�~y2x��J�����M]�C�y9�JH���{�Ά��U�U˒����e���a��U��~�@������i:�
�<��>��B�i�,eyQ��p<"�&Q���;��{�i��*�y�����sg����|q؄�)�s��<��G�\��,�\�e�7�u�g`�rJУB
�i�n0��b�Gy�T.�6�Z��n��ΗKn!���t�?s�L0--��oa]^)��clZQc�״6��ɺ ��Be<W:@�����,�m�/�+ӥ_8�O}o�9$XJ�b�Y���֐�L^p��qn���X��{x籉��,�=)2���e��8��
}�]��G�W�zI��i�d"�ID�=�Pt��l؜IZ(�(��ћ�j�'X�I�PgW�J��)/�ZH~���r��Y+ �R���_�DX�
6E0����SҘ�K-f��tYφ�g��oN}IF8Hx?x��_������g@�����x��|"���I����Au-P��L+��H�?��Ȝ�RM���o�(�0��1��T]�q�'	���y��F��q�wnY���4)��,�5�:]2��:Y��{Xr�?sB\�Ff�}�8��uI�A��J��}#C�S��1��J[���C��W��k�{���9�@8�zԝ�U5�7k����'i�ݼ'�/��B3�l��?B��j����\�?es�c-C51���Jq�`������?z�洮"��K�#�)	�������6�LM����l�bgF|iرF��ۿj!{,��(�0�~2|�+�-���0}��
:fC��<|?&��4�2��Y�͚L��S9���Ȍ���:��55���S���3��H.WJM�2���S�u�
�{(Fw?΢_�c��R}�U��%��nQI�%"����v�q7$�&]L��'*��of�_+���ѧ執&H�23!@��c� L\�)����E_٧,�GLn���l$|�*/��h�6l^� �nD��Fc0�6���z��3n`r�i-�s�۞p�v&u��c��m2��NԋƬᵜ��mo�������^վ(�y��:z�T#+9���ʇ���F�to}�Rhm� 5��p&yk�H�-���L�1f��2'߬����.��Dk�\�}��)�[��v��1���.��+e٧�2?�&g��s O}3�sS�N�0�3)�?>N����[`$(�OK2�&<�R���������Mt_Mw�SH�̰�A���r�h������?�6'�ZvV;����rDr&�z)�t�ƌ���#�W�X;9����n��z2F(q��n��M}(ß˫3�g��m�i<��Z<�&�� "a���7�Cf��3c��A��^��]z���U��B���q�6m��:@3P/D�\\mZ��(9�;�:Z}O�O�B�+����]N�(l���w
ފ�?�>��R�f~�H�M�̑p=4�Ba7�}F|>��:�6�w�i9��Q��<͔`��m޴+h���9����%��T����5|F���_�7�f� �D�K"�(.ඇNt*5�̰ΈxmM*�9��o�O�VԢ��b%D���6m^���M�Էp4�e�H���z�aN�,�Q��y�K�$�(�~��e��ם#E���3܇������-VP�D�u����!���T�b�ٖ�u!����N����ݧ�����['��ҹ`QϑnPUK坸����T�U)p ]�pE�����u�D�,�mb�
;jE��;X��-������[�5�a��y�b�����ޢ��O�]�@sni�����Y�CJ;��ѡY��XJҁ��
��UF��S�u@L�+�/��[m&��1�X�A<b��5\���������l\�_�GW9��/�c�'6���X�=�a>��*ef	0��0���e{��I�y?k~�e������ց��,�fҙr3N��ʽ�e6��yD�l��0T"$��2NK��W"(��H��O���:n�j<:H"�C7�S��ԭ�,�F׶�pN]�_fx��)F�yUj���!Q��G�m"��Fܜ�'9x�ӈ�x�߫�X���%� ��7=�skJd�1,�1���os(�3�D��C<�#bE��}fѤ�Ǌ�;L4���D-�_|���6���<��Or��� ��`:PX |��1����K��q��HQ�k���j����f~��]3�8�3��Σ����,��ޯ�U7t�ئ)��3$�څ`׭d�`�Ci�-pD�����!�\�� $�Y�w���l����*���)�J��y*�>�{l�þg�K�x�m��u@��l��h]� ��j)��ۘ�ӈ����B}��.80�C�R�4��e�M��Ӝ�,�XHLL&��Ë��jVӖ���O-��0%�޹'�d�њ�^<�"_
a�fr.�$�f.e���p�%#���EP4$zCj�Ox��R�l�O��	��.�P��4��
'�����o��4��Y 5����5E#�_����z�� �7S,8�5ky��Q���K�:*u�OZ� �A�vQ�0���^�l��2x��m �5yP�-���"$� �T���V�_��̿��z��N�1����}�?nU�$b�A������s�O�f�f��ɀǏ�j8���t��F��q8�&$���ղ݂X����<ۤ �����U�p�E���=�z� �Ў/#9�֕�#E�32��q��*�Ȁ"ի��^��LCsX����M�{�p�i�)&=|#4q������:-�Bqe<&�`�	
������D��ރ�+Q/��&�q\6�l�,��Jr?��"����PO���A�<<���7 m��2g'��/oWk���m�<g"��.6�ݩ�R{�1��݆j�dF�:4"B})�A�x�� sfS,�]LnT�ϰY����.xO��-ޯr�0ə���@ʮ������.Į���7��<��}�j1��?���
/��� F�9�쳋�ԁC:��4y�hZ����h%]/.X�~�4��z�6����s�y76]�� ]t��f:_��(ŊK
8��}�������������0�w�-u?��m%TUǫ|����1Ɣ�d�V�$A�{��1�>r8�'�6�Ќ���l��CqϨc�WAWx�7�d�r�Ƞ=H�Wݜj��2�ɵ�U��
xNkA��, ��%ľ*4O�.E��H�Io%ݓX܅G
��E�7l��f~��OE[�>�X�>=�VoVo��-a��5#� -5&���ǎu�85+Au�E=��8���\��D]�9�q6'�`O��h��6T���=����6�\G����+b�\p��t�0�"zn3X���Ou`	��A��k/��5�~�?��yAa�'�mg��G{@�DlA�H��P��G.��{�q@3��)@cU~ݠ�c�R`�kX�w	�p8�#������[��r��UXy6���@�i>&��W�~��A�`OQ]����P�aO�������ۆ�,H���]���e��0e%F����l�X��/�<F�ܼ'|*í:PF��#Q�*r����1�=�]��q7щ������>��#��D�V������ܩ���f	J���j�p�r�U���߭���ȞK��I������(�@��>$��۱�c�Q�(���W`I��5j��32 �K��un8{V��jK�[NA��]4�M=�s3�����cH5������!p�;9�W�H��j熽�o<&���]�JrC����ϊ��������mx�Q�9�ӫo�t�"��4�}����K؏��X�3�b�^+���Q��9��S�\�� �3�[��eqF K�D��QĹ+��>Hs�M���6<גؚ5v�#���%A�qsЁ��Z�ň��|[nݽ��!�#���ڿeV'���8�4�*�� �yJ�2U
�v
NMzň%m��Alb��"��5��d���<pP�h�T�K_L��W$Rt�tAւX<x]�����?��� �Rm`���ν1h�ԕ����������Aԓ�C,����?�2��EX�KYi+�J�K&�2����@M�>��	E�=�;G��f�WX`J����'�Qg��%��y�A�[�瓄D!����-�c,
��*<z�����ڗ_�i�߅�]��KT�j�:�"PB���n;���T���d����X&� �� DmL\��<�% ���e�S��h/J:�1T|�.�m�P� =2�C�0�ŭxh�A����h�t���cw �1# �ҏ`�j��q���b|;LK.���W,���z:�����j%8�*�6��U�� �ʸ�(��+s�yJȑ�YӮId�/�3��	^ߢ�N�����%	e?p������َ޵v�zx$Yr\X?��_a!�0R	_����_��ꕮ����HE�I�a�3��S�>u�֗j�`��*`�ݧ#=��)�Nܗ	^o�r�*Q*�pԐn���0��S�e~&�v�;��������S.o�<�����������̤[;����7�6��	�[����@aN7���̢Q��f�W;<l̽𓫾b�2��h�(�j�W�IM��ѳ���V���B��XN����$���4H#]�X���=�l#E�<�%���)$����G�v�$��^�Ę1R�=	��b�����f�<��B����Y1E�^�6m��q�����+NQ8FQ�y���X���T���(lKB�4LA��'��6�K(/���(���$[!i��(7���Թ���lF��)˱�O��Q����fل�i|����Ҩ�S�����]�|ݫ���2��3G�ӑO��Iw�0�Vh�q�>�&CX��
1K��aYĆ�����G:֟�Vշ�#�4���Ok��S|�����f��o�_����A\��F��f�[⏫DK9'��ƅ��wdR���>�M�ܮ��^�����p�J}�����X�OX�Oㇻ-ٚV����$uU+2��w�����I�XZbk��n��z�bD��ۨ����e�?�� ��7��nӱ�e�\��8feC"�g��Vk$�v�(w���)��|�� ԫ5]-k�~���5g�$����ƅ�F�F:9�Y����wvK�	/��! �T���կT�D�L ��Q�x!��%��^�k�!Q�	P # aH=��_��	�Q�Iv��4p�����5�͎0S���F̴f���=�I^�N�N�rk6�@F�׺61,�8)9.������r�$�_�↪�����3	\�
Gc~(!�rE��$���w�>!��N��
���}�w�)��&g﹅%W��ò҅��YW
���I�J�2�ToE�- ����`<ܿ�vPI_���� ��<�\�E�3��4_5�\X`Y���d��2d�Q��V<C[So��P��嵑{%����<Z��.��i�K��p�΄΋��l�/��@�f3���rSwu��ު�f��zQt��VH& �*n��M�c)������ �����%���9��a���\;�'Y)�U9��{5QeN�Ot�/����+��J�
��߰^�����ز���ձ�)p.F�0:c&I���l��bC�5A���LV� Q�l٥q;����F��B�a<�,��.M��C����͌�\�Z���E>I���F��$�D���{���a�Hځ?����$u���嗧�w0�G9f<���n~��'Ɗ�d�f�@�a�ߕ��VyeQA	��d9j�9�[0��XGo���I�{�g�4�\0 ��^�EfK�����9h�曓y�x���Or���9q��r��4����CiDox��#��-�":�uYg��Fh���#1,�Y�8��\D���)��������qM�^�mO����Xf���|	�����;	f�W�݆;Ⱦ  ���\��% SwH;)ɋ�gqg�|k�D�DB�!���#��IڼL�$��i@@v�әa�������;$�f�x�>�j�1��T�ς(��*����dP��̼
�?4��5���V�f�M��A���A�X���uU���^�����L��1���ʀ�λ��IL��m]�<1bO8ɫ/�*�2J"����o'�$��D�}"ܒ"��YQ�2&��'�J1�?�9o��6X�� �/f<M��ԭXI�L�U�����������M��p8�B��d�bF6.����`��_���Z	����h����!L�7�F�"2���ο��g���Z� L��K�R��nAl�*��}�u��J>C�_$< ��%�;���E�f2�^T����\�`L�n�1���u�.�3��-�f	�Jo�p}���%n.Xn�n�Kk)Y@b�ѹ^0%�r�+UX�;zng��$h��ޠaO��[��CW�tTy���y������-�#q,�*���V�(����Q��K<l���	Ga�HWM�tԣ[K��pR�|�bgA��41��,W��Z�'��gDp��C+=�B$�l�WYGň��MSց�[<���a$t��o��r�}�EA�� |��6A�RJ':�,��Q�k �H5ƿ�݅��]1zf;^D�"Sf�\�Ֆ�tEJ�uqO�W4=���. !�e��Fd)���7}T�$������q&����Dϵ�O{�!�DV����6o�F��]V�~��ô=׳�?��+ާ��s�kg_k��:�g��={��Η���J.��^{�*��%��BvT3�w��~��K��"�V�ҵ�IJ�GE�������>�|��L���X�E�E�z�h��沃[4vf#�m#)�L�䏈h�=����f��:��D���0O ��YZ�q�T�)��fVx	�FQ�^�mQh9X�^�u��>��=)���d8�rV����]IG��sr�����â�pt���]��B�a�P�'bfF��O�p�~�Jo��;�+�`�	I�ڞM(l�=!&N(��D��-b�WR��ţ��;r���)�e��I��z/�[����xC9�p��c�h]l��A[���.���
����D�����Yxp]��n�<.���o� �n�l�N�#'b�e��'@���P��f��.Ӊ�Fshn)�����a�'�s����YWĻ�p]w�@Le��Ua1J�k/y�3���F���B��y�_��+��n5�����RWqm�ԆxT����}k^���7\��Ѭ)������Zk{,l��0�8Ð\��<�V�<����#������^��.��]�nkS.���m�*b_�m(��LA���6�RpN�]g�,)�m��*(�,,�U�Vd@0��m�w�Hg8F�K[��6��I&/��j|v�m��@�+�M�p�8����"g~	1�S�X��H'���]�%�EL�i�WO��M�a/v�S���VN`����unA�?� {:�x.�������)a~���5%<)�h�:Y*��!mO�����CF�8~]h������y8�ve�	{u�h��C�v��g/i\��
�+�hI��)���,��Խ�3���2ͮV|�͑º��W�c�@�^ú�G4h��#Rt44"����1-�k��0�.[ Z9�/�e L����	���K�ˆ���NE�/�9$�%���M4�hV�q��W�fө}uE����*C0��ӲN���A1h�f]"���Z��l����t>��|Bes*"v���s�hP*�(K|��p���2���W�}0�'0�B.�~/V�jp���O�ߊ/��Zz��|���&L(r5�1Ӄ�hSX�<�wފJ���I�ߜ���N~w���xv�lO�vR%A�=R����C͟����E��U🔩ϧ�����z1�T���:.�Ѿw�Rl�����dڮ������HaT�2Ӽ$�6�0ӂ�.������&��{�2A�_�&�s�s�<�a(+ė Y�1�o�d�i�]� ���q�%�	D{-���ܫ�si�挱 ��D��]�p4��ӸW殭��75,�X���g��e�Izt<�����#�X�S}����A7�H�ϸ<��«M�G�z*��ya����|�bܐc�j�2��
 �е��fc�)�Ѣ�"c!v8�������3��X@�V�Ͷ���=l[Zw��c��u����"Z����l$K	�k�"���=��]�����p���}Gb�(7x$0g��9H	S�EԱ��6�h�E�s����=<��q��6����~��2?%ώYjVt�
Sz�)��[�.IV��Ղ.�/(*ٙ�D�G:t��pN��`�ȅ#B��3vE 'Ͷ-~��� ���&e�*:����Q�`��g8fU\"����5cP�:5�Mf	��<ѡ��:|':���Y���L���jr�Q9z�eW�V�D��X��D	x톥��!����<ˁuV�4I�P���Υ��ŝ�Ph��vL�qwn�����b_R�ҙ���" D��x�éX]#\�� ���k�i{������)q��O����������m�0�ϡ��4����0<yh���j��
��=��
I^�C��_�Ui�5�Q�� ��-ơ��W�(E*p�.�6Œ
������z��w*�����j��{�غ�|Ow��E`3��|��^���0�߇�uWQ�Ŗ˱F������a��Ό#l_���b��5<*<E�O;@�qx�>�:���^>��b��h(P|ƚ���"����@W�!V��|!I;��뫥	8C�"���5��J���t'�9�ݸ�xd��JF��~�f��5�v)`K��1�%͓,H�j��ck�@�PY�rJA}��%#�Yr����A���D��$����F ��`��D7����^���G
}н�{'��z��8�CC�yx�Lk�Z�2�J\h���i@��(Ѽċ��]�̠�Z2Z.�xW+QA�a��3�˱|ԑ|�W�H����{=��:rnޔ�=#��t��z�L��#���'���Xs�[	'C$�%�AY�$�F��Q�K~Z&�{T�_�9�W����o$ì������I�P�!\T>���Z9�V�&����3�9j�z�H���l@6�@�Y\�$�,[���$]�\%��4��}�!�X/�.�E��rG�*p$q)IOI�!���TN7]��E�IU>[j�H��3N�!�@-��_];�6
���VW�� ��Y����Cu<���6��O��4�Ge2MF�'A�?߆���_<��dA�1���^��xݴ��s��܁��k�{��!y�a�<e�o�f,��c�(	}3{ ��hf����� !����B�p/��R�=��d�J�ퟖMc�����,������F�R�ҵ�%������F[4#,6��&#����O��,1�uJ��*�|6^jL��Rl�긃���$�B4�-���;��|�$'U��8Ԉ=9z=+�*Y��,�P�k����N�Y�J�Gh�a2���m�s�����.�#��7�Μ��M��I8~��cߠ��V�
,Px�M ����|O���q�$T��O�(��ߑ�H��n��[�!c�sƝ���9�-CP!�a�}��s}�-��NxP�����ê�I:�f7}M��jW�E�C#�ANw�k0T�,%	���
��=̹n��	G��2V#��Q�H���;�/y��
������Ո��8.�I
Mb�31#�2���'��ɞ�8�W�4�[� �y��%�z�}�3y�;��˫ĚIc��z���j��8|��*�Q��23v$wk<�N�)�		�{�)��Z���
m� rc �⎮"��L�~���N��Ļ|����'�衙����m)��ɂ�5�WZ0�+��q��J �On��%0HTU���~���r�w92��5g�FVPB(۝A��>���D J��sF^�w�u���}ILA9s��f�(���߿g���sN�>f�c��n�֗�؝�`q8����d�z��0����>�[���P�\�<�}�↗�^�ܞ�2��@0��g�Jov{�l��B�|=2H�W���c������mSՈ?ȄZo��X���i�����9:����d��!��x�&�=/[���nm�h."�Kj8���r�	S�Y���LGM7#��>k/D"{z��G�m{��ӹ]������GIp��3�JM����K�.HK̏��r�S���{�W� �g.���L��� c�x�7�[kQGr��P���eP��^�w��X4�9\O��-���h����W($�E��DN��%�D���mΐ���&%]��*M� Ry�dOY�}Xs=�RQl�3w��0��xlw�u�Y��U���FUD��j��b��uX�����]tq��溘��C�����k�9L��Z�����cY�F����������e�/��j�*Շ��������l�J��	=���	CJZuL���a�0���&w��e����?T3n�]��QqE�19W���rJ�U���(҃�S�<뢮�j��.o'�"I�1��g�i�VY����L�Fz;����2������i��?�i����Q�
��8�j`�L�k��1��ml�ъ��'\K�f{w�����O.;h��"�W9��:{�P�d�Yd��u����>��Kz[mt#w/U�*O��Bi��H@G�������k���2JЋ=��V6��4��ڑ`kz��:�����V�o��	�=E��C!�(r+�~MU=R�+��Dp0�D!�[��2��j�;�\�`�m��|Ϧ�3��d��Zd�S������n8���@#���	.*�-�Qp���~�s|���A���e����Q�GǑȌ$:5�Ū9K��3��P�1�⟟h�+4��-	��il}	���	�
ɏ�AB�Z�G,z�&}��*�LW2I�ZG��lF|�f�4@��B�:Ff�������|C����W`,r��9\��i$��o�U��4u��Tʳ3z�)������k>���b�%1a'�er��c�Y�D6Q.X֘���3�$C	Ӕ���F��'�$��j���y �Y�O�i 6��).O}��M֓��Ä����(���C���(�'�v
���1��p�� ����N}p�1mEب�}�Ũ�uD��[��VTᦐ&	5��	�{��6Z�b�\
�m�V�XP��E��w�\e���K����>��ċ�����7����#���=i_��#�N����}�[���Q�]� ��L�K�_��
��������o'��Q"q����-�i��b�%��]�w�ʵ��t�SSNpn�7�+��qf^�u��Nx��(/�ѭ���.:����k�8�&&v����xE&Xk��QS�3>r�tA���;�7�.�@�&�޴���U�{8�����p��!���";���(����!:͠� �b`
+6S#!A0S����4��
��9� ��k	�1��r!���⽢�/�ٷ��[K����~�L[���eW������������� ��O����[�2{Ι�N�p���6�8��"�g��^<J��q�T	�0<��{/O��96y����s"��a=1���+��8Kg�cg�ذ�{��&�{�\��t�<o��͛��ӧ�)-Q3�� ��%G$�%Kpb��Ǹ��3��=��ʍ��?m����"8�e�ĸ�ꮽ��^�}��B��uR��u��ZD���jP;�<�L���7�q*��s����a�G���n�����m�:~�2]��p�"v�����թ�Yk�&��٨���<�L~�"V\�Ť� �8�&�w�@c�Q¨��za�\ᙏ�I	�bU���,g�8�D�ܫ��@"<�OR^��@K��������3�4"$ h�'�R���.J��NSe�b�:�-?�,�Vgt�Y�c
��?P�:1�~	r�G*��M�nd(�v"�,�x-!��a�����[��2�5�!6V�G� �Ӌ����n2�1u�; z<�w��dK�B�(4�[(���^ʱ�h��1�g��WԴ�Y�?�7���O�i��Uv��[���HG�z5���IѮ�=L�F�)�P��>�2�RM�$�P/��K��7�gi�5��2uJ���L\�X�ܛ�d��������a^�M�����1ь� K���~!q��� 
x\^HI��C1�GWh�[bL����-�N��K@�zw�mE�fR=T�����=�Z/(I��CD>G�)G.A�����w�%''�}�}NJ��.ݫ*.���[����`Mu9�m�	���s��kC�P��/f�'`kf�7�	o�f3.�[�/^w�=�;x����x�ߠ�񋣢B�smf�0�j.9�$O�^��$�����F����*���.���}k�6��^�b={��w�aӌ`O�T���>Di7����ؾ�Da��<�h�	�"�d�ͻވ'��6�(�^x��:}�W�eX�N+SҲ��B����Y>�� su�.0F�@�_iMŝ�)�?���;?�a�3c_e0}�5�9�*3ǈ@��y�=b5���g��q�����X�^In&��-�@>�z$�g�"��B�tO�Ã��A���*��Q H�ݿ:�VDbW� ă�p4��Y$�F]pw�gu�{"ѯ�{j"�w�z�$j�0¹�:V�ÿ=��s�o�jZ �+t� ًR�+�;�A���_e�d�;5,t��2��B��_8M��@(2-�ŜH�j%B�~�|$u=�<if�^�{���h!��0���;��L#����o��^����w�b�Z�|�E����P�Y���N��l���AE��U��&�q@|S�Y��Yq<ntD%O�� 8Bjt�[�L����F<���K�p;"1���W?��h�p�'R!�<��X�RX��5Z�����, ;�$�]*���y�����Q�v�dj���Tn���~3��^�k�� �]����k;&����F1�*' z�#ݮ^},�rd���+���8����vVk��G�d~Ԅ�.�T��3�Q��x�9|%�2G9�tw��tI�mTݒm�Lz�r��Dv;�g��h~fK�$ښ�����0��� �q1s�H9��S�Ӻ�yƙ����w"~0���Xb��Q�緷�+P.���|�u�W�O�Т��J���}
<��q�#�Epd��e�Mލ��N�	�ƇD_n�S��w��]B5�&\u��� p��e�c�8⪡�S��(�,�!
bE��U.Q�j���R��$���ժ��[��fi��B�-��2J��m���CK~Ǜ0"��}+1�����u�"�� �;�v��:�~��F�����M?o��]�p�´>/�Aq��*#�RL����BG�Z�yB�� ��S7M@(�䭂�qZU�'gJZ��쳰@£�:7-����l�nv�5��cc�L�j�w�����S����X���ή�[�wp59�l}KR8B���9\���O�I"1YE�Wh�y%t����b��z-U�Xw�[��,�t���_h9��4Egt��4Ebm��"����P�$�w^!~�5����
�W�����N��)#Rي&���v�4[��騶�V���˨=O��Z<X��KI�q��ږ?�YG�*�������b&,��#O�^����Z���_H M�İ-/u����\Ƒ����2���wW(�L�
��g;c#��' �	���WT�~��/�4iZ�b��.�J�3�ǳ�a��� �>��Q�.���y�1�����K�>>�F�/�H��b� �����==����!��j�@�Q��Y��	~ݏAd:�;l�p,-� �OV���Iw�b�)���,˶
(�+�0o>w�K��Z�8F��î��߈Á�9�S^���x��6�y�4;S@A{�`앁+O�Wы�^Zy����c�5��'�o��q9��Ŏ�� 9�N��:eB�H�����%�֥��I�IZ>ʆ�X"7"W���J%�1#
��I�F~yg�Źg���؃�ZwH�-Y�2�Lk-C�\0����u�jo:$�����#x1�H�W9�/D 9u���w��n�T��nb�1�0צ�����o�E��5�I��&u+��A=>��%,j�uF)s2���^gd��`�,�����s\VTg.��*��}�J��6gk�n`����\[wW�jwr;ƿL1=����eA�2O������7=��G�9�4�|Q���0'o���3�Lj6�7O��}-5�+�t�jj2և�nsko��?F�s`�]v$	e}*c�y���]�3�;�|$����|��b?��2��p��Uu���(�}CQ�/�نDC??q��ڶ��������]U���ry�}�:Z�x+
��ri~�y���[C��x���pq`m��Am����1Y/d# B�l�S�?���S�,�{�xR�d�`Lk��5��j�#�Ƥ?Q[[�L�����Ђ�3�Gŷ��(N�/4�V0���u�Zd~�E���I��f�8w{-�fN�~J��. �cb�jD��W�J�r͛��,���X��~�r�"r!���� J�'�vz�W��O�^n|���0�c�Y�=PT�/aǬ^��c����������e��6� �I�l	��*��,��=��فv�;r�/��Z!�?�eØӑS7�b��b��u���'��l�ܤ F<���Ks9h܎�)K��q���;b[�d5k���Mn�C%@Vʨ�	�>��5"�t�D�<bc��2Jj��$�����mz������M6�@aș��~v��y!�Yd�}�C ����c�g�o@|[�=ũ�V�n�g�����j���ǽ!~��2utp��fJd{��ց�>�{ɪ�N/�1uW �]E���YB>!�~{0?�B%���������T���	��ٿݳnL����-�,��h��¤��D�y�x]_[!}�B��U�'Ϡ<�����S�?������j c=1�!���6N��{�)0�PՉ�]�X��i���~��HNm[y�Zf2\�4CRԅ)8��a���V���E�Ȋ�j;��6��%�|l��`�C�Q�>ݔ�1��v��g���.�N��t&>��!�o�a���
��X�/b_zA��LuTb&��]���+Ƴw�鈻�E� ~�����Z1�ߑuAͿ��þ���z�k��>c!W�E{��,r�\�g7L��[�y����H���k�	؛ݟ��+H{�^�#���)}���=4���T-c�#xM�d<�	a� �G0��8�����C��)�p$��GimH�#��^`���S�+'qu����_7$��y�h�j�{�%��C�5|�iEHjDft�DT�����D�t�k�&Ya���4n����Q�u�y)�W�������[��.ϔ�u�[����rɒ�¬��i�:�j%)�E�O"Y��Ca
�;͋�^2텏�h3E�$�Փ�#�-A��!U�Q�1x�H�f�&|P)-����p���X��wg>�K^��"���R��K���J1�ٕ��HE���[���R�(�o�e����$߹��MJlK2zG�`0����$G`������;��c'�N���I��tS4��^��`TGk�ZAq'����=Q߿Lj�7}�R"�����r�Tl=��%�GNGjuo��HmP��Li;�҃.�*|�葹�=gp|@�w%`hV�}�&;Z� p��DFX'���>�.*On��y��P�5���GBm��������807[��@�&eɵ:�*�.;R�}N���i}7p�'0o�0�	C�85�޲����#���& �Ms�3����l�5��Py��HU`v���P��Fj2���������!
'���P�^1cF(A^�h�>�䖼8����!m���@�)�/��d��u�^�|�����B/T#j�k1�B#�\9�_������Q�1%�r)�9�XQ����YOp�@1��z�5�3��2#�)�c��$�E�[' dsNj�E~��n����X�4�{�=mN/�u/U�wl����(��_���� E[��ke|��_�YZ�U�>{' S��F��lcC+�`���W~�>,�vM��L����ߪ�6�M�N�^)����[�(iyZ5z"�#���H�t5f�(���7]�}2�$>2�LO�g�m=&d���{��H4|5pɋ�h��dϛ(��AL��i|7Xd����D:���~
�*�4|3�����~��"�(H� ;QG?���z�q+����t>�%�]�$��Pջ�Ne\B�.=�ֹ�6q�}������pHA�/����r�W��� �u>{����Sf�G/��I����
��è�,������z{PŮ��,(��d"��dj�_��v�$Y�����
4x��M[�
|����8D�9�� ��T�M�^A�"��=�O,��<[�Z��x>�ˢ`�S8.`��ABZ%"�_z	.%�}P��
FQ���xc��+�����	f�������Fq�se�(��#X��*y����q{� ��E�� ���X���T�Vi8�A[�����%�Q`Fa��d�B�6:E���ѐL.���w/�=��������[���|Hh(�{�W������{�?�V����Qė�~���$�Կԅ�zT�P�ד���ި'#Dģ2���лt����Betl����:A�T�0�0Pj^��B���_	�\Yy���Tc�8/m��͠���e�l�v0i�������v�Ȩ�i�eި�x�j�u�B)�+
�<��ܣ�<�V�W��=��s����|o9����|> ��a�472���-����]Bw&G}������l���L�}��)�1b�*�Z,��6B(*��PGÿGI�
��g`^��ߊ�?3!A�FC�fL��%RW����zAc������OIs1�!�+ �d9�y�I�m#9�?����� R8�E�Xl�IƖgM�aps�	��Hs�&��Q��[�cQ������Tj�9�:ޝ��c#+/.��vGMVu!���,��k�9��6��[�c�0.�} �iT���H���3��@��C��˄xU�O���MWb�=�Z�5_L?�4�qb�3�o�=�}� +f+J�7$g<c�78��H�v�F9-��b�����|&��\~}���a��MkmXU���cQ�~��I�Mt]1�ɑ@Z��{O�:h�G)��sf�U�6� ���1N���n�tGS�����E�������F�����RC<�2�g�}(7>zF�Q�.�������(5JF�y]�h����$I�f��jZ�18L�x k�8|���t�Ɔ�[�k�M|��i�
�r��")����R�~���P����S�Y�t�>�̂P�!��at�� J�j�Q��f�0��p��J�'�̾l���sr�Г�-��gȄ0����X٤#;�y%��ơ T3R�̶Đ�"�B��7�:�S<��ї\,t�t1���1��mz���XY�c �.�Z�Z�X�+	�?�*T'y�����$3�����+0��s�A���w]�����		EIv#�b���,�zd�c�*L�%����x��Q(v-��Eo�'���vO��)�<i��)>Iyτ�j���M���K'vɬF�D4�l/d�4�gV���/yq��8���q��J��K-��7��z�����q�I��^�d�ɜ�F�@�G_���T�<�?��n�ӂ�UI�r�D2�� �<�l�G���)�7 ��:� sϽ޼��O��S�R�S��OA����5t���f�R��?�	��!�w@�ٙ�/�ܳ�O:�֕ˋ���X���&a�+�ܫ�<�a�5��8`���������?K�d�v��SD_zim:kj��EC�������F�?N��v�%P��fF����.���W����n�yX����>��+$�U{]W�Ū���UbK{W�tH ���w�z���L"2S(]��6��M��Vt�h���V���I N6EB�6�gGe�*���7����P�
m�H:�������$�z3WU�tA;n�&<�&�;&9ŝf�2l\��W���W�Jl��s��#CF�Ĩ+Ӝ&�x������n�Gk�Z�̈I�e3x�S��A��3_t$&ɟG��N=���7���%�l��p�PQ���"0�ss8z67���?笗t55���2�	k֖afQ��S��IU)��1��qPf���s�4�M�>)�$��0
���|%�<U{i42I�K,闯P���A�"�����:���逛$!KְSXwb�=���wc���=c��ܮљ��s㵵�-�׷����}�\s͞AP��Q�eN��J'��b��� ыR�t�ܹv��|���Zd����Q�wŪ4߅?b���ꀜ��;�%����ɋ_�ْ_}S}HZR��|;�+@?D0J���Z�tX7R��HP�O�E����������fU&W/��\-���#ZҬ'��v�ͩe�}@�'2�E\�AE*h�!= 0*V"d
�㏩(�Z@,���ez'	�Lj�ˎ�� ���IE�jcC�|�}�e����,�E2��3+I���*g�ժǎ�{�34�������s�v���;�A�Ѥ���&r�H�f�Ƃ{h�-R֖^�a�S�	��S��˟�$���QJ��aW�-/� )���MP`�){eZT��gV�$��cf0� `��Q����,d�����VLT߶�"QZd1� @׻x���?��L5���b�p���m�ٿ	x��L�������
�^�I����u���wǧx�骿}I���\�;����P���a��F�٢#��ii��rD$�M��5�K�:�N��
���%{o�'�
��)�iL�i�68�;>�Eތ�;�C�X9d	�����pjH8�%�;������e�=�m.��Yx�܌֗Ï)�Q,��M��'����K9x���S�dα�t��ď4������aI�_*"��n����%euy|��PG$>�`�+YJ��m �Ǿ��L�_X��w�Dx��:���D���sS��~v>�lNl4	���"�ױoܨ�\�[�^1I�D�$��,��<R�uŹli�pS�G��5u�ǹ~^�ͪ�}�E0cج	����E�ܖ)	a���O2Y;�A:_9�-�{���c�����b�k0"�TZ�M5�Q�>��\%�������;C�=Q���]b�T��e�v bo�y"���}�����z�P#�K]��`������z�5{���(��r��qĠ �Q�}6gN�[���ʤ��#���J�H�T-��*�����mJ�V��E��R\d)%BwRGB��8��9xq�
��|~
;{�YF=�҆Z��ɢ��;BMJvdb�U���,O������èɛl}e��P�aR�^GJD_�Vv���������E�Z��G���"N��m.Z��T�� �� p��L�@M��^j�0DX�dp�,C\�ЧSd��I�ָ#�r�R�j'�����Y�E?h��l6dO�ӥ��6�(��	N��g�-�wۋ��\+���?���g�U�X�KB^����&v��4��'͡��Y�up-=�a���ڬ���o1����]�k�ިٜ�͔F��]M����Yjxٯ~L�hJi�I�S�LU�T�[��L���S�d�>Ԗ�5���S7,��o�ot�iEԈ��K%�H#��G��Ak�w�I����y �
�)nI�4��h}Ca~�vŽG���`қ,��~9{f7k5�Vq7� ��	L^� �J�ƾWJ)�8d�x���6�J끸" 9|지ާQ4)�49������/#�t�zD�߳tY�^��<7�lSr��C�b�����ꠌ����yF&�9�b'
9Id�������P?�:�����
!����B���Q�Z��C��7�Pһn�����*̜7B��.3x��`2E�8���$��Y����:��9��Ö,��)�ZF�'��H����X��A�e�6���2a����*��&�����Q�dy�m.� x<K~���o���$��P+��o'
�w>�b����9˸I�n��y����	���R�3N�:�Vu۟���	�J06��Ϥ����y ��:�s$	e�o�����䥬)��:���ŀӬ&x����\���=D۩3�� �9�t+f�;�R(_X��vH]\�^��j�%�����t@י�D���i)�E�?{1��pƄ�
Y*>���q�ߚ�:,xz
�9�	7`�ne<���q�>gyau0�k��X���K7ё(9�G��N ��̗*�����uۅz����>3�cx ΎqxM�B�m�6��c{Fd��W� c�+�Fkc�4���I�+��7V�1��ʋ�V��<��� ���y@4�I��JzG��N�ؖN�Dw�`�B����$� <���*���M��yx�~���K�_��i)�� Z���^��������i>�b��1���P^�mS
BN}���l̰㤟i�@ �j�S54n�A�S����L���gIZ_����=�漒����<�NÙ��U�5a�4=�� .�>a�w�U�N��v����	��GL�(^|�e-c�ImMׇ��`Y ������ݍ��G٣���4�J�y���3��h�G[/{H]6mk��|����&�I�t1j�t��.��T8^P���Ҧ��hl�~�CV��Z�� �l�$���O/�}��:L�����*� |�.�Tt��6�uo�<�\t�f���9ꝅ�"p/{������lP���Wo�%ykg{�%��ƼD�N�m��o�7Q���å��4�ˢ��35��x��q
Q���_��O?�1G�6!�GAm*�	ɍ$�\�9���yk�:t&^�DF*��Z�JW;�<��;{�B�AY�pz��M����:�ɈcLԃŖ��[܍MU1U�� *�*<^+��5��oq�vl�V��v�����&Eb<No�a�W66��[U���m���l֧�3RI����s����w^Ӟt��=՞=��~+�/�v�/�q��e��ݰXq�S��~������¢U��H���Dvy�'Y��)�L����}��+N�N���Z|�s w�B��Ŏ".V�K���p;�����S��׳��e�{�ׇE(�s/��2A�m�Q(�5nu4&��������⾿�����V�1?�������<N,�FfT��>�i�:ܚϴ�p�K�2�	_#���Y礅-ۘ���S�M��חٖkzn�`A��/1woՄ���zr&l.�h
��<��?tP��1;\){z}s�
��v �ƇQ�|�Dy
^YTJ�瀄S��_�����Ƹۊ�4�d��nX�ٝ�j$��l���x�����_,�� �ƻn6?����q���U$�iQ�]�
�3���)�!�//�r�3�G���T{c�ѣ�k�Ǣ��u t���C�ߞ~�<ƹz�V��I�ĭ6n���ޜhR���
v'��P̜��
b�^zUO킿{c��EcR��Z��/cT>�El������[ut!,��yr��D����-Dɓ]�a*�1�br�-��^�^�O����+�uwy䟁J ����c�,h���C�19?0�2��1s�����<@���^�C[7���-��Vv�1� �T�[HD�����ؗ�+����L(BZ�~�{L�_c_����6:�"�CE��B؀'A 3JY&}�=�B�0��@���ǗY���<�ٵ���e��j�:,��Oݍ<��� ��ԩ�-Bb�|��&�c���^a:�V/b-~z�y9)�pEϕ2s�r��)��4��%QJ��k����N����R�bVf�KYT8�'�av �X[���Ԟ�[l��~<����J+��}��X���wPA��?� �N]3LIs�FhCBW.���f����8����r@ت�^� ��nK�o�F���M�u�A����Q�Y�볎g���=������vRSJ��~�����A�6����'!�58`s�U+"��=��G�T��X��l�p�9_�a8إ5M�z��=t}c���W���~�_$���{����?����L�]��\���m #c�O�<�$	���+��bk�A�f���,������,�����pTF'�Y(]��˙�u��,I[PN���Ɨ�ɫz���ͼv�4��k�vk��gn�iT�����X��pAz�e��톨���D�� �Ҳn0�ST��
EJ9�N�Һ�}2�u+.�\�! (m���0��/k����uδ~ƵN�^�[�V�L1�V��.���M��C)�;'�3���B��G�a@�J�#�����:���<r=6��Z� [>�\7uM�ѫ+IG���S�E`CJa�o�K�O_
�do�li�d�{��`��fpvi>���%g��/��ejN�|-�D�`3eЩ�h��NDt�1V	kˆ�����l�.��'�p��Ƭ�Vc��g�°���̯��a��b�>)��uvy�&�L��h�Fv��-Y��G�-�S��<qav��ć@5���-1�����YR�v��y� 2R!9丄z��� ��vc_B���0��� ��&�S���g�	��Ր��O��nniD��e7%Ed�Tʺ�����o{5� ��n������ْ�_�x2�0�k[��rDQ5�͖wؚ�R�	���S�Ȏn��)�E�I�J������`SLxtQ��[�3�yM�f��G����~�k�Uj߽[5ڼ��m���1�w�q��U�+���i��k�YnKnp�yQ�8�(���
m��U�唹�I�b�qR@�#KAʽ[�����Ɛ̊�)���/�i�.�?*�a��V�&�G��sO�s�ͻ��,���qܰ,�>�������B"nܺ/������[~@��)�V�v�����}��yK�j�W�>ޣ�	0�+L./h��;���crӬ}8�AƲQP6m��..Ͷ�O�f�l�-�t��S��%y�Ev��9�*u�Jw9�{u ӕ\�b���Vw��k��`xa�k��,y��P�4���ēpb��.Lh6�ǌ2�b�����ɬG��,��*K�߭i�Uҝ�:� 8�yR"�Ga`�~u+Q��ok�t+ܠ$Zo����H���R��::+X@�����F\�t��L ��g*�R`.hz�fk�ծ�b����c����Y90�dU%�͸Ē���K׌c�������+g��E�A�0C���$������K��J��7GL���h��D�ڋ�#C2�h.,ݾ������d�H��m�~�Ë�Arv�Ow����25�f<.F%��'�|'�	P���͙,�/|b��j�[�w�_F]����4��BT����������c �}��3��ѐ`���-[�S��;WGn^!Z�q��8��d@�1�"cb�c���	f�٫%*9�Q��9h)o�il�f����#���=�3�4�0�f��vEb�o��>��b��}l�Rc&So#�����UaF�N&���@<�-�����|hxȭM��r���`wg��צ��v�ۜ�H�B��Ɩ)V��]�>�w�u��2���u}� 0��P�Z���l���r��._���9�[�Apd��џ}�R��
8U+m�Aʑs�ك#Hۙ�hՅ�<�� [C��j��v��.��p�H����j"m����L>fD^��)"$/�P[�1w�X��\v��ҫ珏�R�$0ȣ^Н"H�8#��[�%ǵ��ا3��e�ªצ�ӂ�?\vI���mEj���̕�^<�;(�ҾE>��=c^��f��;�tIq�P������nIMN8�}VMg&�I-�i������a&��]�Q��g��k��(�;y��:O�Мe�}����	�%�yܿ�CM<������(�^�jZ����ʷ����$T�g!OL�2�IES�9��4q�ma���\S���Y��1���a&bWL~����w-hl]�R��'�볝0�O[#wH�@��pV ڸ(�'���q����A3؇��y"v-�9�����W��m|T���4X�4��A�	���T<�+ ,Dn�s8[�"}o`s��(nv�]��%6d�4�dմL]��)d��<�ixR:���G��1�y��/�J$
���k��F����~�V&E�+n����a��acL��>(��5��Y`����T�<���H<�$�A�d}�:�m��M��C�/J�,Km�Bt���������'������<2&��ؚ� ������%��{�t�+/\{R�W��w��`N���{-����%�T��;b���y~(�ֳjk�W��q����*Dw����I�W4��K_{ֆ��w@��7Ac� ��J���v�>7���ҫ@d���T�w;��z�)�����NV*�h�>��TD|פ��	���r�I��9yF���z���C��B��<fkE�+7���Q&\����0��5����^�M��_�n٩r~l�1����鎺���R���\k�U^cA�Okz��SN ����ɼ�;�;�@����h}+�o��|Q�.������dI�Ds�ײkSlQǲ��D�kS��������j%<�-��y��kP� $H��&�|����Y� �GF��7
��e��@z�M��/��~؃R�Ս��-ڿ�̝c�Z��K)���r���*`��T9*�C=���hD��j%m���.�
����� �&R���m��rؒ���c�}YAP��?����&{T�)�E�K�9�<���5\�� ��Y4�ha�)���Ȍ����q����{nL�Z�����uAX�>_�|W�|*�Cz��XC���p������T����bFI/�4s��M�����`�g��=�c�
jA_�+�K�v}������h�����[���`�5��F+�`B)��-�+�sb9�#��W���gڳ#����MC˱.}\�Y��o �T�#@�t°���(-D��>u��xުFH��\����O=C�M@���k���	)F����Q�й�Q.#���������\����u�X����:ݾ�R�X0[_�5mj��\���i��g��i�l@���[S2�F���X�tQw-�c߲�{jE���G����俦�	6D�7��4f���T�'~S}�7-Nm	s/>ؗkv���q ��1�侞�0�ׯ�����1�-���<��;3���C*c�p������0K~���;��yaR�>�5Ҿ8�X���|�G�Cl�J���9�z��;}�L\hm�*��C ��������}�%l(~z���	�@�+�(��)F袗ɧ��}����Z��y3Bqڙ�hk-��E���#,���n_t��|��B��(��P��>pIy����4�_Q�Q`�=�����	&�3�%˜��o�U���#e�OB�Ѿ��A�pq��RpW.<����7��}jF�w����2]�'���뷝(�����S��pjtz��#��3�,Z��ax�!�nB.���bd���Ye!ռR���J����ξ�~���O�~��$\�h����R�m�lU&��)��b�C��'=�JP�%C����3��w˛��{v��C��[_R��a��A]ع�5n��A�$�8���h�Kj�KH�MC)�
�^��ᇣ/�#\�r�H��di��b�zh.�ټ���vF�I������:��,�a�+��iYf�p��U������oQ)�Z5A��2]1hh%c�vn�DD=ʽ���"�5d��
�����P�1��l~��sb1s"�<��ױk�����	���	O�"���8ģ����MK�z�����7k�vbsK5Q�\���j��݈{� nx3�{+bܸ��<�Z������T����lHA%� %{M��s��ttzl����naU.�ب�F�gC8o69v#2mo�2m��&w���o�.ǚPtԢ�)H1��d��D�@�7��{�-20�|�u��xC�[P����_|;��Nң堃�,�#P!ٿ#,�������Xl(���1��o{���3_���_Mm�N�~�4�������ܴ�~�i�wm�'��6��p��H�rm�ĺqJ�e'�� �	-RgD0"���ti��>j����9z�g��Ӊg�a��m�$��2��� f�����PK���a�1��L0�^�G�4Y�l4�	�i4R9�=3�"�nN��ը��j�n��Ҏ�*���5���xL�H]lB� �rkՈ���tj���W8�d2�D&88��剹�nb�bh�ܘV�*�s'��
ӽ�tl����_�{�m���2�һ��_�FS8TS�=M��?��-̅=�f�Sd�����4=�y��������o��7�iEǝ�_�3�QE
�Q>6~��1�|��3�
C֏�=�Ā�H��U-����ƾ�l��}���_�' ��?�@�O�R�V"g��V�P��)���&�G�����o6>Σ�ǭ�?u�<���H��%��H9��\O��D��w�3�����/��F�f�i���Sb��僝iv�%�������]֤
$/i�:Y�����!��1��á�z��nC��F��?�pK�,W�3 ��\��:Q�O������`|RBm���z��v-�Q�V��tަ �ړ�����#s6H����E������_�a��P��
 ���������wp�&r��E���bc���A�����]{���:��-|�c��\�`G�W����C�s�驼(5G�^��S�2������r`����B�URزͫ�X��� @��MrO�@��~GA*����+(����R�%�Px4l�$�_?FB��q�@m���"�g�1�!�D+M�ģד�v�	�ٶ/��I;�{t����Zq*,��h���Ք����䉦�]��I�)��/{�C^kHʑ�UIZ����;�G����o*i4����UgQ����tpʜ!���v�x��s�q�[�����\?3f�ѡ侘yrꋡ���#�bu�
��vj]��䏜�؉Xc��h����55��SrCq��}G����ֱ�m`JT{����Lm`��͂;���h�����Z��)~O��k��bC]�y��EM��2�^/��ZRG��7�!NV#v`c�et�,S�]��@0�#A�X}��)4�Dpe>4f=�6Y��X�~�aV�F����6Q���l�qS{�0���ܵVg/���Ç�V꯰0N��n�f�����G�k�6DE�����啹#��	fLc�U=�=�7��ݻ��:�j��{�fýI��U�|���Or��
�䩮���g*�}��i7��{�̍t�h���;�j]�C~Ԛw��b .a����Z�h�����W��K"����i����� %E�����ԛ��׻�!�gP~c�����vC��T�̮?�x��V	
M�=�LG�h��j��!��o˶�z!�}�j��8<M�K���m�6�B�R����ܛ�Y�Ѫ�m}�����JK���2�lC��z"�#nq#�
�ÿｨ�nZ��|u{7Cw�P_�H��׬kMet���#�>&�o�f�Oq�@�i�%��:P�.(������-����e�����%0�PS��j4�2i��P��؂�
q���Gz�Iʼϖ�/ h��)��^��]��ur��o������(Sd���nP��@>[ͤ۱�C�@�Uo44�p�4Ė^�:�ia3)ø����U��UM���%���?����`f����Z���dc���iz�P�,�|JX
Fd�QT�V��Cx�\e��Co��!8�cfV�˚P�Z]�W�B1y;�ê9����ZD���^��9�F��u�[K��1p3 �0���8�ߨ"���dí����L^V'�O\�H�ߊ�һ�n�G1P\!�O�K-F����	׀$�>+��&���M= V����f�fd[���(��(z�=��R�[�N�(�ĩGx�%���N�{��wT0L���Jڎ�~����P[Tةk���6�T@��5q��]��9%ܘ	0p��V g$� ��S���o���#�3�h�l���Za��^��vI��m}
Kҹ�'	-�ry��Qr!��cZ�|i���4f̊_)��T[�g頤�a6h�C4#uy|�E'it�� Jh�f@�S���xʛ"�����桋�_�&+�;�ص�E�("��EyWc���r}��tn�KP�N�lv�!�:k!�c�?)"����%�ҿ;��*�zNf{_�t�T�uRo�Q}�fw�O�����B�����^&�Х������^m�4yجVk�,)��͚3������	��Y� �3!��=������nZ�4>T�9�5͈^t�E�G<��C�Oi��v�D�%�{!�x���=�9�xg���j��pI2Zz9��5����J
t�	X�lg7I��Z�9�O�5�����Ea���a�-��F7��$S(�2&$����.q�+-��:��D�@M��J߸ظL&���0��q���E�i��>߆e��aTk�#A��@BBAF~���6�b���	���M��պYo��p���ѡ��[�C��nW��q��!9c.�%k�G���'��&ۤ����R/�	���T�.龌�!}eO��|��0�S�@蟍���\���p�Q��J� ����H�(�xV�
#Hsm�p��'�S�R'K�4`V��9�')��3:��;�]�l��+�a��eY��@X)`D���^W���Z|�7^);!��0����T7��B��7"qF�<�A�@��ݱK�]Ǥ頶�����x�	�ߣb��k��T��
�,���F�ޝmn���ג�hz�	h��dr$�����1��^Y�0�L�d%+���^��*�5�$bu�K�qh1�9��}��1��k�$�R��u�q��w��w�F�׿����^H�}Wb{���]�k�)�U�ƃ4�N�W��@�iӹ�$�kZ�32�_��/t^�n1��,��Z�~O
P0we�䌕���x,�O��,J5Y�Q�����˯��/&�^:,ar��\`����f��H\`KVQ��x���'�f�xs�6�Ӣ�F�b�u ̽ʭ.�)�]PŮ�;*Y�0�k4�����3�O8��8s�҈��z�G�]
��
���T0��d�?��O��������qŨ�v��!�ܹ�[�(�N��0�X����w2��FQ�o�;�&�"�l(�ο@#cO���O"<*��:�xx�fsEwD�h�jC�`��U�W���|����`_�v&������������;5/P�p���yq��� ���U���qG��YmrǬ�jK���|����S�"�P��S�c�E
�]��B�@}��u�N/�0h�J��A������uu�nd�a5[7��Y�C���q7/q.kV�~����RZ�Lܡ�=��vd�׺�zs"�Z����F0�󳉹q������[%-4<��<�o%_k����<���H�����i�ג72���n��=P<B,�d^H�/#�����]��^}���\4)���&��RS�.��5�")�H^��`���Q��&f�bh��A���`ُ������]E5E�K�������`� =�]�jX���������(�V�[�Y��ʔ:ƞ���J�>��� ^��)IWbdMk����u4oI�ܥ�*��k�Lu�ݗ\L��T�'���	��������9�*�/9/�6��1���u 9k�WU��jJ����4��\�<(��lau�K�)]���=��WPЅ8βIM6�Y?�iOvQ�
k��P���R:N��rl�9HDG�l_(�k?���>ۂ�0�m�R
G~)�,aA�մɛEC��<�\���ϥc�O���B��ӝ����Q��p��D(����0�y��c+��ݽ�%nOҭ�{E���l-�ϐ���؎����|,�D��ԭ��"]=�13%����"�D�>~gnN��AZ�����M��)}_*��H(d��I�j&G�U���1#��m<�� /<&Q&�k�ǲw����D��0�d�zZ��x<	T�������[��y �[P�)O�m�)s�Da�J��k�5b��WPc�����IUolۧ�Ig�T�QYH?x�!$�����bQ\�![� �}#|�8t)2��������u�,"8*��g��ƻ�┾��n�4!��}�}@����ȅ��1��:)�,7���7�p�BG��VTذm��N��'����8a��XX�G�1&{%�+��:�G��l���=!~��^g^~��Q',�;��K�a�ʶ��:��V6,�W��6��q���4
jJ�_J
�q�-�o������*'���*DyG��}WQ��!�m���n'�R͈�c�~��Z�pa�*̚��*���w"]N�s�)#�D6�	v|ρ16�T27Wu[Y���?�(�Z�ӋY�׊՗t�y;�b��l�;�龵����5bFU�<�s��9k<0�H_I!��|?�{������H��ȼew0�_#	垃a��Ozf}�h��О2��9݁���2���:�1�Z���~2* ��ҡr1�Eq�FԳQ$��7�*=d���3B޺u���$)�߇�s+I7�nǙXMށ�S�e}07��`�tUZ��\�r�Ϸb�R��~������ACkձ��#�췧.Z}�ӵ�$�o�/�|+��b��D�[h�.]�Ї�֣�>EQ�U�ZE�Џu��2�vF}�c�+P�: ��9.�X���09����G;+��R��WT�|]�ͩlK����kY(��O�9<Q:W�ÏA�k?Hf��i��_yW�������n3�i?�"��]C�F� ��xt�9��Q���!�iT'Ï��4��cd0d�u`�ړ��k�-PsMsyF��������U��(LHֹ��U�@Q�9tڸ����ANF-��sh�y�Hp�Av��EU��R�}4�??>M���Y��5CT]]���Љ'��HГ�"��LT�9�O��ַ�e�x�ƿ0���|��0 �[�dg.W�^�-\��E�Y�t�� ���)���8�[Ԥ0��tO�M��Q��kh���h�(L;�C���Aa����p��$sK�#n8��T5Q1K��8��T 5I������Di	�T�����۸��b��h�_��-�w����U���?t=g\���DV��Җ�Y��m�&B�m����c�v�:i�Q2~�\�k��ů��9����<SV���1�0�@}���r�g�:�'��IS���J� �9�1�k�-�b�#.)@�$�e>%�Um����(�>�������?� C�IK"ۧH^�P@�;�$
PW�қ{��q��v�־�^� �cݙ���G4=���7J�]g�ԎX��Ob��"�Ym���7���?d~٤(�)u���z
Sn�T$>�Sf:e�~���N5��|G�҄l�2�v2��%)��zNا�Zt��
&���ᇏ��ǻ4��̫�����+I���wl�����K�A��U�qX/����C�a8k�W��<VC��%UӅ1�uGFѹ>ށ��#΁����ao�A�Á2H.�f��� P�Ъɴ*ᒏO9�������i��F�q@5������=��V؁h=�Tq�L5u�����F?�
�D�4���t������U����{��.�Rf���#���y�L��h�=T,�4�v�.+���?�x��/_�^�� 5"2ᕎ��L��z��C0LI �rc��r�dO������/���?�g���O�?V�Sz��Da���P��F��H�'�H{W_%�ㄏ0��߀��Yx�9n(�U��J�����$P2��@k���;z�F�͋���WV�a��bz�V��W%��NIOl��C�Ӆf�W�2�������+R��I	 1�C��G-O�͢�0C�NvN�H��K�O��*"bzӥ9(���\BJ	�^�1(��L��dP�6�����r�����R7rvl�Ix���к�@*�� �.�1�zr�W�'�Gܥ�/9���#d+ʊ����nE���{j�)����hk�����%Fo\��+�M��ɢ���Y(o@�<k�� 	����C��>
�q-��=6�"^��/���,�_e
f��6�=(�;>�a�S�f�*�"�勗���#j�"����-��軤���;_/�i|zNK�d�qB�Cn��֊��z�w���:#��y/��T�}�YE_�M%ו�Yw����l]��/��#iC�'��OJ��{�"����4
u!$}?�=��KnOd �nF��K��r�&}�
�A�9���e8����+h	�}�-���\3iמ[�<�ْ�1�;����ĝྕ#�m���q����Ows�<A��ART��Cŷ����	�+.D��"8�Q� t�m�$�>���*<T��~���A۶�QgPh$��):gT;�����IC;sX��"�;��M���$	+��M<K8�Y/�(�NW��2���5����Շ�R���%��\�Y��kzQ�B�Z�(���ʰ�F;�Aߺ�J#�����52�B5��{�tJ���p�y���ߘ}�f��ҭ�V3�/��l���b\g����o�����w����ڇ9��4�ɟ�I�7����l9��c�D>z��$x�6+,x��PL�G�ғ�Up��ڣ���bN&��u(�s�����8wt�}$�u<9S�Q;�CK�s�0�&ͼkp��h��W��T�0`fA�6��� ��7r!Y�9�?pG�Ia�q�]�^��ZM}ɾ�y�j�!P��s#$�ߺ���`�ݲp<'{:_1f���e��m�t������rCm��b�ؖ^"�,STת�C�80W�o�F��4�ݞ��%W�����i�1�6.���.�#`��X���*꾌���&�K����T�5�ͨ����ڇԗ��+�����|X
?mk�S�z7����Z�}!��N�Gq��3B4J<t���{~����� ��FU
Q¼!� Mȡ9������;)5ۑM8��bw*�m�0\Y���U�Mڣ(��=0$�4f=�~���i�N�=ܯ�� ��勇Ʀ�5pPp��}y.�`P�,�%Zy�4D!����"<u��P��$g��������&\�=�sCƽٺ� ���҉�Fn~���F�8�������`�O^�2qOK��Xo�}�b�Y��P�ue./ �#��Ֆ~����a�$�KGz�Ö�?����i609�6Q\�:��
�hp,Ϻ�e�-����'ն:K�B�CVa�����=�</� O��RI,�EG�~ѐO$��4?]�@{}�����
/���%,4UVp{�� U��|
-S�!bQ��}��U�m�a ����8u�W�u(�O@cwJ���I��FM��� P�!�XSS�a��5�Λ�*�չ!��8���q�Jq�٤t�뻌<ח�|Ԕ��� �q�z�t�L�ڶN	J^*���k�����|ޠ���,BBm����}��-����9�����͇{�]����,h�e�[X��f�<Zvh���Ac�U�E��D͂sş�v��(���Ff��T�ݦSw����b:_i��RL�;��\ʰ���V�>��Qӹ��٦�i�^)��x���Տf,�	-�؍8'|A[�tǝ\3�ɇ8���z�S����0e�Nĩ�s��/�I|����%>U�7IYx3\�9q�|L����`+�(��|�MFpo�����@���6�_w�=���~Fx$$�f����<�h<Β�����f�A�e/����+����L.��dM���A
�<�hO�R���u'�o�\eZ[׌�T� C .l]��
B�Ū�e�/X�y}�[�AH���)C�x��C*�3���Э4M��r���џ����� ���ԡY�J��V��`���v��Ro�&��!oo�����kn��o�d_������js��ca<"����'0Ŵw9@/�(>��:���/��1m�2޻i'0�>LD���Y�l��kF� ��~Spp/��9A�m��'<*�D�W*��ԗ��_�C?�����ػ�)>������k��i9ᝩ�m�&��t��X3Y�P���0�Y '�O��̌��=�#��4�`�1��i�?R���u?&:v�m/{���d���3��kw���@տ�w�-�G-ˏ���.��.r�[�>���u��D+�XH��0���)��7���6��paI�б�w�O�-o0SB]�\}ŏ�5�4��YƄ�i`�3d����;e��� ���ET��q/=�0��o��x5��=��~I~8煟}���嬶��u��h�mA:����fW�v�/�	�ܖN�:���y![x¦����&%h�H�����K3�<��]�'���2�.��j{�������5�3d+`$��O�b}��yOd�Aa���29&��_L����3�B*]4XP���}<�V��Y�#{S�T0�T��D����Ҷ��l (�P���Z�4�94�*���4��-x���r0�����`NwF�G�������RU�ȱ�$g�5�	�p���������Y׸o�����!X��cK�;�q�^3��+�n�x9�X���W��o�;S�]��f��	Tu�j+�^0/JӕͭT��$umG�����dIh���ܦ��V{g���T�Q�%O�B��a5e�^���E�1��e���!h�s ^��	��eu�r�3g�"�w�hX�T��ۥvFl���#w� &���ڍ�O�]���,2�7仹ig�+C3���.��M3v׏lK&RQ��Z�������زm Vy9`�7�]��0��X�Wj��͌!��B��]��4&��j�w�'䅢u��}�=p/T�b3��&!0~R��& ��/�9 �>��w�ۛW9C����=��T�@,(b"��9D��fY�}WT'�1FF����z&�ĥ�3R0.��� j�=���f=�sN{�����!H�^b��N�_��
�M���F�>M��?��I�@(C�����U_�m	��y��N�{]OE��Km��;��\jkRjmQ�K�I�> cV?D1�a�Z!��9\&{1YՐF>$1I����v�����3�Ê|��������wJ�����a�ƭ4��P_ s��J�B��!d�����h전�F��؉!���.�4�_����$H���P�c4�8�ޏ����m�~O�y��f�֡�~@R��j��R�"��G��3yX�O�-3���-K�{>�F�*D����}P:	H8��M��A�+�yD=�(��H��?��|fU�JęT�(ƹ|�1B����3�?A)�=SX*�8}0駶�q2p�I����P]�w�;��5ٚ��[����x�ti�R1��;�e�?J��v�5�Ͷ2x�4n�qV(}�5��ҧ|E�ren��gd�Z}��0m<��W?,��;��/u�ŕԖ;J����#B�_r�k�G���)����A���L�\C[�16cUb�X�	]H{���!|�e�ªx��6�Ԩ̭-߅�07�����<S)5_��Yʣ�/:�U�jr[�
���l���q���k�d��%4,�Aֹ��nS�K����3��$�TJ�l]���qߊG�S�:���U��?=�wݸ]<��P���:�)�A���E�]��p��/Q6�_�L��|�M��&)@,) �UY�4N��%[膇�@t.�;iG�^�{X�{꺲�E�5+2��ɘ�-��ވ�Z�ɕ��`�F�a��Ed/E��y�Sm��G�r������ȫ�$��,��C�O�d�]F*�X���Xx�����g�mR|r���R�Lr���w^�.L�,2��p�X[KLj�N��)���rpl�x�����I��٤�Y���.���)��o4��DTwp��(6�q�I1��p���+Ȼ��4�2�Y��:��/�i.�
{���>�a~%Z��^�bK���Q
0&�-1Ǌ�H�'��"�w.�3�5"��������f�v�5���Cw��V����B���I9�� ���ݵXDFػ���)�3T`d~0i
G��_`�B : �v�3�_�3����+u�=�{N�V����R�^}@F�t�"(;�3Ug�e޿E7�B����lŃ< ��P>�Γ���I����=0Ƽh���ZD��x�~�‡�b���db� Y��o7a�@*�>��б,:t��H������b�=tY����[�N��~D�Y󚺜��Cx4`T�/yQ���Y�ͺPRF�QF�3F�7��fyO [Xc������@�{D�-"n�b�jQֺ�$19*l8Kz�p1p �|��_=��R9sFd\OA�cq�=�n�}��6pJ��X�����cDd}P�5c!�H�41uNX�;.4�$��&�J�C������'(�͎锩6�h��t�i�!��;�f�V�h�G��R2ʋ�٦}�dϏ@��� ���+�N@���<JS�*ڙlp��"v �&�$��v �T�U*3�*gmg
:>�R��П5�?\rڞo�{��M��k4���<zs.��#��9Ζ�`��˻B�H:�{x�})`� 锪�v�Y��ռ,�Ĺ�������؀������!�g�l����P, M��xP�J��]�i{W���_�lk�nZ5?��������qg�u.���I2I�2��4�:I��u�A���T�yi[~\�-���A��]s�{yq�
�۩<gh���}�k<��gz>Yb+��18�C��{b��Ac����=�#��*����mW�a��6}��i`��	���zȏ�w�ؿ6�F{��֭�Ttz��Q��D�2	�6��B�=-��O_�]��_�n)���*����N"w��u����E;���������F� (�1c&�Y��mH��-ܪ�|��"1�-��e�ݴᨒ:~��53�QV�Ij���i� aϲ����s ���c�L������I�Eg�jQ�
Ƹ�
'9@��dʴ�YD�dQ�Lټ�
��4z���� b&hı��{�e���ͫ��snl����<*q��Nkz���Rb�w%f}��)��/s�~UעjJ���	��M��K��5y!;�`�p߀�$ }�Ov��`r����5�����aj�*L�}�[(�n1zH�]�?l�X��P�ș$�|�����O�}���B��e$�s��,���K��Y�C�����,������3THn4'�0��N*�r�U�D�_ށ�%G���U���'����F��~��J�l��x�?�dD��=�<�aL���֬nu��8@"j�Kk�Ѿ(F��������0��:w��?�×���)�� S����'���zFד�8�,��*�&c��u�š��?GSI� _�#?52�9�#i�n):�.��Sٻ�d���j����Lɪ�y�K3B���Ȁ�B�2<3D���W�
��^7A�~���Ӗ3:zPi۴d���!'���Dez:Tğ�Ws�E���&BI7��Ƶ�.�q�Ľj�c#"�㗆��+co���M�K������]��Y��^�Cm�;,��&W�~�Tq�]���Z �"2ɖ�^l�R�?ҿ�3v,?�/�ڢ�n@D�ֺ���`�q���D2�'��%dIuV_j�l��񃲚�z{���T�w�W��+7�������iK˫]1X����{��B�`��i]v��m��&�h)K�5�Wo�W���o+�X��`�Xw�h�Ԥ.����={�����ǈkY��ԑ�G�TiT� �\�Vrs'bsR`��ۍ}�#u�kt%���٤K�ϔUt;�g�ǭ��|�WA�ou�(ؿ\����p��R9����'q�NWD����@Y*�;W�G�|�}�5�c��p��?��4�
Rrɶ��=�$Z��y�d$P5v���	���@�6?�mN��.�:3�Η*q���'<�lx	D1w�;�s��Yh�g��q�u�8��?��G��8޻�XۑӞ�\��yp\�ޟ����O�]b�*D�DIO�0�_�L&��}"^}{��8��w��B�W��/��d��I�;E�n]��;׍i9���o�	� �)|�|���;�B�xm��Ll��i�D+��x-7߰�*�FT}���1�i)��X�����E6\�y4�#oN)�$�\���z�?� ����2W�#U�"�IA'�B=C�.��}�1��"�>��q U3l��5@>�!=>5�d k�Q�g+qn�Z��N��$H7՘�ӗ�)���������4�_��tE+?������Ƃ�-�k��g	�q%s�����>WF�㽐��T-_U�G�n�rYF�a�B�M�QZfNk���H�xV���\ ��^-���D�7O=W �&�%�xW����! ?�bBbDA󻕊����ϊ���أZ������N㏅�����Q���3�L:�怌q�"yjNП1ɢ֖.p)�e쬖ޜ��nF��x;"N�@XA��|����U����Ƶ2W�T�6;I�nrp��%	�kj��;Ҋ~E�K�����DuP�
2��|��GG�c�ƹ�h74�.�`�Ơ5�a�M��u�?W�����$2tíJXJzla��m#f CG&���'�(o��!؃�g��(M�U�f#6߰��YDa���p"��(�j������.I�n����OSz�e�}bX�T����� �U��}f��iitq�]���K���q����0�ɥn�;U���[�Ӎsp	��H����U����=�Fs��|�������T�[����<m���#J*�'�	t��;��%B�A¶W �\�P���Ȋ���a�S��q=���6�7���>���%>a����3�𡝫[�*u�|v�׷��0 ȍ[����S8������a3s���lP$J�t;c.v��*T}���,�U���w��8�J�f��	C�����WF�����f�w��%h�]�D�Y����A�m�f�GK�\Т�͞�"C�Q�chh�d�?G�c�wH��ya|�� ��C<:�/4ʶ�2牲�C#d43]5`�:�/E�K��c�������)Ǐܵx�c<��ѾU�KI�����i��*vp�yDFӱc�?��y���7�?$1���_l��ԇ���V���/��!6���΁�R쨖V�ct3s��A�}@&������b��-sV&���@�$��O_���V��z%��R3��\U��|}"�޻&��F[x�p#��8!=;t�`#�wV���Oo�]�+>djKzo�蹖�|�4�/ϓ���k�a����&3��RPFM�wU�xO'���1ob����Z���,7C���>�N��]PX;4pc��L�J�Ӻ���@S$�Z�+�R����nBi	vW}�'f�^�٠(� &�$SA;h~ՠj�� ��ݲy5I��͡�p<�H�&^'�~�D�	 �7E�D;Hc:Lh\��!�!]x�*�5����+D����k��.�3}Y�Ӟ���&n�]t�����&%J9�~��������籝�!���6�4N�x��!��������[�_��*���SNӄ�P#��Ȳ��>��DD�ɭ�BGclIuiBj�Ԫ�g��"��&BX�FZ�q��G�D���]��ݵEt;�6��!6cn��F��g&!
M�滷&\.m���z��:����*�#O�C��EM\��b�fS��[�ٙ)� #�T�H�s=���c�??$oXy���%��.�01��!w�L�J�5U�i��0֏�k�p���RJٹq�m���&�ڏ{��M3Mi�g����⚠����qV��+���C��%�*��-"@_q���,�p�)FM6��>z�mح�o짓��d��N@��>o]���/�}y��������!��6U��~���Z��Xߢ��:H�N�Qy�z��wܼF��HS'Xa��:i@��a��0�����<P�� �nj@T:պ�aqOBݠMI��s[��k/
q��YO�:�N�
����e�̚��v����'�8QUeQ=�	n�3�ż 4UC����?�Ϙ�]�L�s����|���ӑ�=}:�� E���묵^�f�յ��(�R��UU�
3����Ev��c3�93p����(\�����(�7�JЕ,�;�]3v�ؗ��-�|?���gg��b��`�6a5���}��[o!/�*�z��*Q��ۅ��v�ܾ���$� ^	nąjk:̤�	*|n���<�o��a�d�`Ę�-�|���<��a���\�M}«>��	o>޷��\3�����]������L���L�&�L��f�h�����nTW��ٽ��a�&>�;�Ő\��#j:k�\�VtⅣ�X
y���97��rY3)LՍK�sJ�F�����U���|�ߟ<^W��pk����K�/G+��8�o��?�VG�_1GVa�p��;�K�"(e�܏񀺴����/��;}�9kP�N����D�
��"�i����<
�a��҂���v����3Z-�C�rCؠp$������LFx����v)��Ū�h��^���I$6�`��5�����ԉ���W���	����W��Jj������^���֥]�+��ö>�s@h��������:�V� �/W�Mr�����U�h0���]��w��vg	�9;�'�H��g-��.�1� !�#Ұ��X"R%)��љ!�(4M�B��o��J:�a��R��r�^gO��B��M����ԬI�v���rT#>>B[|+�-�#�n�u���X������
�x�e��+e���V���So����[m��9ui���$_��l�0������͔uvuA�6x�;��t��7$.�s�e�v��9�uq���v2�}��6��y�Ԩ����9�3�*��5�Uz?�~4�aW�M��7�W\���E�_���<Bys�o���C���!j������*Ǎ/�3�er�Fo0��ł�Ο3�gG�W�7]��g�,�}\m���U��8<��:q����'��R�5`��>���D��
b���4���p�m	�DL�G���Da0�H�:���'�[Ϲ��V��2�.�LI��������f���8�=Nl�s�o��H~����,���4[�zH���[��Y�,��%���b��!�j��7�ް@��*�}p'lXl1}��о��x!��T=�hy������䯸�yQ�!�s����>��?�(%�
\!��q'�)Q-�.��M ���T~�(�s�R6�lUn�g�%���,|"�Z��.f�ZCP�2�7y�8�����EU�㥯�ɰ$ko�B�èK��(G�j�a8��oʂ�1�L%AJ3�<�P��Yn�m�zw���Us�/(~�e��g�)@~��T�8T�Pl���m�[T��&�$��'�� k���8,�Nл��}�`h�"6��2R��:��`;q�kQ*5z=�4z�̻4�[�bp vWk@�T)�?��Α�IU�_bv\1�Ľ�X�4 7#�_A�1�1��栎�h�忟������p:ë9�כV~i3�NM�ɿW�+K5�"K7�b��hx�9��Y-y�z�$����;����73����|�����`�ޞ
��LN3 GЊF�y�pm�?M _7y����۠����#����(]D�{�X�9�m#��Bg���h��}��}�aB�{��[���8�$��d�����Y������wo�4�z���{̮B���|4�) ȃ
u��6|���ԤQ'��B�<���%6�r�WX&(	��m��{4kV��	!>��f �.ώA�_D�/b������tf��"�A��2��a�#~XܡX�1B���>����V��� 	�Sc��(�"�V��~J�t\ ��x�⿮U�X"����+2l�y�"�T`?M�FY��Q���BB��u��Iݠ2�g�OHY��ѥ˒Y��X��{6�,w9;��m�Y���m��zT�HQ���*�,���7����Q?�r�S%4�V� Rj0�9�r�)���m;�s��;|tA�m�i ��)��6�b�q��($9����i���^:� =��8f_h��`.j��B�c*ʏ���5?���u�����܌(C[XN��6j�*�B�F�Í �U�_�9��Q*/���\]5l�eY�12�L�?���tw����8�x�́1�]JU赑���i��7;�9���_���o�s�ԃ1X	ev�l�+��leo�ݍ��V��Bx����
���eLf\*t�,�MPb2?B�/1؂l<Q��dF*�*U�ȵ{ۿ)��ʲW���i���wd�9�f�f��W�g�����i�S����%��a*e
t6m��PRH�6�tx )��#;��˜���;�rO��B��w�U��͇�y�`�*mc>g�O$X>�Oc�N~Y�Y�T�b��ﲝ�ql��|��f�N���s��*\}yPESC��B"��jS�������N�K�%�hW����N�c/4冭�Vf*�Z}�[�����jEGr��'n��=��x��":�����mN����V����*��"�ZJ�yt�1��)��i�Uu��/�3C5���6d2	�`ZE��6x�c�XZy����t�Jb��w�� O���{*&� �`��$T]%G���΢�Yf��{�jC��o2 [�`U�'��g�dOC\����$ �i�lIa�uu}M��q#�VY��9L�ؑ���`��Oy�)=��S�n7������a6�`[W�����]U�S�3��[�bɍ�ҕN'���B�����x�~(�I�Q�ݶ��!ٕփ"X]Δ�(� �Y9�{��p%��a�hWٵ�L��X&���:�
�O;�'�c�.�i�\�L)˲�593o�P�N���.2�DSlϧ�Q��`�9��1�e���Ӕ�٠��f-�\^n	�R��ۄ��Ґ�oY���(�v��ۻힷЉU6y'}E~n{?�tc�t�:���%�EncA�_�0�#�e�uno4����뎙�]���M��`qz�ءM��'H����0i<�+���F��N�ݧ��A/R��-H�Q#�IHk�M�u7�B�E��*#�����d�$$�+�+�����:���o��=th�/����
`IZ]^�&�d��%�5oJ�늖B$��?���+:k}��C��4t:�oAɞʡΥ���1w��q*�ʭ�*7�����!�r��0<'����%a��A�����A�a�9���]D��lrz�}{�h����*R�X�s���+)qnh��d�߈�Ħu��V�>A��QK�}�K�����nB�T]aPI�c����K��]r���ġ.����7��|\}�ժ�i���'�mI̲)�m��ƃ��Gϛ�I�&��`�,-�j��"X!��ĕ��p^C����T凛 �_X����h���~Ј�0g.sB��:;M��T��>u����upJ�,�!
h�oG	�t���L��"�:���#)=~�ǖ4�0d'�-2��޿���`x+�*%7��~ơb�"�S=��}m��{x�"����b,HHe�a+� a��:[A���6D��"�|L����Y�iti��ڄ=�x�K(�~�R�����y�mW�����{��|4�6�=x)�efۋ��>�!q��|�+�;:m�����b�7&�ǈk���<�FsY�2SSQr:xRBg�L�k$�ק+���x�=���񿗥�tUU���9Yf9�aJF�*����gr/e�v���]��Kn� �#zv�Jy^Q7�<�r�#�H�����8n�p�z0��P�j9��R�>+��`4_��~D�~~��b�V�|�Ieq'��)�t����ҩ�;����Af@O \O�po�'���� ;�2�lqG���(�i'�����?N�����5+�������*�\Z��"�x�X~�q���ܤ�̃B���н�{��PV����2@> kYGvx��LWkȹ����Qyp���-�f�$ԏ�����ųx9��idJ+�|M0���f_9�U��B��}3&�'o0���SC�Z�>'kэ��F�)g��������.�_3,�uYw��Զ\�R�as�eYچU�<ǝ��׸Lk)aU �3�]ߓC5xg1���Bؤ���qN4bV���LI�Dn쪘4}X�b(]�2���E�L�dJ~��Q�����r�#̯�t��a�V ���; �/�W�Ϻ�j�����V-^��x�����s)]�^��B9����K/1��J�|�BW�b�+N��8#��:����6ޅ*��1ЭSMY�4��+�Ǥ�,z��;�=4���������^֘�	�,�zo���!{��潾�h�M#tM�3��v��P��'pI�z�#ȉ�Z�T9��QĆ|���r�K����c�Ϋ����"HXϻ�����>)�~�8*f�|:��\�q�COJ.��%�c5�f��u����O��!�m��oYp�)�
��=2t#q�1	����q&�	��� md"6��P�7���/��~�_��P��'(�瘼"�c�Y��߽1�SV��ь�CE���"U�=�zi,���qS#����@K��vͿ���4t	��Vr�G���7��M\ڨ��#��o�I��f��[�����7��kg���,g���`(1����ˀ���S!i�\4� G�r�w�4���S���^�VT�X��uk}P>���fjA�l��clP��'��xK�ޒ��U!�_�>M�Ҟ�gӹ��6�S��dr��Du��q� f�n+:r�f7��TXT�gٸ��v�Cq:�Fl�,zPq�+��^�Q����<1 |
4d6�C��q��;��ʜ� �.�KP�f�b���ޣ�+9�����ޞR��v?3�G���S�}��St�O۽ eN$��zg�h��|{l�!Q�Z�3�Ѧ#�!x���/�PxAOMz@.'!�^z$_v0'�,H�(bb�K
�0���nk2?5S�&K4(� ��g�^r����y�C3�ΐF�_W��$Rd�Y{����+�H1T�K���w��Di��v�vr#KMe̊B�	0�\|������X�Uؓ�uێ�ǟ�\ҜR��P�GMZ��%��D�U����3T���M0���v��T��4��.��G}��NO0�"�� ϱ�p?ȶD�����Zw���.��SFDk:e��ia�Zm`VB=E�{�����NK<υ��Hlv�F�B��h��Qi|�����[����.�~��Cx�y������i=-Ǟ$�8�) ���VH����gZDN����~���\��J �1�Pt��w�oq�,������jN�D��� �̧�-}���.���|��c�&����`m �>4;],��,;�h��,��Y��Z��&�.��D��b��8����UH�
�Uک��1�!g����Ya>�����V���R��ߦ���l3��Q�P��hj��F�a�a��V���|q�DU`��蛍h=o���</�p⧵�6�0���>��,�@S��9�[���}46B3ISpHu?$�.�qOr�jU�&]�� ��w[ߊP�JOV�����1�c���6�F����`��s���N�pF��<�QY�	�jf�%�R C2�"����9oC��Vm�hoJ�}����~C��q�f�(_rߞ��PiW���o�EH��-kH�H�%��;Nۣ��ѯn�<)>�v�"��u)�9Qyi��_��X���uK� �r!�^�C
�{�ˀ�fP˛��k˝FS�&���Z�����;��;8v�=��eŦ��k�		�� &7C r	�}��a��+�r����������^r�Э�/���U�<�@tבs}OPίy�5��F�����3B�0���Øg%@i���kR�zV}�~��5~�Z�b�TH�S�;��g7�a��͓0���q�U��9I�� H��!c,��9bEi�Y��-���m~k��f�[�d$�]��Q�fݜE�
d1�1!?�	~��L0~w�mi�ZD����Z��T���,@���BRQjX�!�WY0���;� ms�J'��H��\P����>�xQ�ݿ�)��]"X�M�e1`C��M�b����[T����9=�;�|�IV~B�1���'%�1�����.�1/��"C4y������Sp���z�#]�A9����\�5	X�rK@r6\��ۮ:�o�U]�JX��s�;�JJCY8 q�����el� ���a�F������UpW�\o���2P��>6v�M�����'��_F��f��2>73�EZ^�xe�T������A��C�VE�?{'�	)�(��C=q`�:A�U�r�A�l?S_����s�l"C�e �=]*�@�Qq��X�w0ٙ2
UC�r��c���Pӓ�M!@�]L���T�z�h�e:�r�s�6�1(�z����_�9�@`�=�,P���~��e��[	H�+���k�o�]�&��I��2�uq��<�]�s�m�ɮL�Y�WVF1١j{��03��M�����,?�>gf�n#],%B��R���fxgY]�m��՟�Y#�Kk���T�>�}��|�F{/�o��j�Q�)��#_g�Q�Uȉ�+)_�ǟ���`�@�m�Ճ���=(�o��k5���Aћj^,_T]	�{�a_�TNU��jU�a������e���(���C4��5��J�;��451��߂���f����מT-�9�,B���"�T���Rˁd�]�[03��t a`�1���6����i���\����0�/��WWZ`)�d��B��9� �(����Ƹ�����:
���{E	�
���1��������7+��l�8����ޥ�*���k	��*u�εt7���pV�ɂ����!ʐ�ٱ8#�`9,غC��T �t��V9�����g�M�mkj�:Pz��'�/ز��Q]��x�#���B�ș-T_�L�* �F�}�JE"�g�ì��(8������h
]���_bD��hOs����a+ �a�;<� �JF�ċ�V;��IZ,�O����L�u�9Eh��&Zd�ݜ�>�_��x>2�c+kƮ1���C�*�P�]w�m}h#��
��NU��8͆�w�r�FmJ�ˢ���0R���`�XF�)�>_7sg~�0#G�k��a<�I��%������.���"���6q!��Щ��&{��y���d������=W�����z��#�$gB�
��H����
h*��你iff�^@�xrN�+�4��ЎI%\��[M�}�r�o� *l&P XӢKȝg)��RZ��\�A�0�U`������G�%�M�61n�,V�9k�NT;)v�$a+�Ad�3��j2�sE�xgP=(�O��Э��;����wc�<�n�Y<�]�;��	}�`Z�q9$5��Wv�n7:�'���F�d�'�0���?���(`MSv�ҫ>0!�vY�ɰ̧��!'	��}�'�Q_�$F��H/Iz_��j��
�����w�Iw^������|�
��s�y_��wQ[�7<��bJ���kX��'�Ց���Jl�qB��">���	'��d�w�-�h�2 �p��O5�j�iQbnպ蔅�(.*z:��+H4�.�&�]"]2���+^x\��p����u�֚{�,��
:جձ��R�4Ṕnߜy�&��gT�d������1P
���Zag�m؋�#a����J ��e'�i&B�8,��l+far�oaHg$�G]
�r�PpM�v�C�۷� ʝh�L*�S�x���0S/nb�l�L����j�0��^�b����i��%3��ml<�N� ����!b�j���҂��\(e�4N��O��v���>�舄u��y3��K<P��y�A����s�e��6�]��ܯ���b$]��=/�8�b���	P� ��R�oB�'f�:�,31ڻ�&�ET/��[)4���~	7��_��y��b�7�fP��h���4��\V^�ara�)aH����~!��2�v@���A3x��h���2[|��DڶH�����f7�rT��k�5�]��C�pu������o�f��{�#��Dc�	�"M�1�ћ��S��Ṏa��fń/MO�ǣh��%�D�'���:f/k7����jӱ~`Z$(D��AQ�>�^��I͒S��S�*t�8w�]r�S��#H�h����`�.���2���0l�鴪�����
'ܑZ?�F���GR|ѻ~.�E3郦4cAv?�t��p��(�+�{���_��`�G��|G��̶�����P(��C\z�sn�-*��%2q���6C	�L�3� �Om�:ĔfX|��������Ѵâ]�����b���*�{���lR���"Է�b>ɬ2T�
�C%�J��u�A�d��z��^һY)[q$8J��*���..&q�BB����[�XQ#L�d����#�����'׍d곌cx/��܁K��m�4���$ی�X�R��L��3�mF��Б��M�$C�)P=R������bb�dR�'�qK��� P��m�P��s�­'�fM��L?��f���3x�{����֊���!�4
�b�::4�V�&u/�{��,>s3=�/��S9��v쯃;��f��Ô�6��\b�}T�iK�dB`�g�sZ7́�G��5-��j*c
�n����p�AQ�E���@�+�_�:9��&;q �u�:$݇��#��h7���)�)�S�5ׁ������h�@T&8J�F��Z��e�re�b��]E�w#3L��A������2�t��Il����=*@
j���oi{�iU�׏�V��t��Fd_�����OZ,��>7� ��]2.nJ�?��������y����"}�����9���mE����p�p-N���̻ S3�\�`BO�L�(�&� O��p(��ٝu��~V�w%o�ۖ+RտoI�У���\�cp����p�*��E��o$Ӛi[�,���Q04~� 1G�ܩ%w��)[s�X�w��yۉF�R�/�k�d����<����Vb�|�Ͼ�*2�����;ۭ���?f=彮k�J�I�?��i��)�18*#�?�zoI6(4YNh��ok�C���!���8���
�%���L�!�@��/�P��Q���o~۰���,q�Qq�k���'g��Ѷ�w�����'��6(��k�sB_�R&�]u��Z����kɓ}\�?����C`4�ڣ���B���ܩ�G�%�-~0�w"�+�g�MB���v:?C *0�
]�<ꎪn��w�C��:�c���a����D�R����ԑ�ϐ9�\�fKh9i{��F����$�g��dxdM�O�d�e� ���	��L�Kq��e6.n�Ј�C��1��+��%i���FG��uq(��v| �Ɍ�*����0l�~_�2��i��z!�Ð�z�6t\Y{n�q*�\��N%*�ֻ���+��}ð��D�^k}�����Wh-��#�?`��E��3�r�:ٰRv��L؛k��V�
��1
���  d�6d�tE�쾱A����!$�����c���k�������O�#���%��6��ِ��h�ɣo���ḓx �&�Nբ�r%}���È�_i��Zq���ȥp^���t����F��<�E"�l'�4!U��~R���#��Ԃ緲>��42]�������;�)D�#���_�>6�w̏�R���/��?O�/�|YR�| �	���+f�Q'���k���#d�G��w[���}jRw�&��0�HT(�����㓤u����
Y�v�%��ڭ.�F.�k`�X������(��5��͘�ӳ�[��z�f�J����8j,�P2��b=l;�k��+K�Yt�P6�&#�t�/C;�-��;mڎWH���#<]�j���TnY�Zc�)zr	5T��/��RF`a���ܳ$�RR��@mWE�lS�㞑f1���AEST�j�1zLwX��)X̄ż��;������pc����ݧDy"'�����������^>h��7p�;�Nan�^R��D�������v*��].ܛb:����Mz��]q#a4���z������%n���1r	}^�g:qU�DͰ���\��u�j���tՎs�ׄ�����N �麲˴���b:w�*����a���%�5����������i!U�战A�5l-��]! ���i�yYwQ�����?����c��GH�%�c��x=�8l�Zp�'bw�U]��;�y1O�&ڳş�����`\>pD�������6��Y�U��U�����\ؘæi$�UXՄ�	#���L/���i
`�t��!�f��ï����R�߉}���"���m�Y̹�	�_,#K}�׳�󌃋��?�3�4�j�m�Rg� U�}�?�j��,����Y�� ��J���F��F����P\-�F77j0��_�<�ʆ�ʊ��uӠ�:u�k:�����7�|�7}
�n��-}���>��8�x�������x������[}Y{������\ƶ�D�φ��%���o����/�$Y��Q�L5c�f5�DvuL.���O�uƁ*��Un��$��\z�ʊM����YH��K�vl�ڢ�}�dO:�U�45PC�>R�U�8���%�G�M:�k�Q�5�-K��������k���Ȑ;�X�c�҇��!�}z̓]C��k,]R%t�$�z.���*���IhS�� I��X�w��-�%q7�aP<���y�-�SW��{9�⠙"2��ǹ�ǐ=����B�Gl!��eq2�o7�x�3�\�^a�Ɉ�֡��e� �v��t��O�#��,;N��R���Ggs�g0�q�:S&��:W�w��o'���/w29��5�]���榑e�*Wo�p'��nז��@o�W{
�S��X�����tI%P8�࿛q\دMiʟW4����	6#�XS+'�����*q�f9�$��.B�
Ek��Y��B�y5G}�R"I��6��F��Qp"(�_T�l7T1"�q M���p�QZ��C��<t8Mi!�IU ��I�c�򄪫�v�ڹ�(S�c16��U�[�b��Z�/#�^�E'�$h3�]`<d'�Q����A���eQ
?��K�-���`9*��F�xs��TkTh�R/��ؕ�KS܎�ĕ�Q�-����+��º.`�N�}/��0�D����`�O��Zqz1��&(':w>�N��Q^��8)xX(����<)��
�ڢέ��v~�\����D0���c[=��
2a� !'"��a0�,�!OQ�a�o~��],���-h�� G�p\n>�0��աL(�oH��1P�`��Q���n~����]��{����*f"L{���^�)p��N�Dh�%�h�˞��N�-/Z���6�6Iό�%�7��ny�1��]��۔��`B{U<t���&�fEz ��2b�q@m/��G�����n�%�x���Z*��������N��K�Rѷ�LFY\fZ-:(;�M ��,\Ƹ�aA���B��h���Y1\c[�"W�x�}N��:fE(|*�@�V�{�-�a�[�g��#w��T�i	8��IcǋÌT���5��A�{a	ǉ��$��$��^<L��+!�J������2�e&�Q��֣����?(��1��I�V���\�@����[�Vdm58/w+1HH�ƺ{�sIoo�����<�i�j�������� M4N}eJ{c�57�^��YXR�6�S�w��*v!���q�f88��ӧ�!O�f
A�|�Os�^��w13ϴ��ϵ�{�4��g�AЦ��b*J��속�84�$�
M�\4s��贕��_��b��l��ko�����/���'l���zN���áy
��/�:��(��k���l��4�D��7n[iY��trq����+B�$mj�0r��*�pT�,����<��z����7t"ƨ�3o�g_��`J�if`	��>������"&�Q�X"1�:�G��4wLR�Od]rRɫFŗx�!��aO{2)�P!��?���TQ>��e�2��o���f�'�]�>U��OBh�Xq���3\����.5�߉��G��<�q{[m��G<b8Vq
��A��ǈ�{D8P��a�=�xU�w����8	��4�(�J��h��G���O*sbJ*�@�T&q�5���y�"�- h��"��@7XGc�ּa��%�1�?{$*���.�z���W���1F�}�ve�X�5���KH���������>J���.*O�0��0��0o�� B~H'�2b�SJU��lgң�v�f��8����H>o��&yL}E!-�zKc�`��1SI�&���'���sv��z��m չ4��޼fj���"\
5`�%^���-��!s�������\M�d�Y�w��3'M��l��`)�Aԇ�{�>��J{�Vc[>��C�zu0�K,$�D^��Y�|�&��i0@�P��eXgf_��`~l�-����;�l�NE.�f�;/P�2�)��0��ST��q�+a_d�Τ��s2��w�R��J����\յ��>��w�d�r<ŘÑ�ۯr˰�^�ޣ��u�\z2����3(�ۇy�7W�è����.ɯ>#1 e,�g����tTƦ3qND�-'���{����ʍ����,+Z^{�����(];��:!��n�W�b���,��4�̫��k��*�����Tky�מ_
�#��ݕ�@�(�z���K�]�Q�)�ݜ����O΋�3�+�
�a���_�,y!��v�s�B����p#�Q=�)I�����݌�+�?�~'ޓT��|X�s��	���+��95���5�}�D�u��z���m�� ��M�����]J���.�tQ��z F��"墵�@��c��o���L�m�6��Ȃ�����l�`t	lQ]�-5#$�TU�9+"Ŋ*	�������`�Fw��!��^lsh����	�����U���OQe.[���Ec�57�����$Hhŏ�Ap�H��o5��N �$峠��=�V�|��[y�,V����JM� �bE�����7�4Ԟ�?���0��N����z+d$�_exQ�u�m����o���5�r�]^��6��Y��������&}���-����?�R"��3�{o?3��@h��}~
����xj�1��S��2���Iq��Y���i��?��A��%�19�Y�A���(�c�B�evȷ��ٳ9�.��M�ⰨM�^������<]q6���>�w	$5<k�2[:�޲�Տ6��*͝;�S_O�%�Xe�!b�_�xtB�B@I7�\Y�����.Yo�1�3���Y�o� o��η�Q!�	���:&֩�P/E�H��.�㪯��\!�z��ɡ��O/~P2����>��;�5�j��RLvNx�{�*��9I����o#�,OS����������i����R�`�CB*?pFV�2z�wW�ڳ޷D��KR��-E5b���P5<� +�r�ut�^[6G������~+Тr]��!I_�\�G�m��{H�AjQ���}�E�#��pɰ��B�v��Y�����y�Q�K���_bZ����K�J>|���Ö���Dk-.f0�G{��oC���Q>N>@3�ڢꬑ�1b����&c�g�����/O��i���z�cc�A�䇟4@`O����w=�p2e����[���;u�q:a�D|%���9a}Oh�I���ƺ�G �wkG��Y%o�]M񊤘�(���(6�+3�����`x�o��-+�<�B+��:�\�3�~�ҫ��%����}f@*��H�J`��뜭�f���ZF]�d����4�W�~U\�Lҕ�Dcz�
.��w���9y�A����:��{1#�9��3��[��|���C���4�\;�6��.�4@Jڏ�-��j�g��ۧ)R��ȋ��\X��o��*�*G�����Y"I�@�5"�V��Zځ\���
���z�vlj����c�v
S�A��)��,P�������X�i��wc[d��P�k�J��\�5�d�@�[?aJSqO}P�E��޲`*��x�WDަ�B	�����Ц��+�V@M_�	g�����sU��j��|N~���h:18q��ʩ�`�6?:5{
T��4���B�-�?|���R:1�>�Y(����H���?� $�P?=#ۃ�ɁƱ-�N��V��ZN�ˎ���/�އ�2��<N�놞b@!B�/�;j6S2��������
��W(K\4d<0��+�G���4E�����)���T�ݾ��<P(W���yӰ���b�+��]������ݑxe��R�5��a�Do�yo�nJs��rCR姵�?��	�[3�{�Y��@�\@�5�s����kk�*�+g�����F�L���1A�z}3���;�a�$��\��:����o�ȣ�KJ:�u��1�i��?b��b�x=�T'J�}#SN�ނݪ�5��g{Qg�$�?s%DS��R(yV�4j��7Qqk��ǭ�m��@��} D�8U�nd 1���4�uK�v��g؟�!������Hbrɺ��t~�Qpȇ���J�Mܬ��	�ؿ��s��u�J�.ϙ���Q�e延����k��9>C�ӯ<g�h��HQv���ʝt�u]����:|�%�d��?��z����-2+�l,
�%�E,�jj���c�tUږ�ƃ�sˋ��ETA&r��w#=��4�,���>^� [���ٱ�YX������n�E\ժ�7Ӿ'w�.�yqc�/WIݨ�=0�t�N/���0BI�dIJd��wt���בֿ�!h�Ι�1�4$��eu{�H���ya|����-�3���9�"iwpG�O�'"����
f���?X�&`y$�0@lM�X:
f������w[�PvE��n��%d���Ÿ�WR�\5�y~�NZ�'���%�3�f�Y��5����ϗ��6��	_t`��.و����C�c��R�%���Jod�O{њ���P������Q�p�B��w''�Jm共��JA��f���������)�ߔ�� 4c5�݌7�4����ؙ�J,e�����	���Y�ո���[���r�[�FhH����ܘ�WP����??rKEW�[;��wF�A>�+�w����Ď.dj̟��$�:]��^L*吕 ��*��l;*`��kNTF���/��q/t}/b�p�X���T�%d�]7��4W��U\Ix	F<q$�����O^Y���u�(��#I��*���R3Qi��.Fs�<�0 �H�:M�Vn�����oWdpǽ�	8xa��,�	��.`��e����Z����<EEi6$� L������Q$��c��9�����Q�s�T$j������-��F>}WƑ�d5v���'���*��q��+���=gK����������J�,����Pؿ��٥���i� ��jS^�-�2��T��lZx-���Y����2G�I))�t�=��u|��i���c/��������!_���ќF��L���;�n�m��5(�]��f��s�=,H�>�[�*yB�BD'~����:�=j���KN��:Ya���&=�q0��ښ����QA�,-2?�wW^��B���!��u�#�Q��&Y�ړ�a�����gCd��w=��86��U՘@tC���Y0#����!��E��'P�'���@Q����J~�s9����ؔ
5�Z�P/�iY���Ѿ�s�yw���k���_fE�|����E��{G>e��}�	64K���;��/��8~�<t��|�.�o��X���4��^�
�x:+4�z�Ū%�;C�KV����!6?Y���_0v����5�R�ٽ�w>k;K�8f��ޛ�fmK�" ��>�mC�3YQ������ٝ��Bb���0OZ��F�^��+��P��W���xɲ��=y(̗�A�4U`B�+rE?N��~�~Ä��HU��,�����o"x}s�H��Bs"آ(:<�D��j*n��>B"e��0��}'���X9y���6ⷓ���վ[yՔ�uSAԋQ��<~Z	MTچ�E.�7��rNrh��Vٱ&(8�Pmm��+���l؝Կt���{�_�|K�}c�LM��*s8FF;�A:�a�Jژ���� �܀!$�F�����hj�g)��E�|6���6�g~7T�e�C,�y����A�@Vܤ�� ��<L��<0�qG�ߜ@������}V]�H�z<f�9�t��r�b�{{Ս�q�jM�{��5���4"���W\��9��r��'��,���h���$��%A�ܩA+zs��ǚ�,��*�m�Q�1m��g�oyw̞@v&Ģ�w�8�0A�A[�����<����, i��O��2��w�m�����,V2 .=0Jx�Pԝc�x_<�G"�X�E ��h�&�%y��ǝ.$?�nБ���Ȳ�T��2�p�1vJx�=�l�ɣ�]!."Ų�驉TK~�#��}srQ+c�JC��� 'N%�=�O�b�nvM�"c����*�*HXu��߱7N�����S<d�?O�����:`m���G���<���|$����+S�.�Q_�ʭ*�n�ֲ��*�8�YU6���f�SIә}�=����͸��8U�x+��K��;�F!y�U0&�o0��r�0�y�}�[���d��ͧ�y��Zh��Gl�g� ��az�7���G;�4Ms��k�xR�[M��.㏟���<Wv���$����e��x~��֯�N�˲�9����� �P8��3D����Cpi^(�\�CN���}8Ɩ( u/Z��::��U4-�pZ�ɪ�'��1����HZ��󢨨=˓��@$�a�	00��J	�br��X���atg#Q�E�������������c`5�)v��2��.;�Z�?�NM��Y���Y������Q���#��d+��r�uf@�~�h>��h�� ��n��*OG���{DV�?	�}�ڰA`'�B�ol��!O��,���ii��-�P��L�^��)�:��f�r}ή�%jp<��˛�I�r�u�ژm?�W���v^�����#�|�.�>���<��įH�ɐ��i���hw~D0�%T�j0��Q�vջ�B�Їa�����Pq�~�?cD����;�Zx@��e�����ϸX�����X�y1{yT�X�`�h[H9������� �$��E�-zc�'���7����p�����>*u#)�3�@L�����Д��#���;�Y�"��#�{R����2]D��n�L�`C��a�[K�JZ�N�ͣ�
,͎A�����/e�����ƥr�nTf�P��Պ?ߝM�)�����[3!�r�C���eǼ}���"��uaP���j��̈́1l�� �(��U�m���H����q��6���lQq#�?qm���0���{��AL�E��J�ǃU'�m��Zx~��pX���m�O����\�uͷ�e�n��^e3�Fڳ����%��t�рϝHp{��>�g�C�eP�7��B葒&�0a>Iu���ձ��ƴ�: ��i�خ�n4{zz���=��픇6@��cM��Q��u[��ᜡ�C��׺t�
=+Ζ����ۚU�M�Bi���<�Qy
`�j�+s(�4i?��/,�]�����.���p� L�6cjO��)�i�}�X�_������9B�Ҏ ��`=�7H�U��S�S�G��1�1�0sE͌�]^r�4$�	Ve��C��|�(r���|�D"5v�����ރي���(�~�Q'b��\�(w
�C�>��w��KlL'[#�Z�'�|��4B��w�v�	ښ�Q��'/z��w;�d��2���1���j�9��=��"<���֪a��U����Q���������7��-��:f�Sn�S��.�@�R�pG�c:>Y�Z�]o��N�9R�.^��ͲPtU����(�B`'PC#���V���y���d�Tb���s)F���b�S������Z��H����}1���=�9S(�gK8�������x>��~�˭/���[��an���f����ZȤ4�?T�刧��Kk-��D�':�(y<���Z�@��V&{՝(��gʵ����8h20�*_�(�
ZO�ʨy|
��	��!�b梤�5G/2t@�'��#�v���
�9�$Xp"��p� Vd�6y)p�[���T���C�~D-�Q�4�����$Ϫ����٭B���wX���i��uF���=Z~V��Ӛw:��;Z�5DI�Pk+4k��^熥& �Nڔs�G!��1���h?��I�zZ���@+x�2�_]�G�/%��8����H&�9�w�
Г�X��\�_��C�������l.�� v�0!�nIJ�6�NA�<���e�����|�����Pei!!��E�*�z����7a��t��[� 4�l�a�� |��~��翷���Q�S̾+�?ݼ�w�NӄO��6?�z|uI���
�c� �u�����E�2P�'��MrRɩ���
Fh�݆���6.��u�v��ؕ�m��6�����Q�ԀV/�3;=�M`&N�v�>~������%���h�sO b.S�r���Wi���͛`�(32�U���j˳NT��n���>>� }(Q��"5w-}�e.>E��^J[F��JI/ʃe7A�e�m�椥�{���d붫^��?�t���r�$���l+І�N���p���Z����\6dv����+}��*�k�T��$i�����~�Ӗ��$l׀���[MՋ�������J�Y��7�f<����d�� @=ж��x��j[VռP�l���ܕ˰Y[�#�M�iC��e.��E�����`%��G��Wݘ�Tn*�� �K�f�&n��i	y>��Lq�T�O���[䵹���	��V��BZb�@_Mj��޿.�9�d�~4���]>� �5p9��_~"`��ȫ�%��
�FUi�t�k!0���Ơ�z^x_�Mw����&��A��R֩V/��#e�?�Z���o�8�� s[�puS��V;��?��lڻ�ld��r�'h�̈́�ێ4P�c��V�b�Ch����V�]�GO4 ZP�PgiV����W��3J O�0����RT���
E� ,#��M��p#Zϵ�Cf�W�9�z��g�ñ��'�fl�Y(�[���Eb�2�N��I�EO��'K��x.=��������3MؙD�L�jD����X;��Ug=�s[ܜ#���9�#@T+��3w)Jq��4�ѯ<v����.��w�͏����&Q�@$�uuJ���|5#��'���ot|�V<HM����w�;EL������/Mf�EH��p�D��9;��0�ᏏΣ���C�w����KO�٬w|�U����ZC�G2� ��&',�ht.î��T�\׸B���D�0G׋��Qo�+�\^a2�+q��/����(ȥbz��zyPM�s�x���]���U����,���3rO�Yj�sJ`��P��	_��A��Z�-�2߭D��E�`��\��`��os�#�̅�#��δ�*���વ��~�����lu�<�`Q�9�8B�qck�E!3�\Zv[��I��1��,�*n⺧Bd(��%T�,�i2+�'ֵ�y�I_�l͐�7�b�y�k�ԆNe�@��4M̤C���7���ܟ����>~��V4�X��#l�`W����l��X�gY.e|�~�9s�!����EB+�f����I'*�����dC,���� �&�#on�/�Y���cX+�J'Q�ڌ{{9��E*E��T_-���' ����H$�s��~�$����<�p��+�pu�MC�F�߬Kӷ�P'�VNf�����71�\�/]��ip���1W�5�!��L�R����d�3�1�q��`A�i�%G��,1�7r5�2x��xe�X��J�/��ڎ�Ǵ�ܭ�KMdX�G�MxP<�U0a�kyʓ7�`��\��Kbj��f��82���{�t��GZ�y��}�����d\�{e�x��ad�f4�']�ˢ��k{��-E[r za�J��	W�f�à�$��
v�n�4Mx��!�!~@'����H�_���[׉��{�Ha���~6�ų\b���\
�Q �`S�>�A�����D��@��y*�/,��S.5��摧�ƛa���M�^E��t	�D�f!{&߈TGj؆�
����;[�R��y�R7BW�4x/b��!==k W<ώ�r��х0Q'�xؕ�y ��ԩ��L�G-M+Z�����������e��J�-T(LT+�'�d~�"0���$�gZ����VT_��v,�H�O��4��u�$8d�^򷅿n�~�~v��n�n�Z
4�_�T�$_��kZ4c@B?8���6
�%p"�rUkk@�� ���Q^9t����PxA�OdB�$�m��y��=
�*,�Ҕ{�*�,�����9�c8o��e���sѾ�eԬć��r��Q�H�h�/�{쥂���^���GL���4B�u#FA"�4�)�~�=�Nc�2T�^xs�s|��%���8��f�Q�۴��A</�X�{r:u1# ��͆ٻ�O�q�Hm�D�q�Ϗ߿5�`]�2�$�t�;c�y���ѝ���bo����jƵ������Sg�۝^^`lPq�]�ϊ��+��h|�|%�`�2GL����Y'�n�3i/���-l"ϚM?^�q�ƃs���k9�y�����k�<Tl�k�(�lP���.aUe8]����(���F�C]E� ��YY��'��ݏ7�[,�[�6��|��\��6�b,�x���:�4����7��{;����V�<wO�߱�D-�.�ru�I�x�=�̝H�Fp���Qu8(IAK0�,:��
�q6���b*���;��n�pl�
ѳ$;.f�Z�&���1��[��摶k�:�! �򇝖�sӸ82H�FD����pxp�'2tT!����v�yW�ݣ���/6��r3���5Sޙ6�b�Z���*�V����JJ~fݖ���f�|��!�)�#'�zH���������$R�:ib�+�M�!U-2ޞ��do��G��$> �զ@�5N���7�gd�l�����ȅ9��.���n ����߻K��aZj7��x�KD�
3?f<Z���r0t;
�ŚU�'c�4�:{<\;%=wT���&7;ذ�	�3Pf���/�DAN�n�9����/��G}���y���2�L���'�un�k5�4���0�k������=$|�8���8L��&�eF�G�-����cJ����;��2�'�����4�i�O��OZ�R`1�N��j�ӎ�;=*,��0�=�%�4s�-$��/�9V�;�7z�Ei(0�� �,,FY�"�}�����3,�������V��!2'	x-�*o*�&��E��g�Yo�E��Ƈ���������������X��X�r�³qܾ�+�b��Ƹ�˽~:�j!���+F~����;ۡܚ�C�0�ׂ�Ƹ2���j�\��k�u�$9!D��o�==���W�;�"S��~��y�v�6�	�wE��l�|�`r�S&2�c�O_������ݞPVr��<*��U�U`W3dp#�U���I��q��B���q�8j�a��8��aAPT����F*dv�q�G�4�41{M��4�{���L�WN�D��a�o�v.|D��+��$��;��*��<����l�B�0��UV̿b�k�?)�'�E�tϭ�
��E21����֗*t��3?]álJ�����ڳ��+WHPAd~t��2�c+P}�4=�՗ ��K�s5-�b(.v�2������x�^�K������>I3�s��Xnm��kJ�5��+��{�bvj���N���Ñ��\���S��ѢK�s������c�����g������'/�T��'��4"8��@v��ԕ��KK�[�3GP����)q�"��h��?-���)J�sg?��/O�dq8F��h��p-�^����/�زEk���~v"IP�#�ʾ/٘H��bΜ&$s\MG���)����K����r�� ��(���=�gb(��Ӭ��ޅx6%��<���@*�5OP-6�d����t\	���}�T�MM=�V���&�hڼ}Ơ�a�Ug�9�Ov��)��A�̍���R���x�I�����`�j0� �4���kg�+3�1E���k
��̻3��<��O���jǢ�����I�]�t��������'g�?�1��EK&T�WxK�H)5mG�����E�G|��:������S����L7g�12YK"�./��k[�f.����:��lCk9let1�E���:�� 27I�8���[�c��h��"&�&JupEi�C�x�ug �%�"�GE9�e���K���Fa��h��yr��i9C
s݅�枿���C�\���*������Զ�$ �g�S0����͎10���Df'(���
���1'`5��h �viB�c`�z� ��L+�����r0�[nf�0���������@�\U��% t�6��ĥ}G�,>ZA��M�	c����uS����C_,@��`8���į�^�^��)�3���X�i"h��C��<�R�g+�tǚdX<����ַ�f1Q@�I�I~WcSf4�ZV8�����B�̲$%��
gg�!��*�;[FH�/���q�'�ece7�>�RϹ�:���z��ϥ���yd~eeu�r)pQ�7��sLՔ[������!�Gd��3$�J�d,����gs���:=����
�g���D�
��aHqj����Q�3��U�*q+�+�<d�g�Xh��������s�ae��f='�]��������U~wAҥ���"����"0i����TK��f8���p�P���&l�%B�(7AP�)K9M`9��<�Q��rq��4%4��{Q�rQ��@\�~��n����^�ȯl?a������2!LSb;m��r�:z��S���8#U��,��2iWt��>��~���^�~�`�e8�V�⛋�t�h�T�B�SN��0���J�}]&�2��T����,�e��X��2%����v�=j(w�j���1�<��}0Gv�g��!y��B�4�[���	�m��苍}pDh�v�7<-)O%×���F��m�,�'��H�ӭ�)� ~��v�A#}�k����R.�4c;�c��C4nM�̂��p�ID��m����L�v�>���{Zr�LB�/�ZI�mX/x�W�>��\E[� &�D�Sg��2��.Дk���z@�
6Z&�)H�x��l�����c�%r\�!Ugym#���A�!#WcZY�Գμ��5@Ίuw���i) #M��.��V���	����ʭ�`*8Ԧd���:��+A��&9�*��@���S%;'�W��tl�E���c#j�v���eν0��Ԡ+���bKPr�S^F�]�e
9r�݈Z�4��?o��ٜ��q��
�$0��R���<a���"�����$w��S>�(�8����߽����ޡ��p�+��p����+K;�����.���I�tﬢ٬������}n�7��sB�*X�i���ǈ�ƒf+U��S{N������M�g���O�e�M��B��-�ʍ{�EUc�� S�f;��=n�8��X0,��n��T��(��i�|b�p�(�퇷�>y�G�o�|�ʎ�^࡮ʜ���x��A�~�u
��M'�=ߋ�L�\�XiY�X�[�6 � 7��u�t��8^����B�����B��\l�gh:�oI���c��/�r����Z��΃˥:���̆`�ӱ�a	�$}�`���Z�ief<��8%m����Mj�.i �0���ֈ�X>��s/Ͱ���e��� l.I��T!e�E \{dQ���܁�#Q\�F4b2����0������B��m�՚Ciݹ�h�B������u�J¬�(����r��B	-��Ҧ=Q��6�Xe���k���J�J�p������I��@���T�����8�%���.Ng�L�Id�R�iP�WC�@x��s��H�ۮ��!.�Yq����-~�9�����ݪY�� ~2�������K�Ϋő	ΐ���}���$Lׄc?鍱�9��~'���$H���58I�"�	""�W�F=E����5;�S9��%w�t���'E�lG��ju�1��,ăVF�5�3�=�y4čg[=�j��#uW��8���my�qhkֳ�l	[?�a������͚�T�� F�u�`�I��f�����s>KE�Q�$⭑;8�iT�t����t|����<�4."W�(�n4��`/ֶ�G�^+�(1�$X%�K5�B���ӈHص�n��F��U	�BUÍ5��杨
��R��-����Tl�)�Z�5@ңA�t��;xK���Ji��Z�P9I5_Ś�����6�L�h�i�l��̚f�U{��<Ⱥ������:�Xw]��r���X������F	Y:���0��9�m��'��m@�m� 8Jan&L��ƙ����D#K��2���3<�$~c7wd$%.��bl��h������r��~���-��/�7k7�5�ȁ�8�.~�O��k�M��n����X;D[�4	<b>���mj�
z��/FI�UF6����]��z�W&+���/ϓ���t����k>��ĸ�j�d믪�q�(p����$r��E�}=Z�<�-,<��̌x�;���j�q�!э��٫Yos�<�	�r50Z�$`�K[��x���V�<d�b�|66��Ѵ�5~�{A2�&�cv�1@5�5�׻S��ũܙm�ق;%Ԙ|5/`\p�����龒ށ��]NR0��|8�r7�c po>M��C@��Z~�%�!�������'������*�w��Ґ����hbt;�l!���
8��+��b�\[Z��\��P�BX'�x�~��9�߈������I�F|�̳��y!�&�� WΨx���E��ka��t���{�"ʚ��va2OW������rupr��f�G�dD��]H^%�َ�?����;�A-I���n�ۜ�7� z3��J1���X�c�`���6�Æ�R�,R>Ea�8�P�g�/�E.��y�4)�Ǹ����vb��kP����6�%%��j�6u�Y`#�&�Y��#����L��g�{�B���#�qоV�׏u�F7�L)hN*��.zt�ѱ�U��]m��]yٲ�%���Vj7b�%��+��?F*q�v����KRcrJ����c�:Z]�� �yO�.;|'N�`��U~ڟˊV~�2�,
��~�
ˆ���3x6p���I�����f�mp�L���O޺:����:�&7%��l�y�bG;�drO?gSH�R��p �	VD�4P^i�?�|�}h�@ʹIr��ԾU��� �qX���O
G�тOoC�TR��+�	�\��	��n�Ç K�h�������~���Ս�b�ʏɄ�e�ȥ��M��W�j��W$��G)%�|�����Q�Ć��i��.�1��[�s��RYl��k"X�D?�Oz��U�����_��4�ǫ�r��e@	��E�C&�)�G�?�p��4՝��j)���0����l<g����x��F�%����u��ݕ9_lz}J�ɮ{O5XQrd��&F锻����,�Y����m���k5Џ�a,#~%/l����Q�B`�E@/��dD����Y�JR�]5a�~��\���~/1��ѡ���ϗ��E��!�Z�KS���AV|��]r	%�O�T���0ڼ�0~���<ʈ���/����1X �-����徟c��t��l5ǪN��s��ݝc7�Cp�g�_X�<�XD�ڣ�� ��9��h��e	v��qbB��K~�$���HL�l��R΀�j���<r����@�M2�9��;�<���`��n]9i�J�+�V� ���9�$F��hGΡ|�;ؤ8k\���a�f7c�3Ӏyj  ±I�������`7C�R�w$�B���
;J�/V�{���#��k��^T�X�m�ƣY��;
�9}���fm>6�+�~V�D��(�������G|�zҩZ�pnu�%Eb�p}��������*�vņ��y��J���"���e �'�2X�e�Z��M�.�ĥ��n��iУ��t��p�r�1�l��"����|����ό\|�h��u����&q����Q�C�NbJ�����%�ެ���a ��P~�C~u�c;s��R�J|(�OŢ�G����{��`z���?�����詥����g9,�H$���!�P�H�^�1;|��'���k�#��O,�փΡ@�Q��3f�z�]����H����$�d�+H�(�I���i�Ƴ�$>*@�G+j��9�ῡ�!Z*g��=������� ����]����k+%��m�&F�=k��g�E�׺�pESR�������0����̤��3+W�~H�|~d�Q��-�τ�S����*@�#��b4����<�K�W� FM��3����>s��|TPfZ;Y���}�L��?�@�����H��`D�nR�(q��p�ᕌ���l}����06@\����!�jn���i)Hmg$Yrq����
����i D����%l[	���h>��+��8 �3���߃�BO؊!}O4Y%� ���|K�ͅ��}V|��	9��k��P��%O�e^{OJ� ���U��Į�v�wHe��ˀ|��8��^������z��4l�z1aA#��f�k�ڎ��US�T�c�������v�!(�?�R��?�]��Z/R�����M|]�E�Xj�D0[p�%q'/{īi�% YT�dE������-n/��x��71���*؂C}m�i|C�Ђ��ԣ�1�c:�5���k��djF!�2UD�&�;��z�0g�Z�u_bcj�o�m�VMT�L���ʯ���T��5���J�J�|F%��҃ॹ b2�Ӫ@�,��LTg�{Q�����
��������Jv,Ʈk��Vu��'4�Ku��G�29��@!�3&�WxDc1N�U9M����~�Ӊ�r��s�Jʖ�t�V6���L$@WA0�kn��{+)����2kK/:�`�+t3�)b�R�ہ1{0k]�����ZM��g�s4_�d�����me��+?u*9��ސ�<�F��V2J9 f%�t����x�ᖌkEm���1���m�R薕�7�I�N��ˢ���fc%�b0�>��3��턠��ۄY��`0�C�|:d���':^ν�����)��Ҏ�1���g{��=��zN��ʍY
��G4��gc�9�M������Kf���1*jm��;>Tع9S�Rj3���/5�U����׻(�A�@���W����!U����d/���c }i��w�9����wg�É�y�n��*/�g�v�t�ؼP�j �ɉE�e'��^-���v��D=��$`��+���ՠTRՍ�!L�]U����_0p�	L>�.������S�25f��p�\I�iq���*���_*B�IU��͒�t�m2��B�����c��GR�LɾLx���P?zSYr��&� ���K��B#y����1��޴A[�]o7�/Q6i�5��q�g��9̈́񴋸*�Ʒ���z�^[�y�K��R���F�9޺2�V��Z��2�q3v":3'�#�O#�$1&%�~���~�h���U��7�i?�;��GE�pC����:��� ��H\��l�O:�cz
��Z(�I��j��n��xo��q��Zˆ�hy��6{}���O��|�I�h�V��_���`�8��@y��(�|��#�b��/rf��<aeԜ��d�1�ovh��AT1�,� �O�����2@5=���ʥׄ�����?���z	RP�F���.�s*Sk@���I��gf� ��al���H��K�<ZY���6mŷkI��Y,�
�MZ� ��q JӥŴ:w�4�:�'���;��!˧��N�PQן[�>��U��ڏ(A�����O�Z�V`�Ցf�Ƕ5ޯ:��0���ō��	�[e��,�Ҥ"��^�%��� b�XJG`*�ΊA����`ö�iÌ�>��i��g��5SA�_��&��R�|+Q�5�s��:~%��W͗0�/^�X�w�N�Az�֎n��ތօnX�,�t���R�>�W��p	w� ����T��%l=/��iT�����#��;N��E����nSeV���u���fa95�aM�;pm�$��Il�B	�I_*__��6��� @��$d�}�e9J ����i"�/ ��?i:b�.e�c�@%%el��KZG��)cE�������A��"*�o�i�J�<�Do�/�TΣ�ܐ���-�k0��9d���K]��$b�Р�(9=���¼�:!�}qv\�9 �7_�
m��W2��.��n�s�9�����w��� >�O�[�H0D�wG��ą�EA��d~x���`\�\(4�c�܃� (��|�\���/�������2C8ޤ����G��x�����p@�׽F7%9�5�f?�jp*F�@���6��|�����e�
�(ԭ����c
V |�EY��ˇt�$�Բ��v�P邌mr� �U:"�J����$54t=zة�P�����������~��_|jC��vq��n�V��n=��\���8'��ISׅ6�
Y7cظ8Ck7�������Ē]5ŭؼ����'��Q�p*�nu�����Ԣ,w��i�9Gݨ�®��{եܰ�X���q���}��U_���X��M��d5�G(@�Ng����' �����r�#��r�yӘ,����e��Ā���X�=�Is/:�RZ�uk�f�r�C��i(�(!MҺ���Q�A��t�t'�2��+��k��������p�������QF���*�eu�u�`�3t��ͼl6��!��(~Q�hb�m�@��Ajfg���	�Byӹ��s Rba/�1�m�Ku�j=uQ��$z.=%�����hYŐ�x�0��*��u�T�����;�8f��ڈޭ�7x�n��4o[*<a���r% ����煥�K@����������.��xĻ{Н	���v(�8�İ��q/�,�X��o񪞝'�s�b��B�~��q�9򪳅���[���}��>�4,ZT��@�v�BA�±�y����W=	Ց�<9��?����X�dٷ���	�ТK�qis���`�� ����e���	��Ëg�8���ɍ�c�+hE��7q�O ��Iz���a���̙���D�����u@�0[-��0�N>Q�'��]��!V�^K�HA��BP�kF�b|[��z�((O5-�뗧���Z=b�ܸ��,��A�Q�9i$�~�	��0�����Y�� pU�=Z\�g��Zd��=8id9���yu {��!�aS�y",-����������������5�<u�p\��}A�dV�ՇNr�P��R�f��]��dD����'+%T���\]5"'8�9��֓��.���Q��+g���Hq~��@_~k7߅R�9V�~�;��Yݶj�ރ5g`���:6U�AmG��O�<�X�E?=<
	a��~���b���\��C?.���,6N���'˓�������������$!K.�:��v;���o�Gj�`6����$���<+Mc�lu�AA�1�9R��HS֦D"1�9�HA�7l?��͉��Cv���w�X�D巹S^���|�ߞB2t�&�rL]��%)����iuF��IP�I�
��|V��`�.�2Sɻ)�#SnB�!]��^���t"#(؏{�D�'T����g>���1���g!�T�"��S���زqz���vn8�����i	[b�Xn�'�peǐæېoƆc�-3ų�NɃ�SK�;��Sjv��E{d8K�N��i�́ ���>��b$�Xo��;}V�FϽ�eU�cx?m�R����4�o$������-��p�h7����L|�6�(��ׇo��E�����ԧ�~M �y���v}��t��,V��L8�~�c;6�)�|s�S	K��S~QȾ��a֏00��Y�a]��@n	�%=���xo���z>�
�'��q����;��+G���������~���p�cU�����������(jwrםH䖔�6e��~c��K1L���/=��D�/���篑7B����G䃶��)�+C��X��`�dvn����V��5')u�R�6zP�p]Z��?vT9��+�B�2��3���!:��H`%�2� N�rC����Y��Q��Jrs� ~q�\�ć���hn� �}YFD�Z��@\$e�V�!�5?� �q���Y:O��S%�~��.[��,�roW�r������P18B��
�M �y��qc������<��x�9U�*�Q̢��^%���]"���9��dM��E��e��瑱��f����Or�_zIV+��������AV&������>�7���lb�['�?X5va�x�����2D��'sI(�		�G�
�eiU8JN���D��к<H����C��� ��[AZ��q}�������[�M�9 XM=��x�'�>^�A(mj�B�l��,R]��؛e���LPbv��$���������=��e�e�Z)���R�k��&�����ę�x56[��@�\�P�b�׸�d�IP�o��S���cP�&��	����p�f�&}��8 �pBu�!z��Ȭm%��M��.n��V\C[�!����M0k����O��6A�%H��e��ًvIs�DV�C�;TC���3��2!��$�B8%�	�l|B��W�#H�"�6�QVl��k�!���
���=��",�_��������+�^�''�����;~>�l$���	�^dqF�X�i�f��6hZ�m�C�(�����A�7�1�� �
_(��꽣�3(�����I���Ȫ����A�Z��8ٶ-�2;T���� ��͈%�����w�ݣz!/��d[�
5�3?IL�WO(�26|��9˂���\��J ���0�|1�gY��g�CL��SRJ9����Xr�`�_Gis��Y��9K�?'�R$ PM� ���>��	e�!�j�`��^����-J��b#;�i^Ww�)o s	p옞62�@�{&��>�I��M�z�v��؏0q�2��n�R�'�4��T0�ظ> k{�5�/���t�ܪ��Vh�G-��_Z]*��+t$�`k��?G�(F���� i##�����9�$v��*U>����R�X�� �j+�����y6�/g��K��S9&��
t(#dG	�n���Qz��88/5@b(/�u�h*I	�nM��&����'ډ�p�KT<h�5�nq4�"|���mD�*[,��K=ڷ흤��mϦϣ�������w������\~�v%+�x�Dp���|���/�����78J��quZ?�A,$�5����'I�J}#М�P7��p��H�z�.E��{NW�c�|F����v�婵��JΧD�eC��W$��C����ץ�X��ѕ�7�c���9r%�+b!@)J��\P�:z�t�`5?�C�	�wgݛa�	10U=���y�F[�i��A�S9�C��S��c{�b��RUZ��w}��q������S�=�sOj�ヨ�ͤ�Y9�"�N�fў�_ӎ�4xT�O8�InO7Fn=7�*��c�4���,F�|nn&Ov(&.��Uk�[H�{HD�꘥u����<!����S�f~���j���v���f���ԡ��Q�05��夜w 	��X`ku���J�Gh1�a�B��}�=>�='h�GB�1�j�Kg�&Ϧ+NW�%b���}3}���݌K"����Yd���9>���+��|�z�NE��9�r+��C��������D��|	GB�����/�;�r�X��S�oz�����9������hA�?������-�9��#��4�ٓ(��4�C���n28`�&�
t�mC�G#�n�����ˎ�r��i�r�\NYjp�B:\��j����2�ۻZ���/�?o�U綥��s�.02�uj�ե)�m6�$j>~���H�����	UU�)Zr�ݮ�K��S��jo3����?=�/��ș��+�+����YؠD6��8�����rG�Hu��lv�iS����Z:�Z��nQ�+1����^�-/ڴ�H����|�8vaK/���.�m~p�_�\�O�[Y�}'d�Ѽ���>�?�A�����+�$�k�؄YC#�:��F�������F��aũ�M��
�]Z�	� 1���\�F��<y�-6����ߏ��7�:c �}��-:�\rR��UySܶ�#�EUz��g���=��C&��9I�`
"L�?Ʀ��ýE&�+���:
��NޡK�6����b��J#V�[OTyEN��.2#� r��a��"���7g��Ϸ����kXjW��d��p�DR�ܑ�Տ+�`�+�@52�� �QO����è��`NTт��S�Q�P���]���9V����?}T����(R(T~_R&�S��4�.{�=�'�c�㼰�����]v���²dF�w�^�p7����o���;�3�Z�ʌ�����*�C�~���%d櫍(ej�/\w���纰�>qi���ӂ�p�������t��٥���\8hq��F��^���\k��7&��76��[j��=���~Y��C��r��Ej$���~�B�;4X��I������P�ދ��GHf 
<A�Q;��B�_�n8]o1ǈB��P��u���P�d-w�C���6�㧁�O�1�Ts�;X�s-��q�-����ȡ]H�J��d�Kz�b��f��<�p/����H3�]��F�Ht�}�.�;0l�`���3?�jRv����N)/{?̵��	�]5��Sm��'L<d�� b�r#����6���>�܍xj��zi$���8�b)�0�qH�|��J	��	Q�
�4�#Y�А�g�{��%7;H6cH�M:?[Hg��*d�B��#{0�v�����@��U6��`A�����(��LƗ�� ���ߴ�

?��?u�����}eVyh���R0�4{��nX򓁌1�K/�?�E���5��O�w8厯��=[:(�C�	��x�����|���RN�l]d�s���'~S�����Ç�y&JO;
� �K��XGL�><����\2`R�Z?�'#����^l�S��q!X:����o
�7]���H��t��t��8 '�t�v������aT�A/�i��?�F\9+B�s?��:A{��L�Z�_a��QYP�F�v�M��V��W�"���T$V����4��w��ߞ�����)}���<��{z�?d�$.�w/�C�E�Kuu鐷U/�|�AǍ����d;��>��0�����^G��c��S��R�+%%�U�9���Tn�6����t��T~�^�����c)�Y��Y��p�:l�;$�l|nF�tD��<�Q<p���PE!yWG�m\<E�׳��7-�<�%�:��)�c�Y�'9�e�U��� �R�,��j3��Q�9������c�>C����zl��ء���>2�1��f0���+��Z�,\+�Ń��^ܣ���4�,�	�#9�JM�9��º��5�c#!�+k��1$�@k9��rL~�=j�T��C�����ꎿ��`��!����ot���0R;iU}j�r
�a4!�@��"ld�5�����������_,
5� b��/Z�;�j�Ó�~¡!xc��w����D�,�|��Q����m��##B�<�K�hX������QVs��o�C֠2q�5���m�#�W1L@6�W A��rs'�y��ԉj�p�"~U ��P�<�=�b lᶹ����G%:$�:i���<��>�߂����wpq$,`�{r�:���ad-'�?�2��S��yVB�ܒO$���J���=Ǹ�z��d^sa!k��I��|�����R̳;�kb��YO�^�y9^����Age��OyE�sM��FAQ#,��!H{�-����;��O��o50߫�}�n�f�R��4��Ep�/�?�����3#��-��6R�BV���ާ��Q�W7Qdք
a��`f��ށ'���׌�B�0����B�3��-�6'@��öT�����B��w��F�q�F�h>��縁{���!�K��(}��`X� 08�G�k�hn6�5i�H������e�P頝��C��K@G^T���!�ו$.)���!e6������c�Zi��JWz��"��(]޶x�dUƁ�{_iG�����Q��"wd�R� ����{k�ZJ��/6럔.]~w���¾�]He�9���GR�A�^��J���꾠T.�����,W��N������ʡ%��ҟ���J>�����<#�g�~O;g�Uৌ����W���_0��X;֑��OdP� ���q�@�#&z�c���4�vdص���������ըSS6膈���-��"Ȉ�	���������K��1�gi�e��<�{�hQ�T:�x��㢏��@U�(�kVl�K��]E�O"og	�yK��ן�tg��@?Ӧ�x �Je�����S��)�`��h���fU5�[�9x���J}���d��6-q�٤���&)yF���Q�2��/�׈;����e�'�j�Bh6|�.�	�K��ř�t(����`�V�WTWq�W�J9ݿ�>`�.L�i��w�����T�E*��w��3�c".4�����,?U���Sr�7���D[v�ea�+噯x-�;���IGlՒ���w��+Z�t��:��,,�	��(Nl��2�f�"q8�.����[�2�ߗ{�����1�m�!Gජ�� <j���KИ6�4P���>}�eIC�����|����xW��z_�+c}�U��ٮ���e�(���&�-��#h+�����&�2O�97�˧ea8��`�����P���s�G;�҅@1�^�|z�ֈ�q��oȳ �=^D7��� 1O�Ρ�����<Xt�����PYer��l�Q$*��~�@Iw�ҡL֚������!��m�`���|���Ҟ�>u&�*(��N��p]��;|��֢ʆ���7�0b��]�`�^�&BwN�!�4���c�[���zg����� )���fk��S�������k#I0�L��NI��+ӝ�U�"��w=>	�H]ɽbR	�J^S�(�Y$}]��N�yٓr|>�t�K��
|N��Hـ�o�;,�Mq��&s�m?��?��Q��L�?�t�цb1�@���g:��j��B�FT�W(	���Y�kT�U��UIL�F���몎<�E,�UB
�(���Jt�*�!�Ӽ�$C�/�8>�x�v� *��2h��4a�A���&���\��,k B�$�z�3X=�����0�+��Fh�É����P�$��Lk�$$�~��{p}���ȹ=AJ�����=v�I"!M *�`��#y|]�xB���z85I�@��l���N̽����x��E��*��޷2�\����k���1E���	��c�z�-�=�桲!����h>kyګ�a+�SPCp��W�v���ֿq]?����� �._�����z���6�Q�]��K�S��U�E�����q_w�NQT|�w������P�x�zz�V���<���R��ּ�9�Y>T��Xy�?׻\�DW:����<�
�kEd
(���6%�-���k+����a�K������a~q�A��dg\,՗I�Kܑi�1ֵ�V��0]�?5���M�3c(޽��;"��1�� O䇒X���F��a.�6�uu��P����a!?�w��d$����y��#���w%X%4B��\a�&��KUMIb\���>�\��Uy���1�QX@�8�T�.1�~���!tN��J�k����T����S%��-
C���Ԃ�j�PYf�F���\~�^��3FZx0�]�c�ݭ�b����}��4�w����߉S
{[�������m�S�T/��K�
�j�
���uQ}�0ϼ�&��`�^3��d�������f!�0�Ϲ,.pO.P�L(*⫥��'�B���e�����ޗ	�pu���r�'I���;��$=��.���Q��|�.��ӓ��?떣ƖESa���@�`-��NI���˦�Gl�$f�$o/��!����QL�%<�DO�t��$V�FAs����xOiN����Y#�;ǵȮ�|N�q�rٶbΣ�9,b֗�>���O��jp�Ň�����w�:D���0��_��bh�8�ө4W��,[Q � >U���ԥ���j��Ku��`�$��cL7���r`�Uˊ!�T�� H�֘U&t@�FH q��+�Ҹ��&�{MsYl��p/('�	eDs�'��O[�����F_�IA�t�.�X����G;8��~�Aa�7���HV򡬶I�C�'h� �������,�q$�L��2�&�"��u�y�@��\FͮAH�26���14���\ڵVj��cۂۉ(4}��g�W6��q� ��͋�(����T�#�le�!p^>ݝe��O0LAk��B��3�s�St��E}���:9��e� ��Yp��_��M�"�C)���"Н�Vݘ�ki�@�ɽ���?���ԫsH#<ï׿��r#��Ze���$S�2�$�i;���ʢ������'�\o�n({��`�	��d�u��ǟ�/���yo����Ҥ�p�!:�/H�a6e��eU���`^�4�?6�%7|G�]��XkIw��צ�����'�
�c��?�ƪ�x==t�Bɟ�3�ڠQv�י�i�.��0"�H_��}=X�iX'ra������"���kt�Dq%���Y	��S}y�]�?��8��x�z��py�������q��Lɡ� T֤!����<���Ň�׈=�+��x��D�
{�@yݠxV�`J&`�k-��6h�
��t������
����+R���D
�g�����a�+�w�Lnba�[�А�{���u�=)n���7����'ɴ@�a4�ı}��{��4']�-y�2���G�ʌ�+��!��	���"]a3�%�a���%��LoZի8x�[)	�}���F�)^Al�u'ʑ���A0��}�N3g?֌�c�O&�IW�=K��_����kI�j�V����͏"h?���.�/���hF��g#ܺ�y�dQ����'p��a�[4G��� �6d���H|�_�~��O�,M���X�'cb�A�T���h���PK�#��-']e+r)����������!�9��ڃ��ɝ��X���uw�{s��˸Yڔ��Z��!B�K�4�Y�-�vD���?1l��>��/R}��Ʌ�u�Z|z<��^�'�j��H(y���/f+��<�I�Fp��1�4Gp�q�}��	=F�A�j�"�^���*ʗIX�o�0�g�7������8���G��`�1(.�P&�L�B���l7]��Ӎֺ�s7��;���`�Sǫ�}E���l���Q�w�k0�S�=Hoy�A��	 )����O�M���st��\�50�*~.�?���'X+)]ko-�ݶZ���1_���JK�\��RL6�n�#4�-f�K~���x�Gc�FQ΋�ݟ���^�\���#�<�U�� 9B��T갻z鄙㌬Q˧���mV� *��#�1ԯX<N��D�F����V���b��m_o/�i�@#h4�/��&�&��9}����p�RFoW'��w��*�BڹI�t(>���4Y�4�����9QD��>X��5��aVa����ۺs���P�[��$��?�Tc���b�e��ߕ��],��o������V8��T�U�އ3?��#'�f<���G8�G$n�`X���Ֆ���J$�H�ZD�HCv���;a���ۯ���ˋ!�>�a�q.����� �9w�}�N�MO�y�z4<�r3i���M��]LD�|{�5�0sw��$"pS�0Z`9���&<��)n�+R�i@�ʻ{������S4���	H�����`��5"M`Sɟ�If��:�Gφ}���R�z�]��ՕL����o��	ŜxQ�&[�/7��?��H퐙�`�T���+6�JEfb�'$�j3��Xs�X�8�j�/��a���R��}z�?N�<�<<X��L!n��n�Ϳj!�bٯ�9Ĩ��j'5������.-/Tx�'��h���-F��':y�t��
�z����ъ��;�2�J��g%5wd�'9��3�����;D�jxq��b)��J�̯�G*�7�N)�U��IF�z!�
�����j�R5Zo*�
�L�E�ź�yX���F����l l�88\Ơh�u�HA�ڱ���H��W/�k'��F�arz��sV�H�4O�z����[��j����my~F����I�q����fm�CN��4��;76���J��sܰ0�}�K�y����o��������4Y��gT�<S^���0������m֗fZ������y8��n�m��#ՂY�C0�"bJJ
���N���j�l�n͠�;�@C=p�~<�=A8ڵ�,i��Ƞ����]b���X�`�a�L�g^C�ɣg�Ua�+����c��3�}I���ss���KfT;:q�y>�^(�8L�ř�QLj��,���~(�EM�n�x�x��;*�A��-�]�q���#�{A2�)�M��_���G�?,RdV�qҁ��q-��]w�;x��8�%�D>�$����!j����*cu��ѷB�� ��Ó4ęNo��"�OW{�ϱ�;e2�*���v�	'�.�]������A�8n;v� 
Jְ�y���=n�N�2MN(��ou��-A��ڥC�g�v)@Z�-�&�DA��N��r��d� 0��
G�1^^���rDMi	> �)��2�WMi�n8C���2�����`���A��yL���]
E���ΣU����G�p�>��j!���CI?����s1���+�
��B�1��2{��x��'-0���Q��0kx��t#����!����q�
^��֚l'�� ��v.���	�:�s��%Mb�Kd~;9���<�Y�힖F�F�W�����\e�Z\�\�{�z��y7����Gy��8��d�����3�����6Ф���l�?�յUg!]�o��o�}O?2awDf���)�N^�?(��J��9���Jr����S�z���HD���������Y�X��[�ݷ���GQp�������lY��9�QY����Q�,Dv�>TK+(�d~��M;���~\{���s�ٍn�y�W�%�a����t�.�.8�V"&gG�r����+m�=��݀pi�+lPx;�L{{�I5�	z�v���u��R���{�t��c��3�,����\�r�v���aNIg�� ��he���|�OQ�kD,��:I4Dv�
(��ݸ�mҮ�0���*�Dل(s�6]�0l���� �Z���u�+��0Iq_��9'������^�rw9�/�����cQ���T���z�%\���q��L�tM�h[B�,�qH���&��F:�wW>�_�̜ޮk�[���g'�;��AY!�	�,�^��,Sx�r�@f
R��M���8w(�i��1�!����E=b٢��-r9���ƭ歂Yd#���F��p{:J��8��Ǆl�'�qV���/�Di��׷��dJ M��f\4M^r��?�n�:�\*̳��6�L��U3[S3w� �������Z�#86#����L������$o?+IY����߸H��rF0	���h�O!�>~��@Y�k�f�^*_�@M���un7�M��++�v*�Ծоflu�� ��@6���*^A564=��b�O���M_��t\aIj\�[��ݚ)h�2B��n>u��,��Q6�[��v#���lɤ��߳��4Rj��d�/Ъ�H���[�8*D�����J�c���E������-�I��l`렍�F�'��;�m�Y����G3ʼCr3��2�r	;��}�9	�d���rԫ��� ĄmK\��:��+��Ƽ�<�l%��q2�+B�΅g�MB��.u��O�S�f\�)�:@�l!�)����D1u�&O1�p�n.�/���4�T�5����cׯX!G�%4��2�yO ��ur>�-Ej�؝����:��N�[ɽ8��">�^��s 7nó�w�9�I�� T�wJ��7�+k�-�8� ���>t:1���X�AG2�M6�gLq�蹙�2y�=�Og O���8���PY}IjzK�����B�c�խ�<˽<�[��5�ߏ�d��S^2���`Y����Q����l�Y�_�)=	m<�C��k����H���D��N�߳p��;)U��D��|���� ;�3���=Z ���G�.�x}�8�W�q�#�\4�C9Ka�x�75�lZ���䡭�B��#u�G��T`��qۍ�FL�I��w}����u�	R ltԎ�#�	݅���M���s�{a{�PP�H�Yo!6�G/��5�v�z�k�3��l���X�����ii���	���O�^=�>�KN@����Q�A�vRX}˖Н_ ��v���o������=��\�U�҆��S%���d�;$�M7��7!!s��_o�J뮣g's�:
�t�8�I1���^�=��#%�ՀV����q��.Ҋ���%�>�gX�"�vE��<�al����߱PQ�(.�z>�K�P��^(WtZ!�~g������=�B��@���݈o�x�G��ϋ�G�Q���i����<��� .Io;�U�`�
3�����'�_Ǡ�7�_A�Կw�;9��9o.WX�	�v������$��9Ƌ2J�D���|�R�tay9�3�����]�� ZϦ�rQ76qb����h�1b��>Y���4Q�'���8��~�o籽Y|��(�h&D�]��R	�y0u���'�a�|+���,Y�
-�+�V�C0��cˊ�1�:v@	$�=��}�#ŵP,�:�}i��EKt!�B���������'���6�E_4�!�k��}(�~�9�@8s<�ϩ2����ɪ
;x�lT��5���������O��y	�����@�˯�lu�+}I�|�%���e��� � ��Vq DCI�T����� +�.�%	Vm��|O+Y=��!��$�� �(���Z3�������!�++�i��W�j2b���f���#��S�Y�.Ɗ���XV`�|a[�2�,T�h�@��@�![��@���+/�9π�����K�����<���VG����SW���I��6�OU�3�8�~nLܴ;�������w�ћ�=~<G{�Mpj�V8�/A]m�U��������Ӛl�54�H�|���t�g�>���6���p+p7�q4�{b�v�n"R�0�&��y�n��J(w4�񟋱:f��ˀ������?�]$L4o�m��"��`H��R�My{l����	ͷ�)B���'@������,��������/��͊H�og��a{�f{�RFZqre���"���A;��!�6�aǋ)^�e9}�=�����L�k�B-띆��
Ft[9*���.*:ŗm� Q��=y>������v1�$E����I�|�%2J��l��������� V����W��	��ΰh���Af���#�7��K	�8���+�{�r[{�Z�P��Ψ��.�Jp�����D��SH�cꉋ�hs^@������0	���W��N�WM�1�%���Ǻг��Wu���/G��� S��Yfat�w�R���O�}m��'���Ԣ�"��b�[���^�9��睡�W6fJg:�=�"XM�	������8���w ���g�`�K3��.ؼ4yZbF"�b��ZH�Lk
#�I��M<�S�̋���f��G��5(�;�q��=߂����Ͱ�02I=�x��ut@@������/:���C�	�YP�+"������،Ƀq�8%�5�p��8�E>���}H����67}���pI2� �U�0��'!8�� �_�2T�{�9��"'��<�8/�Ռ6ZUGr5~�LO	+��O��j�7��g�ly�rkt�g�@��v\�M��tCEI�dE�ɟ����;3dΜ����T9�U�?9��ɶHI�Z���?�m�w�mA;��*���P5W�M��M:	�|*l�,Wۇ)��돇�'���^ك��^�|���?u�!��	��ů��=��0m�
�p=8�����5(�(�NI<��ɛ�;�D�h�Mg��m���u��t����&�����^N���)�?��,{�s���.�sR��7�����}FC7�v=ϭ�	3��Md���=�
��Md������xc�%Km�1g:d�.i�|��ЩX����,�o���j��a��iA��C3mQ0�����]<�(��6 ��b}����,/�1Ku�,)=�g�I]�U;�V`A$}TXǍ?����|���HR�+<�K0���fRYמXa�L&Is�z�3��Er	գT@�7I���NlX"R1��5��XF���܏���|-牙\���%o=A/������H�K�i �N4��
�@W�x$��`�ᔽ��77�J(�l��9�xK���<cpȢ����l�S^T��z�k��n�a��M_2�y��b@/�P���8��:��I$�!�q��L�8 S)�1~��)���*��T��n����w�Id��ʻ�����;O����l� � D%OE����CL��l��$����8�h��0Y����l[�i"o{Hr�e;׌��pW�&�Cn���։-rp�:�(S��~�yC���l������m�NX���eq-)N�NI)2JFN��w���;_�0=nO�X�?@�%8%-(�=P��������yD(N���Z��I�^V�M@�3N�0��Zѷ��X�3w��$(�2ء: m����R<fO����Nd�c�V�{69����J�i`Gc��A�.Dp��vrwV-�w9�D�N�1����F�q*w����J
�e[xea|n���,���J�!���x%x���-�1s\�y���T��Nz�A"|���d���+#§Oa��c~�V��H]�!�����w��;p9�L�c��2���5]��2e��׹���z��2�w��I1�̊�A�����ċ�X(���x2���/��9׆ՠ�����p�P#�w��y��u�K��q*=/����y/�^M�_�&'?Y,�f��ro�������tmQ�Q?�Տ�º�G	� ��Z�5�
�
�c��������w��|�p]h;N�j.Wr�`:\za4�"�O�Y���6(C���;�i*�Y���?j?�2Iv�m2�˄�5��{�2{X�ѱ�Q��9����e��L�*1�0�y���ޤl,����/���#��|V�&V�2׍l�KS����~�n@��w�LvE� ��|p�#���.ԩ߸�V�N���+E�ΡmRlLl5�vB��f�_O�U��c�.�ID�#Qa��vH�[E!�{���@zK����%?`[�[�铥�)��rML��,�"��6i0z�7��v/�L+�{h�40{�A�W�콀8�c����P8�"�c}Kt��=5%��+�Fm��r^��Sq��+ݓX����c�U�i�v3���+ֶt����������0���T����Ϸ`��� ��(0�d���F
D���u�6����,��Ta�`��9[H�.�jQV����8!)����;�v�тf\
*�ܜ��a�"�P��97�P����Hx��w[Pm+�ç���0�(b_���ER��ZdϪ5Q�퀝3��Y���>XV�w�ۅ�܂ �J�߇�Q�U�b	;W�]��:��Ҧ�!��~��e-��-�5�k���S�'�.Fbf��pd��I�n��O�:1<\^F��m26�ԟ ��˄�����M�TC�I�i<���d��	sy�sk�Q �e�^�ě�-do�;N3Aƭ�������AϹ���}8��W�X��'$�Ţ�ˆ�Y��P����1����S�8��nM!��ȥ��%���b�X��fp�l��+T~�^�����`zMC(6a���'T��2i�]�5K�������s䪸z@ P�
|s#���g�� ���)�s]cO(�ʛ$��l������=��U��Q3�?�ɑ��j�����!I���&����t����� .������j�8�������P�*��\%�Z����~'vO��5T�6!�Tg��3	m�\���6�H��=�r�U(w�8��ܜc�7�!`�mG�����#��g�m�:}���Ѧ�Qzu���sr�1�Kv���ϼ�#S�z���5M���C��V�-�d���F%���z�hg�����ol{͐9�s�s��Ƀ�{�H������(gz���b�B�U��&4�ѓs{3��¤�7���g]O��]w(�75��L�������Ҕ, �|�95W�v������}�B� zNϜ�Z)/��*e~���çJ!'��zQ)�n;��v衷s2�x�k0#�)!�=�=�r�"�G(���㻫����I��<��ڰ>x�WՖ��s%������dmQ�ٹư��a�]UZ�K[敝���I.�߼}S���|���ը宨����B##Ou��|��x���Ź�v� ��g���i�(+m�O#%���J�w:��.�����n؏��G1�`h��LcBA�q��u��/�`������4��f)@�:����)�JBO��hY�9���0�u��a��0�e�G��R�1�KB�\���d�U�|�U!���l�+��&&gMF�2�����׫vR*���U�䳽_���qY���%�4��!���m�)����EU#�!暿qbO s���0ro�q8ƻU��@��O�..��*,��{e'�8n`s������^-��[L]s~��&�9N��0�_�h���&���,tgFqyơ�=���c�SC��}�}��ˠ7p��$�߲ٴ W�|�	��c� ��]�Q[��)~�V�˛��f�3ot�	R�ݝSi�.%VmhOX�Nb����̔��[�Y���ӓ���{W/\~�Gj��#���If2�N�1B _L�`��?6�N�Q�N��[��9� '�����u0ٱ((�"k}�����Oz��.��t��2e7��;M��;�K��	O����]�g@��2���])�-�7mMr���*K�+�~���8�Xɤ7��y�|���N�EK��?O�q��MiQ= �]�A���Έ��ۺ]��H�,dѮ��mCh������o����Z�.Ñ�v�Q��N�,όvԅ�Y�h�@���*�&Ȧ͛���-*��d�o��S+����l�s6�0'#2(����G"$����7I⤔�[��qBȀ�w	e}���n��+�/tO�)u;���d�z_&'��FR��f��|��/���O,�b�=�(�
�/��}��*�e�����f,	W3��}�A1���;7�7�q�z�@���� �왡�tDTؽB�].2f7=*v{�@���D����ے�������]�wh$�]4>(�yw�C��'�����sS��>}��'�n�Mn	|*���#r�
�G�j��G.�u؆��U�O�9���X`�>x�x�f��W.�	�nYI<v����:/���́!>Cy�aݙb���
Ձ�;����Pᤣ5��bn�m��R�&g/N����)ʇQ��K�9*e܁����t�Y|7�ȣ��h߇��2T�D�t���C�JÂq�#@�*?R�N����;^���<69	����{+R+�1Q��g���j�Bx>�A<>W������k�Fkۧo��-@�#�p��x�������_�B%k!�}��]��:�	���`�d��1(|c��@�>�k�S�X��an��=��$V���
5���9�e<^��r��hC�.o�5
$����7[z��l�G9�im�?�2b)Blu��N��ѭl����vڎq=8�4�q�`�ˠ�H�#o�qy��*���\�Y$4��%�]��� m��ҕ� /�_;5��U�!OJO�~�%���G��@`�"|�n���9)��f�U��'*vU�荁HSJ���Zy�7��z���tU�����
^ȗ#W'm ��f���<�e���Rt�z�Rj��)�uW�7����f1�|lx���6y�MT�	�֨��)MH�+rFOB�%:9
Զ�g���E=����w��LN�*�x1)=r����7mgY�tr�(�|��ttLb�u8��\u���$�	�������Z�I������2��}�:�{�\����Y#Lܧ��"Ό�:8�m�a,�y�^��>�;�.�d�Q���X�wk<��@�5�:�zl����b�����r�r���r��L_��Nt8��Έ��Y�������ךּ�,�7���>f��g�kĘ�Mw�������d���NƉ�,a�f�+� ��y�k����ł��8^gW���m�C��_�M=�,	���Gܷ��zw�2�{�u|�2GVǡ��7�����.6��\�dn��X17kZD��I`��z�%J�{-B(���?1��k��������\X���q����IF������x`�ґ��V)�'��R0F`�����cl�{l��S�)��%���ְ<�E.{�j{OBE�ͦ�f	�m���}9����gƉ�v>]�ePBQ\��u�$�'?,Bt�"������!�8m6RԑĦ�"z�������%�$x�C�:+�RAT�0�5~8�ߌ��|\��� ��:��|te�GL��X�ls �K��Y����e��������c�	݆N �V���<�f��Fa�`S6{a��Wð��a%)����'G��<!z5AeV���g��%�2�W��ف�ͳ)�tf#A/��n�n�3�a5cTl��Z��*�xT�wr	��s<�DV�n3EheY^,��ڬ��$�S��Zo����d�����-|��_U-}�F՞����`�}��x`����e$]��G]�꩗�}�S����?��V��Ed.����-���E��q���3���_F_�=�{�'������IM�5���T���ab鎶����zG�h��f)Z�U���wAO�eF�O���ɚ�-ak=���Nz�^Vz��Fq�P؇o��	:Y�X�7)���E���5pp��&S50ըQ]dY�ׄaR��k��x-Ȗ��P�%��.�K�|~�ۺ~Fq���}Z�eI��H�2��o�o�5�L�(�h�X�c�OW��B�7�VxQ�k2^�~��bӤNtm$�o�����3�;��$�?$𵕶;���%�u5���+��ӧ4������paiHb�$�ּ3D��i,l�b�G��ܝ��G��ek���S�����'u�ݿ��J��g�O��Z �@�

,�{�F�B���eջ�QѪN��g3�,�РQ��5�RP�9[�yѺ��6��`S�1�&{�1��᚜��ى����t&`_�Ld���r�#��-^شoΈ�m��c;&d�X�D���]BgAC)���v6Of�b1�;�u�]�n\V9�_�۽���;��iוa�T*������`=L�T�dq�ii�����J��Bt�c�l#�, �U��I���Gmk´��BY���gIq�����F����tȰy2.�����ʁc���k����u<ݱ��Лk&uZK^���٪��&�K=<M�L܏ŭK9aJLWI臀�/FT��L�Y��|��Eˏv�Qs��p`0� ���(��L��t�6�yLN%t g�)�V5�N(�.�j�ܰC�/����ǰUUnխ�����.}F�ф��*�e*b'^�L�V|�����7��1��Vg�q֣W�a�p�D���	�Yd��9��uȕ'�o��+���M��o(+�<b0cl�Z1��;Y:�[0p4�T�X�3�|m��C�î*9B�S����4�a	�C��խ�4dAX��*oG�A~nĊ���À�+i�^�_��ţ� d�B���N�q�w�tL�lT"���Q���~R�h@�LF�aU9p�	4e�!�hTIN��n���k�����"��Ք��}�����7�+�LMW�3/���݅Q��C-�(�mDڬ�	����/��8@ε����v�u"x#�_>�0��YR��R��LBx�y�wVo�	G�k?Aty`���II^�p���߾�Eq����1x`m��M4�X�f#
�o;��g� �������Ϊ�S�K���)���l���q\s7"��e��G"�F&��̓b(�Z�;=w���k��!�^w�,K"dF��r��3�#ؘHziT���V;ͺ��e�/��W���k� ,���C=�����}<h�v�Ec����[�ި�t���������QTd�W�Z�ү�(֝K9���@�=}��,��vKa���R�4:����Y�]���\�������g���	�PcZ���;یRz?�?�(����
��(@P��٥P�g{��]"-;��
S�ٺ��ǞJ�6���B��~����[g�W�4)D֎�2��g�SH����	�(�����ȁ=0�s��ئ�����~�K�If_���٣�>���V�(�J���/J�f�T��3:qUX��Ԯ���L��1��?�M���T��i�Cl�P���3�r0��h�%#
���E�$ȕ���g�ب�z�b����祣�썍kW����<��IJ5�������/�Ũ�jgS]���@m�������{�1���S=�}R��wB"��!yEVB��Z�wjBKv��:dZ��������4{��3��;�?Q��!Z⧠z��N<S�v�S�%���{v���)86@�����#������-c��"ܑ��ѝ��`;ke(8�S����h���o�:�%�v���ƚz�.��=�v��}d>��Yv2_������&5��O�M��������j`�DY'�(S_�8RT�����.�e�
AV�U�A@�'�F^�q�Ҩ|�&�'��j��0+	�R�&������X���@�6fA��J@jP�w�V��@e�x�����3�:���u�����rT��8�� �a�grh�VIW�>"����7L�����s�?��%$C���	Z�o]^[�a�!�a#U�E)�;����ZAвo�-'�z&J7�5M�*X?�y�{?S�Ab�=U��Yy�7��4�	z�VULH>����L�"�`^��8���**#[�n���67��u�,����c�0 �'X  ����;]XaS��3�im\�{�R�C�.�&�wx��M�Dp;omV�6�p���F.D��Vg��Вk襶�:�5T�H����6�����L�o "����'0S�lK�y��RZ���
V�s����@R%��h����w?3�Uu1��$���	�`���\i����r
<��Y�"���[�o��~�$om�'�i��OgStr�"��Tr����>�tM���<�#��WɹϷ�Ȧ�C�9q��t�2n�-b+��������8��Z��������v�z�A�gi��uzu�P�b����e�9!/)�hkRҠ�����N�|�.�r�dL��۱F�+��G�/�2m�� è��V]�EN�e�y�;�ئ>f�]�j8�&9�L���%!>���ã�\|y���P��o��øN�@���v�h���)��=��������F��dy�)!�p����W������^4��
�-�y5<#���qU��N�E������h��C�������<5�/���+6Rn�%��88���`T�����`3��.�A[i��F&+�?cN�f��C���4P#��]�:Q���-�2�V�=X3��L�zf�|@o��Pz���!��۝Ei�׶g������c`p	I��1J�I�Nc\d<x&�>�^f�E,�9_S�D���'`��P:#^��z�ys�T���������ٖ%e���皗Gwӎ�PE~�V��C����=&�O��e�ℾ���,y�|�;�������ՠ�������6\�|x��	EMh��.g�dJj�t�N�_���:P#�vj K����Q�
�П�<�4A�W#��fI��2�Z7���w�)8�í��Q��W�Q�j&�X+@[Q��!<t>���v���ܡ����u��⟂	�&{?~\�3����Z ���������jq�K�ꊜ�6D͸#0�Fj���&~r�K�ck�u�s��d��Y�'�#J���qH�
�l{���i��a9i-܎'Z'��P?�oL�wN�i�&{��&����_�%�XV��k9�����yf�!��*w�����=�`���]���n���O%�`jR]NR�ǃ�V����t��;'��96��g�� vn��ukS���6�a/��W������@$�羁r�JJ���!~���)���oգPTnl��/$"�f�A�Mn�!�p6������!:��-+�I3�����0#��u�q}�<`����\V�� ��j�^6Zo���<ݽ?lc��Xު7�@E���o�R�_#���r�������k։+��U��'��4�����C�p��4�'��:�2-`��äPeL�#Q�39����A����fQ��d0�OOf�2i�����
G9���D~�q�2g^�-�N��$�ߡ�m�]{��A�ĺ<�_<������f>�#C4��*PGT��}tG��!���L��	4�܁��s���drt+"`b���=��wCty���4+0���u0ՙF�	3^�:�e����,r�=]��Ά� /���A�쁩����c[��Tb��2�n8(y�~���#��K�ڳ$Ya�҅�A)�¤�pT�jJ~`���9�����ڣ���ƶ256F�/{'\M��z�*��Q~`,�}���&��If��~w#������s�O�4ƺӰ�9q�����.M5��zD�Z��.f��G�6�H���uɴOI��,�J�;�YIe~!q�{�榚ʗ���7�(7��U�i{#�^{O��U�R�~��Cq�A�BѼ����4U_rʄk�U0u�$,w-d�D��f�`�x�-��R��cVg��W�4՜�����=E!��,)�<�+�_��%c�{���^0�q
Bg�پ^/�9W�JG%�G2�jo�gtz;�'Wa�p�]������5�@ ͥ��	������{��}1(,�K`6w�8p��6E��ϾyW��ew0��NVɦk����#�:��0xoL��9�YU%FQ�+���d��Mb�2�9{qB�����~ǮP�7�����Z:�|\��&�+\0���;�AЀ�ȱ�;'�G ��|�%�����QGw_�޳�eɢ/� `�-�몁�l�D�	=�-�|��Z=>�?̮��2}���F�E����+'4op~v^B��=�|����d����a�)�N��&�v���ј��/����ίa�7��9��cJ��7�����o�&Ne�����n\6���aZ+�
� M��[��K8;��~����{]����h)˰
-��J�}f����e�+��#���S:'lO쇿�*,6|J�m���<���ͳ��e~3��*IF��>��711#�{N7�� �\��%��պn{�\��7|��&S�o��빴w
+j�t�qtS�#���k
�da��ŵK#�T�R�DF���T=o�˜L��b�C�L[�gG����!�����s�i.�$C��!��=]���G����?;gG�~J[V"��0^0���d�0�iK�ׅ��ߕ��	��"+�`�o������\v�H0�ѫ����s%�+T��~�0��`����	�B�{�+2h�^~��J4������S���g��ٕ������ٿ=����*k�y�O�c�����(bR�Ѱ�W�I��K��f�1@�"2,�iA0����mz߿�i���ő ��0D��AI���]$P�5��D��7�i�ۖ7�= �Y2�Â�\Z�Q�t��R־�x4��Z�O�܀�R�Em��Et���l��\d$�t�R� ��>wW��#R~�57�l��a:@�C�"�LA��)`�wKaQ�ȶ3�:w�v��}f��2�w=ⱴ�A�{��`~I3�\wC�ל��ϗD�������ZA��R#�눞u��-�V�N��If
�	����l�����V���!�}
�(4���$6Ш�j�$D Ї�Yg~�v�r��i�W�g���͡�ݏa�A���Zi6��L�2�a�N!���u��������v8�H�B�&ނih �qπC�FL��˓Im6�s���������?w/��ai|��nL�q���������i+d�l�W%.�\�i�Ef�S����l{���h��+����&�P��׿Js-���&H��jfZ�m�;ՄV�]�a��CP�z2P:���~�h����2��Cт��y ��t&�o��H9�G�#��4���Ѳ�jO���f��B�y~ܒ$�7+�S:����τl��/=��T��7�Nf����k����/�?�e
"�Gj%�=���Q
�� ��v�+�^���B�@��������c}h\�ÿB�4?yt��E�n�o�='��7�Kr���!�[���x����W��mw$�1���B��5��b`&nD*aUC��v��C�ڟ͵Q0�x�g]��n�O�m�->��|`�j=�١ү�h-Dl�
���_����%D>������q�e[(��.�#�K��4��k�����2	�R�e$Er0��`��kV�x5���6b[�}�2ĂO8r��CBHſ2�/� ���ۓ\�0�
�ja�����˯�>���5Yu�*��[��q�k*:�p�w�����S�"/D� ��l��IOٙ
�UP��^�`�J�����:ˮ2R9����<y"/�����x�,��|!q(I�w6��yQJY�ƕl��"
o�(\#P�o����!Z��ۭ�}=:قH l\M��]v ���˵�m��>��z)���*VI��=)���N/(g,E�h���ǧ���;�h�D�k�3g��]�5n����2�eݺ��&�µ��&�����Oyο�7�X ]҇24���Z��?��~�0-�jsv��3)�NPH��&��#�!j:��W=���X�^x͌o�M��.���6P'2�T�ȼlQ
�цJ�{��w3)ƻaQ��'>�>l���Xw�w%��Bi�����.H"k�#e��Cc������������C,.���b���ࣚ�(I�M}A�����+���v��jVp��x�g���d<vc}��=Q��_pĿ�R&ll��4�#�n㱜��ɪ��IE�y��������f9�C,2�*�*!�(�����g]�E
E�tZ�ޮ�w0�'�T?�W�/(�.���y���KrE�,#�j<|�8��:k�-�<ss��U�l�{5��	y�9/sUt�C'G�פѣ�n(����P@'>��5��:=q,>w5��_�����w���:r-pA�^X�1j���_:D�eAh�u��~�E�FXg;�}ue%y���k}����/�<�h
�~�_Z&ƐwYw_�G#`�o�q�?��������\sR���S�.����=��$�<�r��-I9�-�d2�����`>O�"ē�H���xTeh�yHy�2�cY߱����_5�*�惟��TUm��P�Q��D#�{Gy�9��L@�^d6������ޚk6f��J�lK�%f���qʽ&ɬɽ���.|��"C���
��7Ǯ�n	u���L�v���ݳ�\ޢ�@�׌|:�ŷ�{ l���M��\B�ӷЇ�U�A���;,�,_��������gF?�������Ʃ���fw5/��|h��W���2z���@�΅_�Ofl��&l��?0έ���,%Ts��n)	07Xݚ�9�B%^@�u���."�/Si1���/�O��02�9����K����ӵ����Ag��.ch���6bqJ32���b����9�"h��z���1*��ؒ|�O��*.(�V�
�x��P�To� ���?�6[�`tÇ�F�j�IFtGA�*`���<��{���iL�����n�&�*E��f5�0��W8R�(�����v�1��~� ��"�|c�/�}͒B�E���Sb\��������e�"Ռ��֓ł<ftJ�U�v�8'�L���}�����.�t�p�Y�W��� #@C=�V��'��p6�_�y]4�0VH�
��|��x�dw"���V�=�̵/.፹�F����H�^��)$�89�n�-{��! |@7y�c �	�����ȯQl(v�
������D_Q���Y�ޠ7i?W����#�K1˛i�n����ݛ5�Z2-F�"��J��`}2-��ؒy�(?>i��C�C30��&��;Ý�%��bXw��Ud>��S��A���iC�6�Cݫ�#ɮ���2���~|>t���-��C6��(	^u��������Y�J���� ������`����jQF.��*�Lm���O�b�>��|�/�b��6�B��9c��MW���T��徳��tL�u��O�7%���c2f���~`����&*a��������"�ņ~l�ǯ�Kj̩�t�Eן:���{�K�vh��ކ�r�xJ�&p�s��x�\A��?2��A��Z�+ �PW�)�o��b�'�",Dw��@U���p����8�tP@L2Sʋ�#�j��04�%�+{$P�v��;a��/���C��>�#�ܠ;CG�=��
��xؤ-�q�(��~�\_UR���-��p��g������j���W����V,tDUٸ��i=Y?�W��T�B���)��(,���7s�9�����&G�������ML
����įqq��2q�v��6�*�HpjJ���賰�P]���XE�<��/0+��˴�j����	�܅�
��+{E��3���J�h�����Jy������";N�*��0i��Z1P�\W�;f���z��5�;��t�>�jQ��zgż�]�G��.�|�Sd�ѓ��+�w��L?ٿ��8�ѫ<�:]��5� w�b�e�}qD�PB>D1�XJ�NM�|�x�^:��J�
H��鳛f�nu_�_��cͭ�)�J��vg��%�=���=������m�<����߾87��C85����̣z<�P"=(�P���-D;:�g�K�;�O�M�Z;X��� �iT|��<��䭐����D�!(T�?��f6Vzx}�mȖC|6T����(��6CW�� �j\|p���frQ��S�ͣ�Tibg":ƿ]��EmC}�ǳ����7ۛ�~�!<��8�`m_��xC�b��J+._�M�!H��=wUx��ޝ�{}N"oaz�	�伜���t�YZ�۞ƶk� ����~��/�}�B����@��T;���4;���s�����Lr��a��Q�u�]`�8g��C��� �wh<o�9 
	��B�����`� W���"q|F�TV����x��6�I��|n��;8QƔ���j|D�L�kP��"�wb>l������ufŖ�&ڐP[�f�7�a�f3�rIµ~�[���Qj��٘y��wR5_�P�:�.\����A�I1�M|���Y�N���'�D��kb�)z��Y,�7�t�:+X����,�Rߙ�m�k�n�5�x7F�tr�6�Y�/'� "[\Ր�͚����T( �Z� z+W���,����[��a���V���5��,�
�����X�(:OF�E6�ų���!O4�� YUڑ�Q�s������yc��>j]���4������KZՇ�¤�wI��#��ʅ��nx>��00.^!��}�0o�&��,ӿ`N�ޞ焫����X�Ʈ3�A��a6v^�ZVǴ�,n�/9����3�~�c@�T")bc�bG�T
�
�u߳�/7�M�ۨ��R�I�E�&�=g�WL�-�$F5H��x�����=Ylc�*l����Dh�X�c��@�x0�'��x]����ͷr�qj
�l̹#(|�^�� �2���k�Ƌ���l��*��P�rd�?��w�����ڤ�@Ƃj���<����<$��H�d�|�����z���� ]�rSȩ�v��F���"�N�����@���Έ����yu��wO�^"3���T��aE����2#şNd?��֭��g��UH;>\��M�6p�ۺ����ՀI!��M�� Z5��U	F)�O)�H�0������ �JlVh��оv5"N���)v��|^GUE����X7m��7�����ynu�b���^u ����Ș�ly����SɎ������gȤC�ⓔ��UtqS6H�_� e-qWF�a�W~�!��AZ�^PCv�Su5Oc3����q!c�c����9X�:ǂ]�Zݭ���Ymw���1By�~�������w�+!T��-�[�g^Jl�Bܕ�e񎕫�����y�́D�޴_+�)�Z.I�=.�!p� ��,ثw&_(��k4*��(f�qY@�tke�+	��ꖀǀǢ����+#nT̞y�-t��yV��U��X�5��5V���;�F��&�����G<%����ˬ�w��cē�rRY�Z�0�lɨ*'����"]���Sӝ�A2([c�( :����hz�Il��whg[|����TNͷ�e�1
�\�@�����r�RM�b�t���|��Vfi�k��6K�kLRt��]s(�9b���g(�ґ��	�SmO�O!¡��.��A���6���X���=�)Q^LO�{�)��&�y����L?gN0/5N%ϯd>�;�3��D�>m�8�!�2شg+Ò��	�:�֙�&����JNL�I�Q��׵�T_x���ښ˚�̌ǵԷ�������S�T糘��Z����oeE�@��2�&9��(�2���s�F����v�������,X��T������gI=A�d�d�k��@�!=ճ�b32���k6"^Y����df�ĐF�C�M#��9#E��%�b��>�lG&)���XQ��z��Lrc�R��v�=>�5T���%(��DF�l��� �+�umd��jt�M�}СQmo�����O��uD'����T�,�
��S��퉑�>�6Q���i�=J"�(v���T��.��b"��.��`�{D]Vi_l��V���������^�%ڡ�C�H�~�0jFϞ���ړyO!Q	B�L_���̈cv;�rZ���w^�l�Umf�X��!Ek����T����NX�#g>�"^غV<�H2z�����Y�M�c���������L�m�t�ռ�:psu )t�L���'1��y�ަ!Ju����'6�,]��[����c(�,�P4��<��0�`���ǂ)��?��	�8<; Gl��+,x��zt����`	�qI4�C�)Һ��_A�
��Q2�/�ў�����~��
���Q@v������܊�S!Yl/�F�a(�0�1��Q��o�,�D�u�p�9�P�=�=�Q">�?�:��߂<P;�s�ܧ�u�lug���,�͹���V����	�^0rm��������q�](y��3�VLKKN�{�����
��!�*?S�VS`iy�&���b��#�e����-S�}�����������0��}����F�-�=E�����p�I�8����r�=3s���gf[�m}$������9ؼ�Q4.),�Ԡ�Vq��E�K�]���ƻߎ��r����pں��0$����r��p����C�d��Pe5#_m��Y�����1@)�c}��{xq�o�".��y\�k��Q�6V9�T�EP����^���x�wΡ�yk�7�b��m��ݎ�r��*#��>�J�1���Zx環����`�\�_�����M��,i�B�ů����5��V�V�B|�yo�92ʷ�8�{ ��Xo ;��<SS eN�Q� ǡ6%v��K�n��Ƽ'")<��Y	�f�k��iKB]��;�JIX����� �]p�>pf��/jl���	�+Y�+���dX����#z��<k�Y	��s�
�b��<���6n³	q�xF�y"i!�;�C���diE��݉tVh	��V;�mv?��@��)_��g_�������Yc����s	}�=U �J� ɵ^��*	�bp
���]�s���^�*�x��o:�zUYF��j{G�o���1
S�Gi����wr��'K�%\�I�E��u?��d�F�a	N��bL�'I��v	)%�C�z����c�5�\� -�:4�0�߁��oY{��4pZ%8�a�@U�Y�j�P�rML۾�-PpL=o�����2v	yh0�];mr�TP�(�:d4�z�9kX�#ނ�Cy��;���u�䉁/�!<e���k�\&�1�n�?�+���L8���T�Y�+8�r���{�菙����43�,V^Y[)!/=�{��o��A� ���ՃF�(q�+�f���J�lR�P�Z��&�ߞջ�$��Z��ׅ;i�I�&����%�R8�
��ҁ����R��.���\�4U�My������yS9{ԛ���!��t��j��d+�C#}S;�²��jFʺ@;�N�����M��,�����e�<���*����$r��}�@������#տ�\a�0c��}FM	=o�M�Pл��noe0�)z��Y9iP���0)3B�4��	U^�-#Z�h�6�l�k4(bK7Z��C�Pw��h��R;p�=�⯗40�U�!�y"�ws���i�F
��Ae4E.q�W6s�ZuA����th}[��8!Ho�"�#��~�4��J��U��(����ܫE�5��zb����QX;��=^�&���9N�N�����NO)���'k�CY� 3i�"���Ɯc:w9x�5P{ִ��d�s~\I�	k���G{�z��QD)�H����Y�%6�o��:5�2�a%O'9u�c`�1%���oUt'-�$��R��u�E � "�\)�a�	�O�Y���^��ȵA@�n�q�tD�#� P2'-b�{���������jFk~K��/܍�?�J���D9s�q�)~df�ΪT��k�Z"��U��C�P�鈷�|�3<{p�r�4;�����pS$��7 �kT�8,c�ݫ�|�*��RIHWQ�C�"��T���~�}�!�'��f��r+�f�Q�8&;�1�ӉEY��M���˟O���t`߷�V&2�H*�	m�o�h��7|eJW�!�O����Z�J��f���B�hO�^t�m���Q����a$a��C��޳�؊C��Vi���u��L���R�q���C���jJ"'&��t������Z��[0@&�逰��MQ�����+4�/�#�
P�qJx %�����
,���fP�* .�<�u\H��B�RH ��"���+0Y��b�T�c���aB���As0��j�� 3��������,#��Y߃)���)[���d�]����PY���5����kkԧex�c-D��׾���T������D�����^"�3b��� RWE�aQ���-�ٞ37�bG��}x�(�wK�=>�`'l� 3��M�ts~�:�X���	���G��-}��D]y�?����^�{�����H	��-@|���l�@�C߭�-Z=9u��%�Y
Aj� d��wK��ʴW��7��k!焲�(��9좽|���3p)#��ˇ��TB��2��7v���H���Ȣ��]F`
�Qp�=�*��
^3txR���0
a�
��/>L���n9V�Ҝ�%7h��C_��%A�]����(*�~�B�0�[WQ�`�P�'����	��B�K�_��S���(����Q�_��}g��]X�հ7�"b�/^�<�ikNG�ؘ5�h���Q��
�s���sea�~=�+O��)\ en
-��;7^}.g���se�]��si]·헜����@5��P'!�8��($�:�n*������d�=jHv�}��D
�ް�Na<�#7�sIe|\�.l.c�������# ��L��x�\g�Jv�P�V���?f�7:�/��#��o\-[ꀌ��i��4+�@I�fd���?x϶?��*���1.�1���蟸%/j�M?�~�sK�`�L�CL�0��?�𒈵�PT�hAWs9!nØ2�<ѳ�����%�2%~�#��輍�()�:��_�՝���3��� m.sS;����Z"!�&ѨbZ\�Q@��L�MO_�)]pX&?29]��
�5��(��ŧ�'3�G[��d����>]���>0��J?k�	&X����q;j��xʐ\-�!3�6�g�S���:Лz�F>�Y�*�n����7P,[_���;]�<1�h�xA%E����z�����2�on��nt��-Гe�"��5E�Xam*��C��<bF��94jo�A��uԤ�m�ց�1�&�;Л�P�������+)3b������5�/aQ5R�"�@����E(�;�>%�3��W��S���n�r�2���0�ʈ�uݿ�Sy�%�� ��(5�=z��W\F���1fJ�X�~W$d�h�l�ׁ���=Qx�����ۍ���p�FX��x_��{+�~��&_<����5�Nt�̅�~��g�y@>����V%O\R8��yx`�0�������*jw��A���g�5�Ď<�s+�J��nn�8_�+��^�N���8�nV𗌖R?�s���`��g��f��;���?6������0����:i�0i��ZiU[��Fbm��ZwQ	��.6A� j�� q�/?�]���﫼�D�11��b�9wr� ���V&^�u�:�8�\�#c��l�<0��$�=k��k��d[aG�W�D���s��k�D����ht�U��'�LץҦ�����U��d�7z������;���K(s	�	�td�b�K�C�����<q��J��vɓ�l���5q��]�� �M�U�޿|[����Z��lV榦�'P'��&`�$�i)�_�6 +�(m�6�݂"tT���/���Ӆ�� �M����P��������gB��Ʃh�a�4�>�#HLl��~bPK8�k�F�W����|:F#8KH�.�[�[Jr�1\)a�e|_�%A�w���7=װ��+Ч�y���H3θ����Ȥ11����^n��}Y�����&L�6<�|J���l�#�����,��}�*�$���fQ�&0�)� O��ƥ�,�������Z��)Pn�^�t�z�l�c�� ��ۜN�� �`6�J�+L֏���@/_�F��hF����ۆNܑ񽩨��P-}�H=t~Mڭr=�d�Â$��k��xfу�F�ͳ�/�(��D}@1�)�_��r<P��?��dڢ����Tu������#�v|%�g��ھ��c�M͕b!A��T�X��+�m���O5y�8��Ga�7�%T�!��z�Z�����>��ԄP�VI� �Qy~�Xγ"�Y}�*��+��~���a��ǥ��И�FZ?VI��;�{`�[ݜ�@�O��~ջ J�Q�>z3�����Q̆��z�k⛱��@���5���rf6��IØ<�� %U	|�$�*���VhJ�85��jF�,�����bV�w�ө������|��4�yO�*�?�g�����!"wчQ���E'S�� ��R$���5��2�)蠷�%�ŮJP��Oʅ��ꌀA���r�(���A\Pz�R�%;Ts<K�AϿ���BO{����1�j4�" �̊�1��֕���D���[��4�_#��1s���$�U�F�ɞb�ZH��X��V���n�-K��l����>	Q�k�W�/MdᏍט�3ͨ���҉"ώ|������/�,���Y�_�&����
]�4qV
�S�9[�1��p��"N�]�HU�@�c��VЎF��q�| Sj�23�D��*)s`TC4�~җ�� ;?F�x�nJd(^d����������� .�j]U��ۯӚ�=���C].�I՟�Ȝ<m�e-^xP[����Pm���`��˚LV��^�cZ+?C����+��X���xW`��ݹ�e�`,���m��c"o���@]i3&�s|��\�"��mu�_9 �ST���L�麿<�N��&	�fF���=G��P����%^���K�p:��jigl,�o���\�p����X�����e�xq�8��r���	�P��1��͚|��]l�a:�tp�*�*���R��|c`)�1_&z��K�����`�Yq)+T�q��n}@�m�z�f0z,�m��@��/�=�X;�A[�DEUF{�� jLC��u��"���W��+�+�A--y�u'�\̴��2t�$�7j�N�܎b�S�?0�YMy5nB�6 q�#�5�ڊ��hԁ�oH�N�,���;*љjp߭(¨���\|C����#$����T����U��z?d�Q��+tae��x��6:1%Y�t8[��B�ĺ�X�����-��r]ap�= �~����o����Z3���B�VZƏ`�� @�k���B	����B��kΏSB�M$��gf��8�"*����;��C �Yʐ"�En�Q7�KYH�h�:�� L%4ܛ���͔���
9U� �/�x�5i����л	A���@��Nο����OHW=�h���"�o��\�l�u��~�ѯ���*B�@���7�$�y��"C���n�������T�%@�vϗ
��Rb�2ׄ|�M����B�xTr.)�쒸E�,�}T{��]�=��}��L���Ad����FGB�gCE�l}$gI�ĩ�(����,�-�<��Қ7�K�f�b��p6���a%��`��Ĩs�	ۋEyU.���p�2��-%c�<g wp�y��]g(vF�7[���d�p-������I�A�G�T�p[ʜ�p��v�ו�Z��0���p��˹7�@�w`� JaO�?�TK)J�������~_�5�/��59�J�:e~�e��M��5�G�g�0IYsg���5+�)�� PT'�&nGXRH� g�{��(� �?f���@����w~U��I��M�u,֪aPq�7�^��V�8����\���D�@�`eC4���iPCQŠ���'����?�ᮣ��t�ox��d�8���_���"�\��ڿt2��]��(� ���}�5�h�s��PNT�~�����+�s5𘻗�Τ�m�uyEB�8��	��C�*xd�����7G?��ޯ�+Ba�6Y�[��'t+���ǥ,8�AG�K*�/o!j1����j�H.��p6�a<X�9v+,��f��9Ň�?�>^�ZC'���k�,s��4����W䁀��Ir&�t��"�`l���1F� �v�R������ך�JԡU���nPH��c�����r/x��=����@.&�t��c���r��hvz�'� 6��p:�s��x%r�0?C	m5KF���;Ք�1p��x��v^�����8��c!\�h��q:��W��򗻧����9�r�4�j㟉Z6Dz�k�Q��N�ӃН��	�ҋ�by1�(�1ЛҙS_�:/h"�(��f�SZ�j�	Z��t���3���z룞�y�D��Re�ny�F���x��m/���?��pgs31��HN�2�[����j������[�j?�������3�UL��9�܄��s�5��uqe�f��$�k���ٿo��)�JE���,�}�aM����Bk�	ҫm(ۉ`Wd���XT�/�_�LW�`��[���Y7i2��l�����jDta?��]�C�1��k�z�`���j�bP~��+�Iѹx�6�I`�<�n�ip�n����'�cw*p�Vfm:�t`��X��hK��_Ϛ��ӽﳴn���9E��C�����Q��R�.(w�r�&ZP�:sh��j����iK��Bh8(V8�PEz'�^�{K�i�G�u��Op��jV/:U���I5J$$1��Ƌ�T	�oN̫�g�E8��<��]�	�ŉ9�cFkT����C���8;���X��rT"w|�X�������ʐ��><S��vp��צF�|����\�\�X�Kp�-2h�H'�&��!���O]pǃ����q��%�Ų%�mh6��9lŮ Nr'o��f	4� N�ע{�;9`�i���]��>�0��D�����2�a7{t�����@:�투��D����qox߬E�jgo�n�3�������䔥'�gQ�T"���2x�}���v��]U�*����gǆ�4�
!�g2�2`�1h��OqW��ǳ��q�"��P�e��S�gʷ������^�L$$�U���h���m��1�M^Ke��\�xy�bI�(��[��
6��v8j ܷV@b:ڊd�L���ᷰ:j���v���+>"�J���h�g_>����@Sn�՝Yݚ[s�E�b�4K���.ٻn/J�}pB	��ڃ�LTg���1��R�iG�n:g%!o��Y����~���-��m�b%"*L�;�wXI����	��X�e��C���<?���3��)[�\x�υ�.G/��o��%h�w� �΢���n*d�Ν�
�
ŅcA~�7�Z�k�oG=���ٚ�5���Ap��`�$l��|O��[�nZ5��×����s3�^�$G e�\�Y]L�L�?J��l�����&Q�&��pz���>����?�F���7y.V��i9{��C���-ǌ(�t�?��J%@RkEj�>�L��W���h��E�t����'�|P"l�_|Wך���:�R�	�R�YTr���1W��J��:���Ajd-�U��s��NQx��l�"�<I�����_,mP�߶���k��lZ����]fڃ>+�!�}��w2$���>޾�O<Ȣ�3�a�9���%��E�-/��*M�����TuE(ʊ��l��c�r��n�$Ea�g��ݵ7`����Y@"���8�]�bd�>�H-<5Pl߉�ڎ�:��'���pH?Ăz.��b���*XH�1�CD��/�|_!��eSB7��S�����8�����$U�P��=��K�S�����.��=���������� KCU�&- ��R���(>%�7k��rp���I�߬r_D����ʓC)�.�#��ŗ�X��i��4�0>xPo�w;"{�Z�=8�"��n��$��{�"j7�5��6��$�uiĴ�Fi��^ݲ��(����n�^��n��yP�:~���B�:[ιa�w�_��o}�]f�Dp&��������RS���VɈ
�I���$3*J�&��ֱ�L�T��wҮ%���XU�9iO;�m��|��g!خ/�.5�56��R2:�f��m�#�݆�4&�C�Q7�Q��n��ջ� 	�Ou�e�a38H�]�S����/��z��s\Qˮ��b�
�,V&>��V�y
�C�(I�M^+��6a-�Ӎ�乯�o&䛃*�%p�L���1�Sy�2��j�R$,�)4X+���2��Ld3��r���?�	N�Sw������f.}�%��}�ݙ/��5u����L��oo�_x�:���Q���DK�Оg�Va>��������-:��7�����r�ﴶ���ŷ��wx�����a0��BO4�q����N�����E75�,�q1Ѫ���
`"I�+��jDa����@�N����l��mS�w�Ğ��F���f�L�S�B;��D)�q��]X�Q����;��L�U�+���=	=�UNI�׉��%,������6#�ѱ�U�#K�\wU���@R�W�nRJZ�h�Z�Cŗ��iZ����;B��H����z��k.>ߪ� ���R�E�I���Oo���dđ��E7���fY3�: 9�P8
���.� ����c��.���7���_七5���-ۿ�6?�S����n�e�i���^�è�OF��*���6bo��>)��)�+�$�A���9R��e���I���^	�!R�t�O=��&�o��<�\�e����0*� ���<���\��(�d�P�F�T��7f�@p�"�� %��6[V�J����M�Z��
��H��$��m�b�!����7��X��=����a��h-�p�dv�pQ���c��ۓ��S.Nɱ�5n�Y�բ`�.���Vx(1[�
����ru*̠�ؼ�<+HF��L����9;�xU���&�/�J��T3�&kv�F�T�hZ�.�@jyhf�s�lv"�PV.�#�T:L_�����	��&p@�,x���z��a�P}S%Xk>}�H8���2�;a$:s��5x�m�OV3CF�ny���{}I��xoz3M�cǪ��=�m�bs�t�p~z��9�My���>���� �|�7����2S0��T!*˴a7(�m",O���n�>�P(�`l�����H���X���N��2 j���q̣�k#���S^�b8��������~��#���YJ��v���dI�̪�j@�\���R��av�]@Rz�Շ$��L���ێ ��6u5�z��"gT*����k;�ІOtF'>��^�,�V�5R
��|��1�WfO��JƂ#_!��{.ޛ�w6�Nc�o��R�P��(8���R#Ə�,P��Ydǭ��>�7ҁ�~��$|��fg?��;k��Y�D:>HƄ��T(�d�c��c��/au�����?�9���������ĩpk
�S'�W������ra��˜V���œЖ�G����0 �<�OV�>y��	��b�T\{�-/�����ưw96��W�6��;�x�b?n�\%R*GS���"�_��o�y��{�-7���6q����9��t��m�6���9?�cw7�P��U�dWczh��}qU�0�K�T�)]�����Az��i�4$�nk	fZ��n�d��0�R �J���Q������u����+	_�.���^�JDУ>Ӌ6^��q�g�-�qt�TQKh��<��&|e�s�,���wx5N�aK/��lc����7�J�cͷV��Yrak�D9u��ˣ�R����@m��ng���6�-���>&�;T|H�Y���N���h�EM�/��Y:f�3$e�}������"*�~��x�m������猧��yM�_��Q'3(Z�q���u��0 y��q�#/�w�q�6딂�����%_�3�j�f�uk�NM�o�/�?sm�Y����UlDk!��`�ѹ��zP������ŶKD*��L!b�F]aCfIND�d��i�\<��x,�}�Nп)#���2�fs�d�2)�l�9���v�����|����Y>�T�;yY���{�G���H�X5݄{-��ǿ�YI�DęnH�*N�Ʉ��.�������=5�݈�"��-��k�W���q_��&��A���,`	rd@��D�$������y�1����7Q��Y��6֊������m��4�<+��i�A���kF��0rKrh45�MM�eh�۵�݄��q1C#䈀�O��U�!~W#:iB���K˗����.���YlE$Iu��IS�M��xR_먗^��[��9�����7�𖌺4L����C����������8iO��\���%�h��fҩ��Yl�2�|Fc��t�\&۷Pᅊ�~$C7��h� uqwZ��e���Y����auH��b��=Ԇаs��9{��7.Gng	�^�kM�!X��}Ϯ&��K��A���bA�����T1������b�Lv���]Vj��T���-�q}�.�r���$'���^қ
�bO�����~����4�b�]��!c�xkɏ��<D�^[P�-c0i��z�Q���I�4{���
��ϟ��!���dޚ�X���#@A��$��ϳ]��W�A!�K�Cͻ�Ė~φ�畬�m�}X��Dv�@�﷤�I:��
[u
�T����sLϲ�	�r�>�N��-5��5D�s�"so?��W�~�7��X-��y�w�!����]�a��E�?�vm�n��dtj�F�:F1�s�gY�VqN�8���l�V@�Kn3�X�qa�U�?b�Ր ����� 1�3�~\�^q����oS�~!��7r4���s��e!�$��zG�����X��HpvW4�:J$������Z�+���VO�t��.__''*��C[L��Uw�gS\�Q��8�NY�'��� ��)>_Y�0Gvl��vr}x�d%�w�,����-�+?�ZQ�v���1�˘���l1�����n�7px�AhMJL��,g�w�#jg\�i�v۸V�u��T��:�~fł�=GXh�GB�B.����V��s�Gݝ��=<���TU����kN�9HT�h�X��ww�
sK�����"ӰFどF$ 	"\o�%I�xc.��Wf1���Ł������d�x��h�sY��^�)\e�(`pT�@�&�	J��Ol��*!�琲������#�i���2P��n?�R�&e������jc�]��ק���ث��_�eg�Q�{AѮ��)0�N�0���]��2E+���rI�nrWX�{>�^��HZ�0����Qb%�e����	ĺ0H�G��$[ fJ |*>�҅K�����eZ��f�X�ك����{j���#Z�|/�����v�OιX~�L�7c�P���NV֍A+~��]em��H�7_�,�4����WB�ȟ�`�^Wx'��1�+�=P���mq2)4-�v�K]/f���{�&��K�����x�</ɔ}\i�qn�>��̮��Wq���sK�DOM{�����<XC�1�.w�]�|��	�b���ߗn�v_�H� �M�B��%S`�;VG|���e9���g�*�G��	��%C�\�U�ࢇ�X�+�2?/��q��w@�;������`����#��ޚ���~x��}b�{SG^��^&���h�6������%��{lH�`V�����n7�$\	$m@�7ư{d8���.?Mv��*��c�$�npB���S�ߣ?����-I��G)�3�.Fu[�W�D1�^]�6mc	���J��G*O����T�_����z1]����X��:e��=T�"%Ѩ����L�����{˷�9ZШ+�l��*#&D\
���˴s<��������i����G���x`� Y��R�.[�!���jÈйf̩J��� �tɢ�r�Z��AK~1p���.�.��(�?�P�W
9�� �R5�w��UR>W=�����b��O��Rm���X#��I_�ݣ� =n�
N�a�IL�mq�M�ұBv#㵥L����Q������o�48�P�G*4�4�6D�����/��MW0?�L��FY�M���(/j�I�9+d>�ŀ����=fա�4��`�����s���?�j|zv�hN��؁��� ۟�\!�o�B���1U�SN����E�	{�� ��O>����RM�Vf���י$��ѡT����'�hO,>�6���gT_m;���=-�O��uT8�ڵT�ms��J�q�%������3̖���{7��C	VYn,�Y�]��h�2�^R�m�9`�gU�`�9)�/� ��>�����m0���w)�]jW��丯V� �X���r��Firh��*|W6섪p�1l)ݡ�/�v���Y9W�:~���.���o�K������ջ�Z�$ڇ�#r_��ۆ/Rܘ4���}���u5�?hpUr��Z�"���v-���w h����]���h��dSa�!);��){Y�(��1U� 	��O� PƤ�����V���fn*���m����m_�	JŅ������lb��"�����=nI�NW��1��u��MJ�1#[�
�xf�H�3���V�g̥7ewu�Dܒ�n�g���VDhU�O6���mT!�0X>4ޕ	c��P���	����7v�M�J�^x���NNe�ӹr�+�R�C�!�&0(��HZŸV���>��}��'{˪;���:|6��/ja�;���ٍ�Sa��0e!lt-�p�YwJ�{h`Q8�2~yp6B��J��k��?�����C�݇���}4!���պ�8�IERU���� (��B�U�Ua�y�N�n�_F�!S�ˉL�� rNdR����y��r�a�es�eD�)`��5�����Ru��/~�`�m��G5�3|��4;]8w#�Hxi]n�ͽ 6}ch~�c�\z�]ݲ�ILu6n������3���n���k��lLa��/�x(�aF����(ӸU� bn��~���O���x\��$E
�g�\�up��k���������ر�ٍ)|u�5���
�Z֌j.b�h��I%���,��E+�{\�³�4G����˦�jG�Nλ�1@����h�I�K�� ��8����y�_Pi�|vR�'�������^v�7��2.'d7[׫jh�����Ǆ�����m����x�k�9���2��P�8LI��j�`k���nHTU�.�k�-�l��)ѰL�W�m�@܏� �gr��r�2�tǞ�z蜋w)����{�E�W�l2�s��!6��G��P�R�2�����>7t�6v�0���CCW��Ŋ�6�/�*I�R��jҞY���2Y�����������a��7I���d	��j����&�.Vb��f��H���|�<X����ŢwH�N7<Y�Ct��,�@�m�]�Մ���R��6�5)� K*���X]�V2�j��Թ����Pˁ��&�VD�X�O����^ ��j�D�	� �`�Z����$�.+�(��	tt�v���;Bۨ�8��O�w�V�LNG�a�R`mW��{Hޞ��5�Z�\Z���H�6�4�q"u~O��d�^W���N�yэ�b0$7�R}�4��#��[���g�$�W���KL����a~�,�4!d�M)���������Z�g`�:I�鴧O��]\ؾ"�h�*�tQ!��o�&�I���m[��P�-�G�_ի�Oi@��=�B�_V�{i�*O��1��9�@Qg`���q�~��e�����_��
,���YFV8�c�|Y�����@��ӳIr�6���4N�����D��Okmur�~Ul��;�3�����D6�0	2��,����+l�Ֆ��w�8_7�4;�~�s���[g�������*�ny�*T�Nju�9׉Yc��>x4,�}�6,$N�%��l��v�Ho�ȝOk
���������!`����h~��V��Yܯ-t(]`g���CI�%�0LB�,�T1Y�"r�� �pN�"��SOUoP4�>�Nm�5ʫt�MZL��:M���(G�:�h��s�i��,�D�;�ۜd��^�=��ˊx����3�2N	m�	�-�/���(r�B�9���rV�@/��_;�h�z���W��7'WEMi�R��S�<KL������� N=&�����������g<�a��ب����OB-7 ����_0��d�>!T{%�z������1D� ���<XwI<�݅�n�)��m��2�/�~Ԇ�׾�^o�ܖ��\/~�CtP#i��d5��@im��ٔQ=[Rs�OT��3�O�!�R�wԔ|�c���+�p�i�����Źn��'�&�y�:	��8��
r�ږ�<�Gh�?e�#�[[lz,`k0��	����G��XP���/�$�?��U�w�n1���g�*��6�Ӝ7��5���7������'�^j����=�D�B�Y�$K�w�6h��	�NI<���5XCVS@ 
Ĩ�ez�?����x�py�l�bu�!�q%��X�`��y���ۏH���Ba�~Y®���9�L>#W�`����c�)� ����?�F�cٍF<�u)5뀥�<�G�=j�{�	�.��l.%��Y^��6�a�5`\����9t$}	?�w�Q�n��n��r��*Ļa�l������rp~����t-�~��3"���|}���`^VrJ�'�Z��Ԝ�^�y���C_�o�~���)4)w�^��ni+;��W�L��3vLx���WdGV���^8�!6~�q���Zv�(��g���gC1V���eNӖo�9"Ϛ������m�e�ߖ�����D��4<��v[���6T�ؿ�CI.$Ѧ���,	���-*�}�.U4�}�c����I��_Qr_r�LQmCT�R�)�}�`����EzϢ�Hr���G�O��[�lM$�,@�I*U
�W�!(����D6��>��/7��ge����e\��O��\e�0�{/\�1$42v0� �#>��Uj�� ;�O��|�6�P.�mG.0��8��6�s_�i�c������v,S�ŷ���yn��y����hPF�W�����1��oč����0����0���z��8�P)h�FV��ptV��T�=e���Ȃ�n�)���)Ҏ�����QX@Q���̤r�^m�Oָ4���&6�F`3F�D�x'��V�����bk�Vug:�L�n6�.��w����Z=��AOk3�:������+�C�&aG2�w�&�k�Σv�j�u@0��uy۞�{��!��x���x	��P�R%�r蚚I0]�,y�c�AօR>�߃��2�2�<C�Z��n��O�|� ���W�!NH�MkD C�.�7~���1��}Mև�t{�{�}\s��K-l�����S���X��p�6�%D���k��t
����D*��;�"��̣���lS!w��!��#��3 l׹\ܔ�қX̱#*��w�Ho޳�zʻ�7��1|�Dz�����7䘈��scY�!1����sF�F�ݗ�o���s�����G�Kd`뾦�9��1�Uї�����ޡ].iF����HN �R�
�o�>��di��>��//�;Zs�1��{��7��2ky
V�ބ�*����
̷�Zfi;�F��*�Gˌ���Q,�B��#2Бɋ���w^V�n1��]�fih(,l�Q�el��%g˝��f���ÇW�d�Z�%s���7oe&�Ɂ�J���T�g	ƠL7g�0�^��ݮ]g����T��.�]��ò�#m/A��F�~U�N��:�\x/��77��9��TD����hѱ�Um.�,�fw 20�-�7z�j�h׺[��Թb� L�ۥ�W�	�B�Pث�df�h�Y�5i<�[t*�� �kJ(�E�ӛ��hO�/o#��4��3�~�W,��ȱ�ZN�K�����P*F��� Q^l
���[�fY_����G��Xǵ�'	�*�}E��=���d"���PO��ݰ.��hVm�h6���p��E��Ů�ظ���7N�'�a�����
s�َ�oy���^��o�w,�(+x'Ȗ����=�6�,qwdY����mu�A�8�8��8�|�oC0�(O*/��K�w�mco�|���-B�ƚ֎�AM��KiFD�A �v� fA��;#��a��kTo5i������)$k�����K<��ݫaE��x0���F��?��sr�*�^n湿{�����M�����c.i��3}��Mgc�w+�v����S�ȇ�?���,����\��?�e���.�=L����f�X�T2;�z��d��NRȅ4%�&�&)�w���F��t7(΍1�$�.�u�%~qֻ�_�V8� ���k�1j��DΥ�Vǈ�Lܩ����kD�/KI�~�\��$�Y{�\����E��&_MM�S��;g�5��)��&��g�82��f�����^�^�q�T��Y�v�������4�\�YS��C<�q\��,���;�/�q�G? ����Anc�rMB�eѩf�fR���;��3�&`,�� �⡯U?�"##۩�.xS=
�k����Z��ƻ��O�E���W$�I�@IR�$��u��Mx���@.�T���-�>W�i:��˩.�k�Y�Q����$�]JKL9@oAqW���]���a=��8�{b'��`�\y��]w�e�h�Ue�. <�C��7��%�G͌�_�-1U�	|���(��&N����,�*3�P+��m�]��,l��^���AqH��LT�Y��Q���Ӎ)�Lj���&���*����Ҳ�?K�.m�s�AI�L�x���������V�-��t���;�l�3}�og��1H.qm��5g?D�aw��) P,Ɏef�d�M
2o�_oqk��d�C/�y�nlK�H�䂳&s��3�|W�*H
����nR�>X��>�:_�ۣ�Y��]D!|d���&��MηbW����\�� &'tŲ��-wĪ�Q���̝N�F�(ݯB��	�a�1�C��JoPFL}`?.�)l/�I�H����A�i)���pkb�eG��� Uv,�2��x����Ǹ�O,0��+����K�n������<�������)���f�]�����L�5�h�.�sM��DN0���7Or 	+�V��/&�6��yW	�gt�Ub�=�.�+ZS	�q�t�ʵ�	���x��&zL$�bmE��P���2���j����M�gui���N�z���rp�}o�|T�b�'&]
�Hi�)���>�T�sn9R&�v��~~ ������g}��zwǩk�?�"��Ӿ�F �nFn�B!ܩ⊚M�[o���W��F7��8���
�xn?�OX�)�~+�C�J��Y1P�|Sw�+�e���/gw�ܶ/���KB��j��F ���z��kČ`�
_�C�����K��rI�B�2O�%����q��Q�&N��(��	�h���7{���h=�*�P�Z���]f�E��@M�>�g��#�ً!/�,r��p(Q;�9ʢfE@z�WK��-�u�JQI�M��ː]���{� ~+�y~V�zm倩����Y~���P�Pp�S����R?����0P�Q��"��<�I��KM\,���m+�Oo�=YOD�y#��$�t:S&�OD��	��3���$Ş�����[��j_�7��N/��Nܥ�O�D�T~�'n0� ��sch�lN2�3�s�LE��S0����i�z4���E��gA�[�5~�����C}�bw�\qO���H1֗���dkR�Mv�EƨL���x�Q�9�܌�f#��f�]:O`�*���2�KF�)4��p9J�G:Ń�E+�5?R��؝(��u��hv*_�E�JФ-�ʰ����d\HG|���sJt�e��U�����g�;���C��I4��F_���k8f��>QdnwS|1֠������X���k�8G��p�sL����ujA%�p���Q�����{��ګ�4��+^���	Ѷ�o�}�c���%ľ��Jt��
�\5���C���L3-��;V��gh:�K�,X�����_��U�k����q#)8���i�J�Dz<NV����eaj�RDM�~"�R=x�����W���������)J<]�}���x����}GI�x��9�~��-�����S+��W����/�/����KsP��Z�'��wz Sz뾚��T��zh��u9�tMC�qߚ�)�n| wӴVѽ�;Y�RVT9�X:���i��vS'�C
�!�3d�����8؇^MJ�6���%�1��!���^�s�9wx4�T2�Um9\-
-l��ݍY�|)������m��O
�C Wn^PK�d\��0
IBt([5 ����DiȎ`[}%8�@Ih��%���A`�*�L�"�������V�^!C�zq���'��L��q��^�å툖w��ǃ�Y9�h����h�]���㡡g���C�8Ŀ�,�X��}kD�<4�G��!A��2��G�K<�i�@\��1���#�ƒ@���$�8:��-|6�0�n�:3b0.��AB"��q�}��Ň�ąGث�j���l��HL��A��Fr�v;�"u�^�V�����JCC^3����J��v1��e��p/	MW�C��7�`uȻ��|%a�Θ&��n�<����?�� �<:i�b}!��5)@���+h�8�ӓr	8|�}Htj$:k�9�id�����y0��UG[R!|��w)$����3�@{Čy�� ��-�1"l�ɞqvwVώo��>�J[�$�$�e'!�"�#�y��,�2���=�E0�@c�/Z��J�a
\''}F6���S�������ÿ2f�:g���/Ξc+4o/)�s�}^��0���4�!�gs�śB�`��@:� 9��1�E�M�(m���ok/�ׇo1ˈ��~��,����}O����I����%�PѾ1�?���c:{U{�S.)��p����X��MM�XϹ�uqg��v�����י���ʤ�?Ns����~�8y��o%�^��S�2&��
%�R0ֆ�m�0�}���/���~�4�A�?â�V�KĄ��=��&��r0ả����}�6��:��-��U�t�9���b]�d���>ߝO M�%z?��~���[�:b��`�it\d�����%p _�|����{���ED@�m�EG{u�`7���H]��#�뗇�ǉ��ly�@��h��O ��Sf'�KC'��������o��x�e+�\�&�}g��!���ӸB������)��n�@zr�"o���KE����+���'L�<9�4��<�"]�Z�_@^�&�T���+H�&�m�:B*N�H���|:�q��[�Ȟ:r�a��8�
��M��v��ňg�P�C��WP#oU'U7TFA���/�Q�o!)F,Ž��B��3	7�>��jg�����{�4���3����ڟTW?x�g���Z�%h~Q� �e������R�ď$옾w�^�C�K
�4��-��~$��^ľ��`D�z!��,Ѷ �.��*�݉Q�ǳa��쿴�'��qpt��m�,��D񐸧��[��W�����7 �S����{�y���0��KM�!��
���',�:8�rU��V���(b%oW�p{v��ʜ~���@���·�F��ՎV2��̉JR�E�^�P�Uk~��d�"�F6ҳE��u�l��΅�汣�u^ը�B/������o?�Bmd�i�!�3}�tn�񋛻�jAi�B��9��NhX>i��Pw��ڶ�w�ѡ�̛/["#w���$�'O^D^���=�
9�M�!�O�G���7*\��v��HOly��#�"���3nE��̸mGN�rm�� a�QkL?�O�I�dd��^�sF��߿��*!������3���(�F*6̭̒�.Fa���u�r��j�~H�	�0�]�x����4\�����\����4E��s³�L�.���2��w�e�-�W��6��u�E[hLCsM�����t�п���WtXТKy%��q�a��g�5���[�A[9u�W���,�^d٧�c{4:-j��?�.1w[,�"D�l�P�I��ْ��OrX�#
����Ԉ�'���y7ǔ�c���Tt__m�p^Ѭ������ŏ�.S��`����^��?����h1���	�T�,*�����%�S�P�\p6�C_��^�]�|5	��@6O%���6���%F[�.�}�MW��9�L��j��07E�4;�T�0tq�'Z'�W��k��&��V�Q�S�s�zT#�Gc\��rx�,ʃ�=@w:�A�}��]D.T�?pF����R=��%~�}��,��{���$��>`�R���a� �꧑o��w4��T�	7��̉��TI�ʚ�+l������݋�7���.���Gцy��}��s�/�&�_���@��́�Q���jJF��.v�����/���h ����9���V�F�D�ο�?���N�|�ĽN��v%V�}��b~g�t)�F�qh����N�+��8����?P�[�� �
0]����8xG\\�Z�'��R�:'b0j+���������BکLi�A����[�"�Ы�A�c�k7���'��d�ڵ H3E�<�&�Q�����d$[?��l�4cD��U�U�Hn@�C�Ů��= � �6�%-Ѩ
&S�j�e#�~��DÔB�2F��n%�O'��7{F��	5�n7cЏ�+�Z��a��~TZ;�R�>���v��::!�'6���3}N;���GAߜ�+pb5S#�yp�=QF!#X%��1�GQ���˶��*���s��Wu�[Eц�]`�>����>�-��y�db�E��*����(���j���l`�0Ai�r��==�LWt�T�q����$)5�Ƹg����X���uba!��S�?�(��d�����MY�z�͛cx���/5�/���U�fIu��p�����Ơ�E/�p�px������˪H3�.��n��GL��C�-�7�mb1�Z��W�y&&�[E���O̅�Ȁ-?��P���;ެ�a�����!!�r��G�n�-�"��`�A~�J5|wu�X�[��6�$u�rnj�^��*�A�%��9�@ŷ���<�����C���%���.�U��6N� 2�[{�^^ʌd1��y���1I�>eO=*R� I��A/ՎP��(	�r���6�L#q�y!��ϙ
��L��=�pz�>��D��q�Z*U�0P�7��{�]9�D����-U8?�&�������%�>_n��@"X;��<y0��VkH2��ܙ%�7�j��V$�,]����9)�>d{؂]h2`_�j�
��	e��4� n����	_ ��.��>��AVag#^�t�y��SBLa�9#�]�aGyi *�P�s��5p�x��Q��Ot��&�ݦ}�[8 ��6n�w�N�u3��d��!���	K�7	��#~��� y�<ٗXj�Sa3&�����_��J�u�0�w���@G��ʼd�A�,!�h�0��O;�x��׾�����'�|Ki���9'7�g������BT$�udZ��D���(��7]��נF�~���K����DX��̨ڶ��r�A�i��؞�֒�F� AO��ݬ%�[�c��H��4Y�d��������.߆k�c�L|qR��m��/u`ق��L���8��Y���^�dP�Έ`Ӿ��4��{���v6��:8-:��,(�ʫ��)�|KG JQ���Yx��&�~��%33a�xWED���C��z��Ҧ��'e�2�k�j��;�IEL���(��<V�T�.E����h/
���5-O�,��&7
�'p$+�Ds��;�XDo.�@�Z(O>�r�?��[S�d���`]2So�"K�0`��Phħ���P��y�7O9�,�E|��s$�W�lr���=D��9� h�F�� 
��τ{y�={��v�6ƴ�4	�
�Ro�Z���2����A���5Й0�j�|���%��mi6r���� /AKj���rB���n�=������{=�L��;23G`ȒKq�������u
CѸ��4��3�ؕoGxGZҷ_JUWM>�Ck	'&G_j?���G˅�I�Qê��K�RV�L�6�؏��/�LY�/�e��+;+�,_������>)	���7��Z�ԍ�n����I� q�7?`�E@7�M��(�x�;t��fT�~�3�]H(/r�o�;w��A���]��w @��w7vf��k��6cl�oA�h�]q=��Rn�P8�����5�����A�F��W.�%�vS1e4�8��!�;l��Յ�0��u<yU�E���2fĎ �L�0���u�ݝf�;�ɝz�(�a@H���wO0�25�K~��c�7M�"�R�RTo^���F��U��Q�g%u�1�*g�[�E//[�mͨ����b����h7���h\�(;f'Cv�kO�q�,�_|h5�4?V�v�z���l��"'��qނlxq��÷���Wa�)k��e/��מ�V���Bz���t�5�/���\�rVu��d��W�څ�4	�4h�e1�q����m��ځ�בaUe7�)���B�56����O9k=O�`FH��<5hc(a2�z?EE��
q���+B!K�=-7/���bB1�����c>}��+1��Q�P���x��ڈ��.E:AA�1K|geB�sw敜U��_sj<���/Y��V�����LC�A����!�1�6!�0��
�؋*	��@"�)1��⚫�>��{{�ޏMv;[e�T�&jh�|6��o���Zp_y��:�h��K>w����@?�� ��t�->B��{��s�s��g�2�f.qh�g^�I�7/U�͘��	�Ñ:�4��zdy+,��)�t|jO[�t�8�DĈ��P"w�F�A��� ��=��d��:��.(X&q[��M���3��Й�Jѧ�ÿ���=���z��v��\E`�Vu��5T�6^S�p��Ax��xn�������u��Kʫں�nx*�ivoo4�@ގ`��S��A�ݴs��v.H?i��ff�k�E3<��Z3��Cx���t�Bc��˖3x������(����|$���2N�@oM ��3O����OWO��6d�'#�V�^0|-�^��לJ�/�:��>�`��>F��]����\'����A&�$����>�F+�����zٝ��q�4=��|QՅ��+�5f7��ۮF*̌FQL�5�pD�T,��׉Ȧ|����qIB���wQ'i`�G�@)�~#JT1�o�����V�a�9�,;�	�էn�|Z�9��K�dB?�I����tT$"$~��	X�!Ӵ!U���nk���ӂMN����*f��>�0����6	�Ż�$�3܀�y��&��]})&DK���F��>4���!�ObV�9ͫ�R��C�5��{Sg�����יV�Z��\9 I!��";y��ɔ�;�Ǽ�]��q�n�1�o��;���������|��H+��������z9e��I�$�-��d�`(�`�aܐ�TK_�21-����~8��H���k>���2hd�����mm��2��y�Y��g�&���������
HV��a��?��kj�>�>�Q��E�-��FЗ���~颸bA�҅��kE�я�^��ab������b�1�
�����]x�)����z��_悒���q!�Q�Q[6l,<��������p�*2�݃J��Ѫ����/��yNu`�dr��"�"����W|4�M㒉�_�
&Q��WL��rxS�~��v��W���V$�k�D���5�ζ`TE�B2�˃��¦)�=$Љnw�A�[�w lX�Ϗ	�;FI0S��"n��0���rS��4[�%��o��z/�r֠��;{3��㩪�Y`�Y�.Su>�߆��J��Q,5��=o� ��`.u�s�5P���81V�ٌ�5.=�����WqBX��ϕ��Y]�wԯ�ܵci��ߺ���W���� �����>���@W�ґƖ��SѴ4��m���߭(~��ݙڍ1��7��'���^W�$����zL��'Xޣ��sv�	ˌ�9H����z�[NXp�
B,�1�%^��B^�^����o�Ē �n�69�7D2ږՕ0�.#�����g[���ݏ �"JH�_�� ���{K� �9�4Q�:��M�y��ĶV�a�����bU:U�'��m)o!x�[����$�[N���Up��j�m�<~,�S�z�K�K��!����֤2���K���f��j�A�7�"���"<��ĨcG�MU�O}ߋC.�>���!�֘п|�B�,���[�'ܺE��O�O&yN��#pA6d�|P�u�^�|f\�muَcf�g������t?��~����HE���4�xH��yFh��IbQt�o���6�<�}�/����PH�&6l�0%�v��P��^=}V�p����":�+8�Κ/���� ��3<|���Ԉ���mPB:�o��t-r�wc$�c�NP��T������dإaϭa��0�!�/�rN�K�Nܺ6
�%��W���.#T��~��"��[lB��>�x0�*�4�$�+��Ÿ�L$&y����ᾔ��� 	�<(�E�ă!.[�$��a�5-9.:�	nY�6��e��0����&nz"R���� ����=۲���? ��hJw�25���قab�7���Y0[��f�絽�Ƅ2>�z���.�C	Ǝ7��o�Z�݊ոqW8b&�NyR�2�۞h�*h��o:.��f������:�%s��s��8��h�G~�#�&�0�P��S]L	Y�m��Y����� c�7\�1ض���YZ�U��,ʋ���˱S��$dNP��׹��*�2�;f��⾔�*�!yg�3qߌ<J��E
���0�ri]E
���n��\m^���S���Y%�L_R4���~�2��'�ڱ�,V�)�A����9[�+?��gW��޻f��{�m�u�%(O{f�(����P�ʱA�yED�4�w��O���X��kZ�k��B�[	n}������
'n+�4����)dc]&�
(��8���]ߋ� �^����_�FM��.;��Sȿie���E1˼IxU$��d�y��}#�g�]�d�a+�6nQ��U/�ez���}��Y�p�����i��9P�C=^*k��=*��h�s��� 7]�:�ue�0$�n�)��jH&�	()u$�
#�pP�03�/����!��O��@��$��[L�`�KoY�@t\���w�{�Xu�zdl `y:o����� �5�$���y�%¡1b?ځ�M*���&ɊPe����d_
�����%o�b y-��h�ʤ[j������DH��WBP�ŀ�=o.(YS�R�r��)��?�ɺ��r�6�u�P�l�غ���^w��<# �),0k�ኰ����=ϐ�X�������N��t�N|��'�]�M���E��j��K���{X�Z��`�vop_:�-C��W
��v�ʛi&�P�m'��0��ӓ�t����C��Q�+ǃg�d�9�I��M�� �F"j���q����������Ed-���$�8r|efΙ$�
}u ��-�=7t@���dF
��Qu|�j��-��#P;���˚�}掑�5u��Z�ɘYL�ԡ���H:[�5�����uTފ�4�p��T]',N~����<9��֖u����� Җ�AFaVg�F���\4��HЁ����e��H^7[��9a*J�΋DD�Iv��>u�ڀ 4yUȊ�.39��S) )�N��A:�<���6?�@�D �U�tZ�%ow{Qe�`I���)]�nL}9րO0IɬW�q�	U�*����2u������Bcf��S
H��m���=^Kx�Qi4Q�"~Հ.�G�����%a���n��u܆o�I���� W�(��������/��f��D�M��"��<����4���5��R��c��7SX�$�"����7��~��p�b���i��?�d�=L;�C��z	rRn0.��Ι�W�-#��΋^��v\�u�-�4���ԁ��d>b�*�뱓��m~��3��5^���(W%Ye��-xc��o���v��x~�G%�pg�)M�yb"�T<����,N�����0?wtb���E�9�O^*K�i�9F��mQ�\ �-��d���E�p���tj�E]���5�H%Y�S����^v٢�lV�W@�ʓ��;[����'�̎�(\K��r�+�R��"��n��	b��I�W���d}jk�1�Hk��ws�,��{�t;�c&3������Dל7P����z�^��:�/J竔{l��u�Q��� �0��9�ĥ�v[bN����#2/t�4Kl�d&<Q����>@���B(���Cm'LNԊ�u�|�و��I+��[�<����z�dl�L���Mm�6�;��9��/��h��%�f|eQ��r���=h����CU� )s��72�&���6{�����EG�{hۜ�	u�]N;�q�>`BK��_��`���GB�>J|z����@�C�RA<J>��ĳ�ʟsQf}�H=�M2�nO٣Ʊ��R3�,�4d��W2 ��re򨸓t3��qXʷ`j������`��~�ՈT�fv�ܺ�3�fL*�|׆*�x'�mtib����z}eG
�v�N���jц6د�z�|y�`�!�G�-@���������E�r���̝/�G6  �K��P2I� �������d?��B�L��l��e}�!��ΆAsu3�=����I���(a�\���H�4uex:�����;�V�*���*^�fA�_�
��t����~�j����`#���RO�����;�\)4��_��z!Y�~@�'.�]��?@��9o��Tao�wO
�����B��qk��4ݵ}�Y�Oc� *H��P��.N��?��U/b5�QA�J�[{6T����:%��D �2�=�4J���j��ٱ�H(����G����)Ӛ�p.Χ-ZLh(v	;,��ōoxu_�����G;j�h�)1c�%*�6�6[�N'��N{��R���mbVb�&��Q/�?�o[�A�3�!�+8�q��"��#^>��,�i��	�)�O�u��f��5BV�N)�ami��O���(��K�e�X�tۊ�����>���������>���qB�y�XE���A�CF�.��?ϯnn��mmr���	(�}#���ۨ�}'ڥ��Z�gó��%U���㻢w�4�t�w�>���F�!��ԭ�>^�1������.N�B��0����@0���C����h(����A ��,��U���K$��T\����+00NֱT`"PL2ב�#6�LsrkГ���X\Q:��"�2�#ù $9�R(%`�]�Z]L�E� \`{�t��C��Ӳ�0���	 ���]"�����6�gb�b�8�h�C]�6�����٫q[7��4��mH�J@O>��W�$�z���� �k�5HZ����_��Ԋ2�BZ�xs.��\���L�#)�[�D�`pC�<ej|\�X�P�� �,�o��Z����h��ǰ������|dPYed6b:�^��� �E"�	��,07�n&�N�ÚM�"���(�}W5V�+�:L�����a|&����+qxrV�y��ۢKa�2��U��.��7�]����wǳ����"1**G��]��,B�N��]��l����Lm�B?���I�^�dXu��I�V�7����ӧ�;��0��Β}��Ql��6�ѧ�0)�ij{/�M�v�g���{��#4l�]{(����a-�dIr9	��/��#�͈h*°��������.Z�O$��?�5��������w�4���]��d�Nޝ|�1H�R�����L�ӪK4T0�eUn�W��ԅV,�����Dթ�ᲢO�@����.��ѓ���C�T���iy ӌ�ɯ�H�(=5�_���4-�2�<������b�:E�-��X�BΣ{��1x��O���F�/"�k�h�+�&Ɲ��Ax䳵:^Ċ�dw�#�dj}��}ߋ/�ěl�2�J�D"�}���A�~9L��#��p��^�޲N����pP���(��u�ѿ�ʱT�];��-���Ew��B59���{���u��4d���zC�[!�V�K�t���`5m���_���V���|G���ʲ��8�N�$����kQ{Ȟ%���=mE��/Lτ�̬(h���F�B�/#�C?-�V��T���3���Sz�gZ�Z9�	����Q���溽j*�"ϴ-���l]�Z�VM�֜Z���h_C����Dȣ���L������&����԰��J`��pO;��]п�*!�x��=��9�[�l���ő�4�X��I[�1n*ռp���٥,���w��kΩ}�l��U�mfT�G���@9ro��y$=3t$���%��`MG��n<�7���Z���P�i�0��0��>�.I�[�	��2�~
�?N���d���;�ܙO>�6�w4������\.������Т� P��\��BQ���G�x�0^e3�C�If�����Fck�	�%���J&N@_7��洫U��!W�=���ʜ�K��u���J�ܩ��Z @9<@���zIx��b�ݝ���Ќ���-�^�����b�.'�[G�� I��1��i�\�V�t�){l�.�E�b9�T�F,8�8���'��x����1�� ���l&"U��#N;�u�N�Eڂ��gN���β��0c�����n��\7p��L��aN�g&�^������gH���:!%�d�~�cvW��)������z��XU�C >��U=��zL�G����B�����̴g�>�Q=�h�����mi�*�@�0E�"�^�ȺT@D�-nKIK�e��B�?�X����	��'��ԥn<���w^�fdPF���8�N&��3M$�Fsj��$���?��``�x�Xdz�]��-,��:4�@�a�N�j�
�U_-1���M��Z,ud�K٥�f��L�D�*D�
�χL�Q�1��ԝ��P���(�Wӑ�uad�\C�vQٲ9!�#ܿ�]������xݪ���Wo(e�(:�Կc�p}G�_C�kT+�=}$�#�4=~ܯ\�pV7�BaJ$3w���� �tM,6^�p���������a�ޏ�W�U��S�/����W)j�?�y����I
�TO��,o�n�SQ�A���`|��x�,Q����#��5{���������I���}f���
�-�:t�7���{�HºD�Έ>����H��3Ǫ�}G�Ow/�zX�]=]������IwL��7K����4Q������o�cǢ��Le(�Ayw��8�5�,�� Gq��8��L�f�l����d9������8�R�����'�[&�u���AA�����h�ul��'4}��w���I���� �j $�l�.8A�yٔH���� �	����;?Ӿ�P�% �$[Kͺ� �]n;��^�Q�<=�JVw:qZb��d-��
;kާ	I�����x H��U���n����*�N2�y��&��*E�"Dd�a]u��SC���j�R%�%c� <u�D	Re�B�`���e������x�}������Ю~�Υc��	h�RvA�0'�&�9����lx�=^:��`�l)4�lF�c9}(�Lo�[?:�C9��73�V����5�����#jz����T��3s$�����',��Vݝ5�:��' a��z��`�l�ְu>��#�r�vdQ~�{|���Q ك�K�)����[ؠǕ�82�.��/ͻ����Z��=.2*^��~8�3e��ڢ%
��nrw��fq\6x�)V��`�`t	XY��@�a�aXxZ���`*d��7&���fq
��@.1���Z�a�)	�9-�%1v�E�e�Sd�,���D�'�V�'�~S7�Z`��<rj$Ĉ��f{a��Yη �	Q	�D�w�%:���q�
~��V}F��Ɩ���z�r�0S�V�ɱ��	�Y}�-�|,����)��w��3k�n�~u��<b�o�Idc;��E�E=���nD`� ���eQ�Mɡq���!S�)�~�KXWgAY�6<���.�0�6v�o[x/� j���,Q?�P��G��,A!T�dVtcp�VU%2Òa4>h9��K�C6nE���'~nՑm��{��,�Bbh}��b�)N�]
,���⃀SC�cb�_g�K����:��I�i���_�`�Q�_ZŖ"^�&'��}�tK�(���l��?d����J�@:1 ������i���>B�Ɯcߌe���j0J90�_d1��_�a6�P�O�sf8���������q͂��Br��멺ix�&�NT�/��2U��O�V=B(y�0M:
ʟ�M1�&zW��#oL8��1�N���h�N�x�z/	��܌Z�؅!B�{��`_��J��!9����Ǫ�z
��u[�z�Z�����^���r(�������!^%Z,��<�o�G��E�u�C���??`���6_�O
$6˦�'5�Hxl�a��W�+b�c��EЖ6��^�ʪ�&�O�C
����"a�̃lC�&Օ.�wX�6%q�SI�)��1��w3|����r��&"\�l���������4J�MR����$��;�=6�THo��Ο=,QN�M�R��6s��W*��d�X�ww؇�-Ȑ��]̀�h�:FM�]У��s�P���d�|r��a��1!ѻ�Ѥ�j1�i z���RI6>��3�Rb�|׀,U������i�ˡ9C�+K#�#�1��ܜ�X�I��~�JL|�c-J~����g�T���_����oM��2�5u�R?�3���qq�L���z�{e⫄�8���mok��Ċ4+v �At��n�*��J��?}�%M�G�eD��t/����I��ϝ$���i�2��O�+79ͭNU\9]I�3QneA�'��?-�#���̤���
��[z���)���a��㚶�S�e�:yD�V ���8���z%NZ�[u�d����pN�[�t�Mr~�C���)"�!�a�II��z�a
iiW`ȓ�ޣq=`�J�^��6u<dm���2b=s�t<8��L" ���aT��gD�l!��g@��9`�����ox�d�R�te��Ցِ��CDp{�|��F�6�ra����f=���]��asuA��&�=���@���^��s$��(y�;���N�Ko֑�������4^=�us�~�sF���G>���k`q��i[>1���5��WO	����:Y�~&v*�AȘ�W;k5"�����n�訔U��/҂0bea��|����!x���߬z=��L��#&VP�8�85t��а$�w-l;a���OZ�:1�		�zǘ�_.�D�rg1jWu���G����%�\�'b�ͫmk�|����8O��o8��S�ZC�M5��K�6��p]G�Y�8�.`x�:(w�~`u(+s{ߘ/���A�� q{�H��)�B���4a?����7J�C�����˞PS: ^�詛m��d���������7!�a%c��l&<���� a�L6�QS�o�=]�3dcMi,����Ki2��ȷe�V���D���Dj����w!�Iu� �ŗ~� ����{7���9�R��� ����b�K!~E��et}��P"��j�_�FŔ��~Eʩ�k�o)O��-K�9X���s����y�W�bL�H�Ds��x���b���.�VN{��S�qAZRff�r/|� �)s8^0�O�z6��(�#Af��{�C�\�8�����C���ףf�8%�c:Xf��x\p3�Ԁ��Z�w��!��ģ2=��H��E�B��g]�y=�z�T�$��n�]��~h�co4��T&�&��Z,�y�!�Y�Zk�j�G��E l���X;��QƑP5���|��V@b[��t�'3�`��{	��"��ON4+Z*������@�����}�t�h�#�/��&�U�sR�u����g��!%���=��Gð��G	���N�ȣ������l�~e�Ǔ�s��� I<O�Ez���IŞ̴GS[��>���,FS��'hۄ�ށ���ҙ��í�5�����o]sks%߳�ރ�뚾��AE�I<#_O�e̧��l���7��u���_jE5-��á?N*�;��s*���qy&��Y]�TBr����Y~ԇ���x?�i^yj�@�z�%Fyۍ�K˘��ZZ�jz�R�Z��0�����T9�R�o�-r֬nϯ _�'�	M�������E�:ɏ���GiV�~�� *�*A�� �9�����KVnF�=�k%w�����n�8��)��{��lVo���Q�fVg�9}�c��ד+qÒ!�W������zBU�
�.4�a�w=�Ԁ9%�6`'	7�+EC�q%r��{��pY]�1�����_�GrW7���g���V6�x� m�~Vʽ�Їj�tums&�F�fe�>WV���T��
}`��E3�ѽ�n1�L���$�tPF�V���=OI�e
1��XC��53=#*aX��mm���6����y��� ,��4��E��P�Lw��*��L��#ì>T�g�1�y�]�J��67H�g|I�<�C��3�ʓW��f	dN�Q!A�M+_��k���x)6����O��7�J@!KMۘ�#xP�+��@���^�ܥ�G��y�7W3�=���l���
Œ>6Y��z���)��*����ވE:���V'
X�o���U�a?1`P�B�ܥf���Fc�LL?�2��[���05�r��[�_X־r���8BF���9sS[|p������Պ3Q]���=��.�P��n���@��=��He
�o��;��C��@�fH���j�K��I� Ի��UC����g,�L��C�����y���ɝ{�ۼ��a�WZ7�t����+qRx܄�G;	�t9{'m��C7,�B�MǌT��*໘�S��5�`L)��Um��fUݧS�?^z?�_���X�nM����!�G���p��N�$[���F_tx,�� ÕO�.�^w-� �(4I?|�s�`��'ݻ���b�VMsN$��zQ �'�P���rq�����=7눈rL�/:%9���|i^�(T���xriytr�dJ[��!벩��@S1�i
�����8kYh�Y�,�?�2���8�v��h�����z۟m�7>)
���MB�3�vv��o���Vh�N������J4��7����mJ��%P��o��s6U�PS	�U�+,���4���v��d�z�B�D�IȂ6N�N��v_sh�����g�w����e�[k
�ug������4*��Ƨ(W�#_Oj�wM��pTܡv�NV�Κͷh�x��0��"M��L��3Qr����|�;{}��Q�耿��>�{��8���|��d57/ �r �Z����!rzt5�8>?�s�ܣ>x��C=Ь��ڟ��⃥�`t�S���PT�v�|�f�J#��\�h�B�ne|�R�T獕�}�_�z��V�{�DHvF��ԋ���x6�~�nf���ByѿN8?�E�8GD6Org�Ƚs�%�)�J}�h3���vޯqaץ�Z����nEKr���eJ���V5Y� ������rΒ�Q�BC&k�[�[4�a؞���j�'$���"��)�SQi*,f��=��iփ�f�aW�i����_OQZ%+qw�� |�S�"\��Q*�[/'�O.zcAwE�Z�-4�"	ڹq��*/V��#��ѰH��D���h��?bD7	��6��KiLQO� 0���Um�\�6R�_�~&f(f*#v!C�n	 �J�N��p���Nؼ��To�y��>J�%\�2��c��)hR@.2���Tj�*�'֫-����.����mA�	b�tI&N(6M��ʓ�f���R�N�^��[G�:���כ��,��ŞD.fߥ8��,	93D5�7^��̪�[B�iX�ib�w�H�9s>S�*�keֳ�{�I��"��H�.��g=h����˲�J�-MMm�e���Y�u��YI����u[W��wΥ��&�+�K�=bo-�v���;LG�V=
g䨯�T��z i٣���ɜ`�KA�699��az��XĬ��"<�<k龈�(����V-��$j��$sIPs�p����r���a��1�U-����7�#.��#�X�bt���p�T���>�y��$� ��K'�2��Y�6h�r�c��I������gX<����k�t�U7��%qUf:P6O�\�8h�6�e.F�/�$��t���=��ZM�I��Ō#p9È(�Y=U�/9uJwSuf8Ŭ��D�Jc��Ep޾��_��p�g��1 �lR#L��]	3N�G�x���z�]V5�AtlW �I�i ]'�l�������p�"�~��<����m�㔐oR�R3|'�Hu{�p�����EG���o�CI!�?�1Wlw�QsJW�0�R��h���FL�(p��djϜ�"�V�S�[���%
����\wś��҃��`Ϲ5GZ��`ƥή2$���P�a���R��X/�������y� ���L�G�⯏�ǐBi���kx�K��w���[0�BjGYq	�O������[4J5�S��沑�g��O�,�ڦ�R/ڭ����xz>�
a�ٿp��68$!f��jA��#���X��P5��?o6�qT����M?�n���t�a�\�s�Ʀ� �U~�f���^{�]	�
��J*HMD]i�Yg0
�8��g����絒Bɼ{��R��w3��r_ ���0��T��w-�O�>��(����.���ݦ��ǚ����i�
��9��ݞ�$�!{i��H=ˣ��%�h�5�A�x���V���k�@���7��D�Ʊ���Ջ��<:E�W�nL��úE5,�v1,�Z=�6�^�����+;2���h��+/&M;���D������p�N�¼��1ʌ6Xi���0C�����ǲ�%m�\��5��_�����1~y]�j]{�kX�wԳ�j3/6�0�>��)�D�'- E)��5����p�8ÔW�1U�vVh Ѥ��o�<�:��z�. )&A"����� �b�rRh���b�{�@g�Ҙx�;��:{=ag�Ы��G7��o�<wޤfc����$�x'�0��Eo��e;��z�f{V����cܪ�M�Z��MD�.�Z����1�+�+�#�E_$I���ȓ�ԑ��9aI��iߓVc��iNx;l��w�Y+�g�����fn��6�w+�I�z>����R��܃�a��P��$�K��vZ9�f{]��@�ˊBθ��������/`���[ש��2��
��L\w�:ɪM�������M�D�ǣ-C��Hʷ;�o�h(;���Ą�uG�k1b��,|�N��,�M6#N�,z|���a,��xܴIz蘚9������f�y��`�	���*[I`����Q,��g�/�"����W`�[�|���	���E��*'J+��F�l�Y����"s��w10b�t��`\��'%�l�!x�8l��"]�:s�"���M�'@�4D͹���~���R��9"�.C}þ�MҔ�0Φ8����e�l�K ���}D�t��|m��w�v�HH��Ck��w���]�:m�������{ˣL/�\f<d.Bj���y�z��m'a�e�;����kbX$�)ȟ5�������A8�xp��86�JRl`"��.Oi,����W�q�j4����Lv|�ΈN�؅�9q�ƧUH�J>F�;�:��p[�#�(\�"+�<�!�⯉��ل�K�⧜}s 9�X���Mk����?���M~:R�;kX8S��d��� +��!S�;���{��쇽���]"_�������5N�ӂ7�ڼ<�I�.gm��hT������qe�2L����WA��%���33���T��T�h}JTT��d'ԅ(`Au1���N���%>���yӸi��%YA���e��h�S����Z"���<ա�P���o�w݌�}�A^&m�w;�w@;�xjh,k�D�o>����m{�d�F}ZFT����q��:�J�ЙGU%��WR�"Q�Lx����m4����q��5�fW���`�-d2�f�e%FD�k�s3�o�ƥ<�>f=�`�Y��v�S��r��K_5��c�>h8�{P|P�nH�h��$C����2=�H8��@�([��d^O��c�6`7���eWJ��3�r��Z�ɨ��@z_s?�[$R8׮����{�
��t$��H١��^b��.�ʡ�_s�c`��I������:��l�ͬ�]�  �R�&K�Z��k���3k��"!RT�A�L��q&����CE�yu����I@��3�W.,�.e��M��J9�����{O .�#��J���������t8>ķH��s��T��Z�bN�ҝ�p߱J��
�=�ܙ\�iVD>�4���>U��nOn!4��yQ�e���	����F�뾧�b����֬�hR�c2��]Ty	
��f��L/bye_��(�>�|�^�_~
5E.�l|,�|�ac�LCTŚl�����e(�X�����U�s�ߔE�[s(I)����tʭ9�0�����̌g0�*��ڣ�v��n+�9��%!\CA5�«$%H����\�����4�XM��2��G��':`��b������b���V6�an�OGUE(��#u�y�W됋��9�:��������[�E�U�]I<��̓-Q(�R#�|��㉛��;-A]�=��>��1JI/��e�iϰJy+�D��G?�����t48<.�	rd�Ȓ	�u\�Zj�EG�j=�J�`\x�wG�q��b�2��'[�wb�?d1+��^&o�rB�Ȍ�:&�~ R�-�׌o�hy�A�D��Lf�j���U)����󙽍F�*�%�G��b�����)7.�z�J��������a�Z�6���R�M�
�jEA]O�tO���{��x:��$�e6<�1�딿�mGbk��!$�޶�����W�81}�/��@ m�\�|�Dhʙ=��`��K�؎���Rn�r�Rõ����nH�P�ls':�샖{��駬e2��]���b����y|[����txyc�o1m!���N�b�����ʹ�ٞ�	̾O�@U~v��e�OŚ_�K{���F4J��36�Rr�`�$!�U:���F�Џ���	�2䰓���z������:x�S>�%+S���H�)�v��5��t,�w��K��ul?P����Ut}������c��k�M�ovs����^	g(xB������' �n���&/��du�"S����n�7!Uے�}*�1؊��=yx/sY�V��\�Q�8J��<J����x�{zδ�RE|43��w��D�<Tʊ⟐�\X�C��d���IYt���4m�~��~�W�Ͻ�Cq,���+�c��c �B֣�Ƌ׆��h1b�Ul���	81��p�)3��ӧ'k.��0���� �u� �V	�/rQ��Ty���)�\�@�4$��^�cX5���zw��q�X{�|��p�Q"�"cP�*�^���J�xT�*��m��<O�k�`(t�y���W���5�/&�yZ1���z�JBH���R���#,���,u*������CSo\3�#�*OH9�CZ��9;�dH��2Y�m��=��"�CL���1�d��qz��&Hݍ�/?�j�����"�@[X�׊�c��x0{VǶ��,^�2����P��$�7#�l���Ī�i���٩~W/^(]��y5 �}q���j�	�J	�vև%j��<�����J�v˅j��x�y�Sy�x'�R=^uQ̖�D$V��+��	����ȏ��!�*��������˖4Vф��ú�ay>�((�8.�>�^�	:�����
������A�?�$t�'�댪z~6���|�b�9��Ӫ����p�Q: ���9��I`,B\���٢d>�;����%=�ױk~����1�Rns����'P�o�Q��cw��K'K\����8����U|Y5������ ݇���T���ѣDy� ������Ji޻1`^e�W�7�%0��?�+��6(h��/�y$*'�P~�O[=�xyq�:F5[����7�!2�Yki��h�E�|Gh�HW��1��t�+G�C�����������l�)55�xk@�4��q�һ;7��WkA�k/�3u5Xb&���s��?��Ȟ�}hO��߁��S�����/�1fD9�ؼ�C)�;��Y��L�¹C\ ^�☝+$���\���� �t eK����oS���w��J-�ڷ���(I�rP����(��{�<���1J�"��$7�Z5_�	���Wѫ�ύK�3"n'Bj�ɫ�TZHc��Ȧ�bK鶤���'-���ch�^eed�¿�K���X���^2m�.W���ɀ$�P+v�C�ֳ�9��N}��^��"4`��q��K1��錷��P[��v�wWt�,�k�ղW�sͱ"X�� �$Qi}������imI�ȏ���3o{Z%����:��G�����e�~F��io�+��p�Eol�*H���Y��u�d���E����K]������*�&�+{5�A����������l�:ue�@o������$xbO�_�ȸ;+��c��t��Lڔ�ӦK]{���D3�YQpC��\�+�Y���(\��^��� ��0�u�v�KV��2����Ԫ�7}ac�,E���b#��|y�r��yp'������*��&��x� 'E#�$�(Φ9��M�X��;�c�|!F��$l�˪��������+)~���i1�`�?�HZ�=ZT��P?�y��	3��3\����Yd	%�1M�mE&��IتH���t�
�B7J�Th��ONYߞNO9�XRqre�*�FrT�������q��U���:� -������I'=�͔iK��4��l��s�|�̭���r0�J���������Y��!���d���x�8�
�הƥϋ�A�;Oė�J�%�Ͱ�W���}q�),�h�SzmΨ�A�����E}M�	�����YEFw)] `8�T1�?��.�H��`�'�����R����;t}�۱�qAn\Lm���+�����Yq�V7N$=�s�PzD�U�n�I42#�|�#E��_Q�
i|Սp���ާ���EY��Pp�$%��o�cpG�P���)�)K/��u�O���+օ�:�? ������ I �ݙ���󧈱Ez��7�͠]���� �bEN�|f �a��J�D��g�)��w������x�/���-����<�q7�t�sW��[�Y$h����(�,��l�&�� s6�uB�]G6�&*;փ��͋W7��׭;�AfO�~���~�]StW�m ݉��p/����	�|9�+PL�6��^օ���Jw�����m�N���A�q�����+h��\4t���w����R���X��?���)[ ���X{}(^���qW�@�kѰ�s� ��ȱ�����<��c�A:�f��3�U5 ���&Q�!Hh(�;�Q*���Y�]�zʥ���̀�'�p��Ϥ�3�+6������e2	|�n$@��1��ݡ��I9*dS��AI���}u9�rS�\���nh)�#)���� ۮQ�1k�ɓ���m=��c �r����L-A�$�#^��4���Vя�n#�X����ڂ~a_���0{�`�B���=q�ҜVO�sdF��k����-�	�o�/�
W<��r:�-�n��uY`�����%��R�$�|��Q��5֘�G����!n�+,K��3�L���*^7�*�Kb<���V΅��N���)�y+xg�Ò�S���i��)i�3#�i��Bic���qⓕw+�0��s$"�b�Yl��y�w��I�.	+��3���!���7h]!�5֧�t�Sq#�(�Ɋ�D�h�3���,�����j �^Y/�0��~eQ�%��?9s�2��}���'�6�i�#����:(<����:���Ꮵ2�/��J�ݑ��n��j ��;�q@�
{�E�z��×�" �	y#	��^2
�G_��/�G҉�CvS~
k���䘮�t��^��b8��9eS�ˢT�xo&ޅ�%5��WlM+�gr�
�-��=��E����| �zO5%�ᓆ|E&���C��戌�/�n��FFeHEb�y���[	���|X���#8����O�~��ܳE�~Yp$gY���QR>^��
Vˋt�\����pc
ٹ�8��Y�2���kqlD a4L��IU��B�� �a��];�"ʧ�[�s{/�2�!ݮ� �Yǚ4q�߃O���=�{��l=p
"+x��L �_4�t�'�s�Tް����/��^��}�/E�R�T�7uK��K�/����2NY��Y�$:�$� �l��z��G������^���:rC��P�	�)-x���@��w�̂�����vg�r�Ѕ7�=�|XsL��F� �qY7��@<�iBd��@76�5@�G���f������� ɽaR�,����p��H�� :��%�W#�CN�<�İ(�ڡHR���Ͻ��I)#�3t��7d�"�4��N�;c�f
Wb��:8��`�h������\I�}�g1������'n)�o��;^�d�ƥ�9u��
�I}�z�9B�G?�i҈P��5��8|>�mp늦����@��R��~�:^����-����P�R�5W�jQFq�k���ꖻ�x��Xw��Z�L�k��2�t5d#���Q!&�VOU� <N��X�V��I����RM��n�J����:Í�������raCj�N)�h٭@�P�u�"Z7�J+��=as}A4���o�~�R��r�e�=&8�}� ��O�w~5�:���6��2I֫�V=E�$=xaR;_�v���Й��0Z� HU������*
+���7n�9k��ƣ�d�1����䑫m�+,�I'�
�'��tV&<`��]�GX<��̇��`�J��6@�	s�:{І�Q�&~�Mwz�5�u�Y�
hP��E_dЂ�Ȱ�����[\p�m��_bHX�0���G�#Ǻ��?�a,�-_���PùӃ�YK��j���H�@����/� 
$�Lk�W隢��S�n�=Sz�׆�M�i�B����r�ZR'��켢�?�z{a}"{�B��j�%�\��#%�Q3��{�HQD��v�b�N���jT�AG@����L��IB�%C҆y�Ô?��1/��{����"�K�M&��������ְ!G��lOʸP]�0�r�� ������t��K�3�7f�om@����*�bͺ��
�6��/�a�"��`���nX2ks?����(�Uz�=�u����uay�.�����ÄL��2"�o෩^Ș.�y���OS�]c�s��"Sƨ�/xJuQ�,��q��j��ζ��@��l�E�1��oI������?O.��q#ܑFA�x��p���W�͏h����4ud�c�W�w�]֏P*�P���f���.pu�9�s'�?5vSvC�E*���,��d>�,[N%F�V<�O��H�r��ߢ��ܑ鑙n1���V���t�sv�qA���]���ʠ��ѥ	_���ݏ��7*��ƣ�4��n[R0�\�Ľ��}
ue�D�;�[x��$��
�PMΘ�0>oo^�*��ғ����b����H������Pi� �}]�I�T�*³�Ģ	�w=�}xS)�Լ��8����ؖ�x?0�� p2ǵ��
{,��h�e����'�>���줃[1���UCݜ�Pr˸��	Ú��h��@G\�K�_�u��E�kCVG,��|.D�DsyW6����F�9��*k�]D�e��sJa��@�'n\=1���"�&i�2��?�f�)ڨVc��?��,a��XG��sC�t��t�
Wz6p]k���m�~����B��
�C������Z!i̽=-B�!��qʍf��O�%�MKA:�A��hn+'�bP�:v������9��j�_�W{�h��%����[l0��>�l'O�J_� ��#��d�^Frٽ L�V�5�X/������	���8w���\�F�"Ոa6���s�a��l��^~t>Rk��X����7��m���/�Uf)J�
L�ۄ�5�'i�����g(�o�4�����_p���
�����I)��O�Wt��	�d*+��nts��������V|׍�(ab�xv��%1�l����A�����W��!��!&͘���g?�k�:��5l1^_��r�z��S�7��_�Ħ���޶��Z(�YYW2�ZM�
��'��w8ˌҷ9>����	������M{��M_���#-\ǉ��j�+�;�M(X�}F��������K~pF�g=ā�V^*��ހ�V����8��Itv]�
�� "߿{�VE��nՃ��sn�b�9K@�p{�e�oB}����ǽ�X*vqhG�'f���Z�	�d��9YU�\�9����|t�` ۙ���E�8OOSB���}����� Ri~
T�/��ݻ����a�~0�J;�ar��a"�����[�h��'e.����A0Rv�N	������NI#b��Q#�?�9XM���Z����\��߃d��r�ȘMB)��Ld��P$�c	u*E'LBM��Q��ԝ��[;��>��ЬVg�I�l��jCO��H�.��4.ΰ���E"D����JI�	͋EEݾH(�����J�WI�1s��0HB�v 7g@�W��9V����dZv��C��-f��G㮻���&ID����q��t� !��Lӆ�Ƀ�m#�m�<�	�-Z��=4����Ř^?�2J��$�U�2uD�?�j0[%�'��]\1���E��ڢш-�,����+#��u؀��`Ag�<��,l1s�/n�������J�@�:�Q�'�O��~T�9LI����㩸"5�7�
V:I�p����o��m��
̾�ںM�jHcz?�;�����{m��2xgt8��-�DK�Z�=~}5�9TA�� �n�.&��K��vS��8���E��Ƈo Z;��~�����]!%�h�g�w������hq�-e�s$��x(T
�_����f^�{�	���5���02�c�!؁E �����61�$|�ǝ2�&U^��oߣ*�mrY�{����˷���SK�%��T�X��a���#s R��2ǍI��Ε��Nzb��GH
fC��V�k���T�AL	�
���P�{y>B�^[�0�׉_xD殜@!�Õ �|Gr)I�)Б,��d�aDFI�Jm
Q=�Q,��v@8I����주]����|7�H����>B�0�_�xJ�̖����v�d�H�y��Z�~5JGA׀\����S3�#e�!����Yr�c���@k?:�\L7�/���"�x�÷!B)1���|�A"ܜ�د<�����E�U �T�������7������q��=|�(�W��}��JFԨ�T��k�;ҳ�WB���2�	7՟<riI����7�,� ��~n�^5�`�l��],Z9�����l	��l���z'��i�ͯ>�0���!�V�&E��}ߩSI���)Y48L��(v�V[+���D�rj3�˂�Y�mJWI`<���$E�5�!��P��n�QQC�D�njBO�O�s�7�;w�����A9[�����8N�2��0Fd��<K��ǒJUx �.��D&�`�'|1�c.�AR^��O�X󫷸���3s�O�~4�/rbŜ�ʫ�y�s͕����b�ۣ]4������j��I�<�=/9ʿ��V�ꓖK�e�n�,�ٞp�Mτ~h�<�L5WK�F�w�x�ߵt�����"Y.
v"9)\�����YL�"�AK��r�!4��Ε�P.3h���B���գz6'�9BR�rM�>�e��$��m�R�ؼ_>�mVF���nZ-Y���K�yՀQ�q���R=-���X� xfZ��� ?[i�XM	cL���%���oخ���9	������c�e^`tOh (�H3y�ڰ�ư�� ����T��"p%���}I#y`%�}��ObYY�n�uU���3�3'�,�#l۵�o��i�>tl�JWz�Q$
݋�
#�Pj�4�׋7f�R#���A6m���#uo�Q�d1��[[��~[�Ɂ�����<�&%`���7�Sh'I�����lI�#�"u�B-�A'
*�[[B-�l�Y=����+�x����^C��6Y�,q�3�#�`�Q�&�Ԁ������/z�M04գ�U�MM�F�d�B+q�.��ܣ_���#�<,���L<\U�voh��kG
qY��v��9�@K��&�W�b��j»��M�R�0��m����fu��r��#�<t�(W��~7�r�h	������U���|^�F1&F�>����6	0�uJ Qd-����!^���y�9�X���n�����~��e,�O�����Mm���l��#��)��y(]+��q�B�ŕ�3�Z��F��
�CT��Ћ�wj�I�`�^;!�])���!��L�'�9�kp�0ՍJ�F�Z����P��^ߎoXX�>.!�Kdg�7�R�wl�����K!��oh�|D��`���_<E�L��H���l���h��fXҦ�=`u|��!g�10�+S�3vpR��+Q_"����"��1�*B��4�P��[6j/*�82��d�����6�N�d�F��0���Z�+����;'��h㣨>\Gع�ٍ�L�s�d�eEzz�7���t�ϔ��H���ԑ��4�P��5[�^�_@x~&���8"��q�����Ⴟ}�3�;U�m�ܭCGn�?b�ِ�[+�|MJ*�R���E0Ljo�E���$���wEq ��B���0%�S�Tby�v��T�m��X4� 3�I���ύކ�h�_3�$�0�b:scﻎ5�_����R�O	x��$e�6�ӟ�G�c�=.�z8��~�&��%noCz�a�;�*���P^�!��;���
/����~�#�˯��΅�T��5%�N�cm��&���g�1��Z&��Mc��26���!<�6aL���l�h�^���Y*K�6�y�LR����A�7�ݶy�?p��k���ʔ�uV�o2]/}���b��.p�@������2�n��Vj��l��R���f�9I�Pcb���&dB��4W�_8��ެC�G����6}�c녛i�8��h�2JY7��
�/^]��̹pߢÑ+G��ɗV�=(y%<߄�LuŐ��Z\Р}�ѐGP��1��+�z�wK�q���
۽,,�V�+G�/��wCu���y�A\ts�OiP$C�ǙOq�&�$-\nIї�-����[�+�B%#|�~���"B�\L�xf��{����c���X�7�_W�m�\�4%﷊0�zPw�l�������=� �i��qda�H����[WO�!1�w�si�4n��zoʮ݌Ƽ�����8Iő� �.��혈K=��ɵ��v������o[�8��f��P�}����L����H5�>*������4����gk�)�L���wny�"w>I�&�xޯ�/CL"N�OgS��.:�C���u֕�����?���[�7)z,GA���v��%3�:��_�?& ���TKMOn�S�T$~8�=���d�<1*8���FeT#IE�r��~�٣\<?��$�����/������d�������\����%|x��aDP�ˊ��������������]7��kHTj�1��C��Ж�֕Ɂ�ͩ�@k�H7,l�ȵ�yTi�9�&��T���ao�\@ژC1v�g�."�`c��tXiF3�qZNe���X b.��,ֲ������c�r�mJ1̸�-^�R���Y6f*U�c����`���cU�>�$�煣0h�PCˣ�|�Ѱ�eB䷗s,]�TIuc`˵⁭���]�����e@+q�.T�d�S��G�C�i�;k'�k���a+��9h�t�JhϦ����2���툘k�������	����p��������
�,���y���Pu�"���k���F�ޙ�����g��=��:��P�B�zpW��������9�j>��W�=%����-��@���$�n������^�����Ԍߦ*����L�_Tq��
�2�2Fv�4�A������r���Ѭ��_^�v��
������P�?o���0֡ej��?��E�e�3�) W�DT�s�P��T�c?q�F�� �L�����-�6%�~��/����D�6�#.߮j���9�K�ͺx�w�B}���ۿ�}L+�T��l���L..bջ�M�j^��A��h�QP�?p�%˜{SP�0Ɣ\�<h�]��ۙi�m��d�XD}Ql�׶3%����6�</ȸ�x����6�%�W�,�����׋[�#��H}Xn�u�}
XLs�̡<���`�M�G��9z���o8��=0�(NRP�	 F�KnT�r^����Zay��M�H\\�W8,��q;� �3��Vt���M\�߽�[<�(��x���2x4
<v�a����9\��:�.Ջ���_�2@���
P��e���lQ{k=��۰1ȡ��0<X[dji$^p�^�A�{(��$OB�hƛ����"��Y�"U���&�>8)=���go���Eb	{{
��1#?=�]UV�D3�E��=�҇�+0.=g�˴P�Z��T�����qG�ɋ��|L'O����Y*�'X��2z�(�c�ؼ�2�샞_��㹕��Pw��e����?v���i�����z�\L��=9	�S�D	���I�%*o.iW/�Rԙ�$�)�p�́Z��
���(�p�q�����9Q���RQ��Zϊ����r]g�C41s�2q5�gX|��Ө�&�D<�!gf2�<T&W�<�;vBx?K�4���}�����I��:c_� ��������Z���Hj���ĹcEG8�	�<4�|dkqe^S����b���9�e��19�!
�9��4/Ub՜�}^4|m�~
�[Y/^��}/(u"%�a�ӌa,v�NF���m�p��%�3�M����7˟�^ӟ<��ң-��.m�.X�]qD�N�V�A�"qO�8��_�������0������z�h��Ѓg�͌t>k��93|VA7�,�uhAϰ��u��2���n���T�lm<!������@Q��W�����'qgH�R$'�/4v�����@�M�ti[��u�n4C=P̑�F��_�B,H�:��wz��<ר������s�����˕�m�-`X���TS0��OG�O,����Ld��̢�g-�Lf�ClR��9�<�Ky+$-i����ԚRj�Q]�Zq2;(٠G!
���Yw5A2qO��~S洫�lq������~�`Rm	ƣ�q̏�h��ܹ�x/A(B��b��G�֘0Zo
�/j(y�.�s�B� X#�?�{�J6�R=��TR���'���Xv��}��)�ퟴNm�:8�pzL��#�����yn�.��?�R�[�7�+$�x�'�^��g�Kav���e͞�<���uG�d�������
�bT��j�wI�����߳z�[��z�K%y����>XS[�dh,�m{^��s��c�<�~/�*{�|��f�$C���;��ȕ�3w#�uH������D����ڨ<q�h���f�g�ʬ03�eU\�M��-�ž*����e������߽eaz\裩D����u�eӇ��EΖ�f	��@����<oM�V��>WG��<��̼`K�v�_h��rDR�Pi�o�x�����,k����m�Z#�#�^F-�-�I�V�No�w��%q'n!@�<���T���-3�-q�'S��
C��1	�p�[VC,J?J;z��Z���-�J#W�V���?�8���B�؇�H�&��Ν��V���䔧x��䨡�P�my˺��0%�2���G З�M��=fi���!�v7�����,���8X#��j�#�����Lv��Z�����"^r���2�/W��5N|ǰ��ޛH�K��U|��oae��S �w���E�Y�)�@���A�Ե�:G�7��\S9r�*Ѡ~�"�"6�ݹ�ٳ������8� �yk�/׌e�3��]F͆1�m�M,0��kFt�R�ֶ�s�~�ܠ�R�ꂿL�h{T�O��)��� �j�\��f��7d)>!�̨$bbhlΉ�릩�R�b�'P�؇�2[&
�:�t�#����f\�UW�j�"�	�`?<�&&��!}9����̶�Z6�*��=PֿG�c�84���i0�H��@I)������#�P�<�����EcJz�s���H����^��Esju�m��+�F��Dz���**�^�6x�s�Tʢ�-z�]͋����l���;�Á&�:+���U�Z��o�s�	ae�{]*x#1~���DR9T��\L���*����I'b�o�)�.Ǭ��~�%a�u�O�n�H����Ӏ�[k
��4� zε�����T�,2���MzȞ!$"����P���	�XF�u�VHS�c����8�V18�T��^�-� lM'��T�ENu��"9p�*�����|uE׈�,�'�z���z~SrsH�$z���n���@� ���t���T+��q��.��<�������"�C;?߅5<��}68�(��x�\"/Hc"�� �F�����]KY��f3{�}���J7�~�����d5�*��>X*(m����/?�o3[����E�p��l�q�[���)�[��
 oKe|�0=U���'+Xxi�x�g�yE�3#�t��^����S2Ey��a�.<�dl�j�
Q��t1���~�!$,U��LY���kٝ��$Rn�hVT�"�D��}�R�n866��!oyy�grP��2�����n���p ��`�tL}��J/b���ĜjP��0��J�1Y\f}��q1�%���o��t�q��U	r�[��h�E!Q��-�,M�dD�bS<�#��K�A�aqt�5�>�9Y���L�V��Ǒ�D�7�N��|��,;$�����>dI|�Q�i@�X�G�@��A�a��E�FX�-�?d�wWt�/6dq��d�J�^P�-0�3,'�$c�8F �t|��É��:\LO��
���I��,�A^�@��i���G�S:#��9�m�F��.�S��?��K�������M(�# y����ٜ-qA`V��ҁ���3��(9jx����8�r(�d�ˢo��n��$.��z�3�B�i���ǼA \�7�:E��mn��l�'T�����*��^l���7>���@��*��	��Ĕ��Q`Ơ�A�맚�z���J*�g?���!0����ɡ��O��iA��S��-��
�\�*�����9��+6�l��0��0��K��*�;MгѤןk�����Iv:g��X��!�f�����/�=�Et'S�P��s��{˒�%
b)^d|�r����xYRS�At�`�t�[�1�g�[�.*ƺ( 2�G%S �ܜu�@�Ēv��^Q����E/�"(�*�Ő�6m�+-����0���5h���v� ����D=��"iT;I�Г���U�2O�$�
ҟ�4%���1tx-�Gi�R��BC������/���m˩Ɣ<�/�=ה�m�f�>Zf�ߟ�7sU9���q8��R	J��Ut|%�`��7��ȘG#p\���p��'?8w�~���K��I�~6�
������5�:�F*�fz�ٚS/٭�r^��'�����nJ0����Q���[`5�Fޫ�!L��Ds��3���z>��?���K:`t����p���ݭ#:f;�\���y%DD�j�P��:�M�\7���}=`������
?���Ǻ�H|/�A}ʷ�s��mm-�����8D����P�Z��y�� s���2ʧ]V]D)���y�L��B�ԟ�F�tԙ׎�k/�K����V�j!�@�~u��$Z�UF"�ଘ��@�4u��jM��&�-q�
��a���#�V� � �k���$��m{�l���;�_����ye@[Vq���c~Y�o�O7�:�&�E�/8�vk�'$���]�/��"y\C� �\��rݫ�'GI����))J��_�a��U<A~BJ7��u;�SO��՛�	p�����(�E�VCW����}������;R�bD��^ݺy�Χ�Eh�;Hׯv1��u'���A8ԽMn�HI5ޙM��5/�^&
k�ܬ�?J~'�,*�W���-J���+s��c�(M�q�>�=���-P[��}i��z�k�g[k�`�4/O�	��KB��=l2m�N�3��"���o^�8�����f����ܾ��X�Rq쌏A��8�,y'�?�Q�UĂ�b�_vq'�Y�9���'e�J�1�R�*��g�f�!:�rtX�n��; ˆwa��>=�~5�}��'�|w;�4Bv h�Ϊ������&Jxm��T��!|�T��h�˞����jY�S>�Y)T_/ț�3ً�f��]n?O?�j�����+���l�T�)e�<W>�R�&��m~@Vg���:'�άtR���H|~���"��q4O�E�n+2D2�e6_�N���+��vOl�]9������O�[]+|tdz�S�X�%�?I{8G�G[�z�k]� ��ڢ�K6�Z iְ�~!�����۝HzK�8���^%�f[�R_�\���ZJ���_,�w�z�L}:�%0v&�d>�q��>g�h'H��Pmxj�a��B�������aS�{�h g+XRn�ex�K4�C�=o�1l8��}�~�:͈��?`�k|6��63&�ق�ƫ���� ��������k�&j+W�Ý+�xo�ۉ��Ĉ�cn��-cG��x��N� 9BP��!C���	�6�W�(�^l�M�Q�Xݜ����I`�JJq���fѴ��q�w�0��`C�^���4.�������Rw���݂G��؂x��IC�L&�"?D�5�|/cYs��ػK�#�g�3��v�i����]H3�l�;�.�r^D-ٝW���� �0�^�2�R�瘮��8�w�=q,Oq���fZ�?y��)B�k$�?xT|D�;��3��9���,��x�1��b?A�d�޸y��T��7����>þ�u?�{�K<ى*�3ܫ\/��	�Lٙ?=�]�~_�;9y����4��D�_���34�0��<o��h���RQ�GV������Lo���na�s�ў�;�O���Y�%�|͛�Ӟ����ǹ���ɵ,��+�����Z���:�-�]cp3g&�>Jǋ�j����ҿ��e�ɆdV����n\l?�MV�p�gG@Ȧ�jN�E���ԯBk�O��/� ��Z"���B���@Xrt��mN���:o�܃��~���q�v�[X�誘��_���+E�W:)K�1t�,�'b�V{w0bX�D�Y��'�1�����0��D8U
I���Ķ�wur���|��W�Mύ����ΕkD��Ӡze`��֞5����P�� �!Z���Qs��'��e�;��{�1i�kr����,%�"��O�)�s��7H���u�Y|�:�,s��?%�Ql���=��=G��9.���]�E!vr��xƕ�b�o��w��H)���k��<�O��;1Z�������7�����^N���>�+��n��og��%��P5�����e�N��g_�S|N�j���Ū��t��+Z���a_�Л.��O�bF�2�%p:R L��V?X}$�@�x�Kt dy����y�CJ��ea�E��9Ui���=��?�L�
���htq�p�Fg��w���vW��/�~���9X=�
�7~�'T%�C��/���s���p�g5JOKK
�MFo��Q;�B"nX�"d4��b6s;U����2�g8�v�t>�"�{������
�^7�8��w��I�B����*�P���s�E��l���"\��d����C��J��@2m��ͦ�4��1����j��l���Rw�6��,�Ac�K���Q�l����d�fS@�2�Յ��t�UF�/�Œ��N��0����F;�ט����a�4��˟n�p��O�S����X9�n>@��%Ɂ��z�G���j)�gk�����\�@�}8'�|� �^5�4l�Q
$S ���p_}Mt�?�9�p�aHfV��1DB�ߞ�7.��v�
8�`��K���w�E��-׈;��N����,��DC��y�Vצ�f� ̑"��9�6�4sCTV��$����Wv��?���GE��ӯ�ܾ�'��~�~�����g���2��؞��g"�)O�!�A;z��j�?0��+�ER�u�uN2�x�[P��p9<��|�I!S&��w�C:��7�OsQ�u���P�u�MJق���5���|nw]�ow��\_.��n�k�� �����ju�*gv��ۉa�-!�מO�ͳh^Ff�/�D�8l�XW-�k�^������?K�p�_��fPU��D�9RODJI��#&J�l<��w
��83͢S�J!Ah1W�b0$iis��!Ko����Z�N]�Y|����Ɉ�͘�쁺J�E�HqDI�����%�ee�f�����Z�n��F��y�^�����7l�jFY�������f�T��J�=�t��w3�����ً*Az�<�w��Ã�_q�sD��e�!UƩ�1�po��篞h<��"T��,�S��d�����_�ף��
�� �B��=�[��ǎ6�f�O7���6�o�3Vj^�����۪ȚX�v���������n���EI���`�/O�uف��k���C�LT�i}�c`�lK%��3�m->���[H�t�^���{Be�WpKz����D�
�M��Mb�c�|q~��Z�f���?��W�ș�i<Pu"����7>���_�<4��(�6v^�a�2;E��vy@}����i� ��!H�"J1��Ƹ�����"�[��K܂�2����8Yn����]z���vwۊ�F����r�"Obo�I�or���}��s�<����)g*ᒬ�Ӱ�2����ٖ�s�R�I"�ĝR\itI��C� ������>�)'�M�u�J�G�6�g���%P���Ww� 7q��g��h�'x^⑔�W�唟��7���PWZae��e��Oҟ1�U͛�6���I��^]pύu���>F��t�4x,t66���r���#�����?��)����"D��Sև#ϳ�oƤ�\��S�Au��v|62V�F�M �8��I1+M+��f�!pn@s�w�1RҮ�{�I��u�b����e�:�I�3+�+�9��~�5��GįI1yCp74�e��=��<l�	�Ѧ��k���5�H���-s�e$j/�8�� CC��������&	IE�[�<٪����qf9D���W�N�V$3\��z) �J?��8&�O}C�Y�JW>S+��'\�b ����{�R_���!�"Ѿ�K#�Æ�eK�����߆wm�q&˽��	�
��(�Y��9	��6�)�E<D��SjSO�.�	Հ����Y� 
��ؗ���I�����O�\�A��ߒy��]T{C�F)�g�>[�k�X$d}�P�:�I�wX�t>��v���Im䏭曔�����S_Z%��Bd7��e�,��T=*1h)����/�������K��%v1b�^K|�w�/?�t��4�������`�~� z]� ղ*��I*�h8���kK�".&��ch7��ee�r��NKv�o��U�8��a���WV��?�{�4��Bo����(�߇o�0�O�KB�#����h,�1�]gAp����ˢՖŅ5����_ZF��[GW1J\�Yz	���a���K<�Ը��i��0TU��-�Iz��Q�|�G����f@K�̄�/��'��)��P{�W�.#R��-2|N�b���bi�&�n�$���A8Kyϩ�$��H���N����=� �w��5�*���_����k�P�|��@F�;f4�_���)9b���D���� 2.��T�uD�V�.i�_�tӸJ��{Қ�
�+4����=.��w�5yO>+YР�<�W7y`4-9�6��gd10�mtt��ʣ��O	���9Fu��m@�$�#��#��?Y��7�e�,T�C{�r���r�	0��-L����DE�HR�H�ܔ��jX��<(O����F�k{�&iL*��Ӻ��y� �ٲ(�U��3c�����O���%_k���Y?������o�R`'�LnKM50�A��2�մ��!N{!|_(���8Űƅ�����R��}�4��JҀMZ���T��2�����w_�T �!��ͭ�Z^�`$(�4ao|y����P��ZD.���'4 #&��9��mW�:�&6�~`?\$�d;(�b�߁��?���E�ýo�_(Y���e�!h�v�|9��)4��v`A����\��n���6<�ڋ�i����I#$�0��f��?��0���ʚ`�KD���#Q ���I����;�;�uJ�	�����٘�.Y����b���P��K�0���O*l�?�UPc,F�H��y��
��⊢�q<��b�<���T�h�E�~�~��ޢ���ٞ�r�3�L�����Y�.ӧa�l���Ϻ�Q�����\o֙Ӭb�h�§V��dS<c\?o)���~��I���p��;��FW��8����p��f�	� ڿ9`���f��|�݅��J�6�=�� �Eyz˶߹�d����S�f{]Z�-W�s��r�n?��Ǽ��Q%f��� ?,g|qMJ����Ruy�U����d�qd�L�w���qA���^"��(���������Y�.H<\�i�����@u�|<^��Z�jB>|�yI� ���=~M!�E�5K�ŌL�J+�ۨg4B�g����M$�郯�?R�XM�9�_���޵�;�Ђ�����h�c���	��ܥ�1�^��:&�Y&%HX �a����5E�%c���sO�����*�Rz�)�~b��r_�h�ʂ>�x�����.K�#��؂��pB#���#���<^Ü��4ӵ>�[�@���$��SL"�
����v���^��n2>�1ҧ��ȖXNb&$��!^���P�i@�2o���'�2�ĕ�:Z�G�����o�ć[9w��/'�T���������w����4v���RCU]��s���g"1&��Wiv�N�����}��oE��M�����\z���y��eP��z,z��|�zkѝ���8���ke��
�\����Y��JX���U�Z�m��Ү/@��q�_���M' �T�M���#��H��+��E�Ñ�M�mk��@	u��j<��l�SU������䭳�$j���c�Ŏ��L��+������}@�Ke˖L�4�S�˘���� %Z���|�����e�!���Yl�*�@5���� ��dd��g�ۓ����ZL��!���a���#5HU�Ȱ�'Y c@�F%���2Q�j=�����_c�D���"~��c*�|J�	��B�!")�O�0!������އ4d��#����먧ާ��HJ���R���2���P�mK21lĈ(�Fv-r��>ĵ��to=�����f��,q� ���L)���V���	�*��V��)�?@C��.���hJ�U�N��;}K�ҏ��J��ZIy��@�階{\9�އ��:�.���9�����`ގ���(��t?�:���J=S+H��L:�wtq�SĮ�k�7��P�KD=ʁ:�G#����!�B$K��9��(�֢&2@����-�(Cxq�1�?˲��9=��u��c��~d)�U߬�F��`,��p�wK����� v6跎�9D78���T:�I�XKo;�v'^��8%�O��7 z���	FzJ�l���y,�O�TT*�i��'E?Eߴ��F}l �����Ak9i@/�?5x������߻��]׆z�6!��<O����B(�J�=<G���c��jM�J5��䋨��H	�A�}c�>��]-��W�nqC��	���i�,'<{X�s��H����
���X�E6�j��!{��&��L@Υ����Ȉ��0��F���&;�m�Ɓ^�C����Bq灩 ��!���B8��=p�m���;������}�^I�E \QfǬ�{�x�-j�i�TX�
��$tEAw���_ ����<Jߎ�K!{����R$�Ux��#���跠��[<
�"�ć�=�u3�n���_/�"Y|3h=�����+	��h��)��`tF�*I���tnmAz��<n᪮w�K�N����
�?R��'�J:B{�LMLw	4��j ����TY<��:������۔�,՘��3yX`���6)j�gr��O�0o�h�?5ie���wK5��Q;s
��A���£��K�~�haJ���/=s���-��Xwn���n�*�s��� �\�/&b9C��ޥ[C�x8מ��.�s��D�g���>�GH����jQV�d`�4���Wr�a�\[*U��09��<'pdk��%_�n��\I�G�驢2�y���u����D"�1{��C.S���Rz@�J����-������症|3Gr�K�`W���B@���p��D4��)m��� �z����/�Z`��A#q���8q#M��Z�L](#�qM"�+Dr3����s]��OO�j7<>��^=��o$Z��Z�����5��
/�VآW~&�]:�QA�aUc�I�˼��&�4�	!\�X��g � r�9rD���{��$x0՟Z���q���_�UwU!I3���a"�7|��VM�Y̲*��pVt�45O�gns�׬3{��G��c	��':TGd�9�kx�e��:o�rT������zYpT��<�tjj
Ǐ\%���Q?���X��/}����Vs�K�o,��l~���r�V`�ѳӸ8j��Orj���Q���Z��t ���w�=��fW����ns❟]��_qD�c��(eŞ���;V�O� �1�;Eᑰ/ /b2��W_F3x�A�.�C�M%�ó�S��|��0Ӽ�L-%��?5�ͅ
��(��zV_Xj�����vIY��o#|Ğ0M�+H�HKÂkԄ����k=y����(Y_���3�K���#P<S�� ��X�O���*��L/����1��o���s���\��?�.:I?_��(�g�������E��-�j33>�|��Z7���nFn?���D��\�m{�����|�p�s���E�Wf��d���R ��M�a&�(��d���n0Jz���.�6VXv�f��
��l:~F2�R�6�9�j����f#��W*�B���9ش� ^{�_z�~��4%�ՙ�����>��3A����m��
�Ӊ���X���m�i�!��hY��_KQ�2�^P� �0FiP7p�� "�É���Xoq##s?��*>ؙ*����X.�77�F�`mt4�}uZ��\���ĩw����v3'@��'ګP}���!��&��7>���A������ۃ��e�a����O4G�6q�f��9j%w�ۘ���s��C�/8	D�&��44��8'�*�r�v�+�+*P�^N�SK�<Or���1A.c�j�e��ym=�r!V�E���6�o�2\rj��Z�a����{M��y=�4�ԤIĥn�i/%��}^�Zm�45����A�W䤞���3�$ƃϻA���uvY�\�,�Kf!����	%Ϩ�cN�>E/�ueځyX,����
���7��H�÷h���j���QH�v�u��c�,��1q����&��j"�u��VhWF��P�]B�ߏfg�eYAq�B���=���E��V/�8��������;fV������"���<�n���{9�p�����ܓ�����N�Q�76:VGF�G1��+�}�4�V2���:Rh�=C�o3C�b��K�}���?p��G�m{�|/�^B�Pg$\�`��U��uI�8��۱����I��b�*0]��k1�,�Ɗ-�(�!��Q&�ⴖ龭]�ꝿ�L1B�DHHbҔ��z��)�
*{W'�S��7��YM~��|v���L)�{�k:�6h�+1�.�b�x(����b�����&��Q]���W�i���dAR8Ѽ�wX¤(�v���s�ן�K�~V��^k߂�!p�	;�6�X���3�a��̇��wܔ �P1�=��6K �)ke��+�Cs����� S!z�\G\P��8�P�l�~;�-�Atd;�&���O�����:�l��U8�}����W!q�9&}殞��JŴ�*aR���3W	6�~IV+�T(t-@��lwGpg��
Cυ47�|�J#*����ͪNO �#�>*���bh��/=1�E�ڕO�շvNp�|�4a����4�v�v����)H<��M�����뷡8r��6=	D����.h���ԗy�xK�������5~��l�U��P��Gg"���4�}�B�����99m0S0��²EV>�([g��3 �:����+�{T�:Yx;�~�1����́^�E��z,^�(v0���E`[��w(�'��]��������^��R�ԯ�+s��n����%�H�:�ő����TA;�6SS'�<�E@t���p��1]�嫚���}�����v ��T��֜�Z�ы�Ň~��Rz�{g(o��r��_?1L�#kA��_2��y�W6�|�����ƏPP�/"�P� ���ȬT���`eS����D[bIB���P��p����.���yI�gEq�y"�{�Z%\�g�������(M�� �"�+`�RD)�o\c1k�gDz�pRa;��B$�2�m��k��˒YP$�i�eӵ�*�Jr%����1�/��H������(pa���gv��%����p��?���;�߹��\5�����	4�ά9^0�J$r~_:�? �m�4��E���lQ4E8O����~���T�)_!t(�|��}�YU�~/$Ԏ�YȤ��ײ���l�2+�%����G����Vԏ�+f'G�T����E���R��eRwg���C�1w.Cf�-�ڟn�;4���i}�5$w�����5�����)� Z���!�,W�WTG��� G���S*l�rO
K22�9��_����ļ��r���Fs�r�_�`�������%�G�w�Q��u �83����X���M�2T���-���3ٔwXxx]@~�sͬK�K?�r�؃��N��a���N�4,�kp.y�N#>�l\�	1U��M��\�g�Y�bt|� Hg=4�
�F��RFro8�1�b0wܪBp��a�m�`���u;������:i�<>���9]����L��kO����ɖ]V�B`2gN=�G��D�n���؛,X2� -�Tڒe�R_�T�8q\L9��`���rM��<\�J�k' WW��c��Y9���'�ux��|�ؑ�jhz3eʁ)>`&���LtKr��Ʈ����]����}�/|6�,�H��F�77��~Z���huFf�o��5��b��c �d�j�__��m���i�*¤ ޚ�pH+�ve��kzG$�0*�Jvzt��� ���&��U���>3���d:���X�sN����v9�0��V^l����L�+�F�.֓5�fb{�*���D�\J**��k(���I��I��(�]��R1ԫ�>[?-!�p�djSϝ��v���d]p�c!W:�E�=G1hG��S�2g�Aj������j�I�T)y����C�v6�	,���V--'�yl��$O$΍�#�>���#%���Hd�w�^�渽Y��
ߪ��k��=��'հ}դXB�z����f����Mr�xc���שּ(��V��5�.�
���^�oм�$�gO����dd��$�S'�p(��� ����v�;�����'��5@�<9®D?�^"�0��C�zmVz�����ܥK���Ǡ��[��H7;"�����F4�NA��5s��xD�sjut��~/�"ؕ꯫߰�9�	���^��L�	��0��	�-]uJ}�Xl�:�7��:�2%�Vێi���;%�dv���.@���Rگ��k�U`-�ձ���݂����W���?�n��&{*6|��Ȏ`��ߚpcȈ\Fv����A�YeE����r�t��ԧot��Q��E�I�C#�%�IS&�3j픹\��%�D��T4P�
��ҫ+Y"���[Ʈ��c�h��y��]���6�kj��o:�`BH<��q�Ӂ�e���_b]�"���[[ ��M+�Q�]��9��'��t�BW:T8\����}oa/B����r�̬Q��k6��U����9�c3�0��[��������mm�����;i�6�/���P�+��E����a�K�!]N�;��jM��UFdc����L z[�Jy�����|4�㔵��T$T[c������qYU/b�H��]"�ԔN�b�U	L&K�+�03j��̲*�0BN�u��5� bcC$Dߢ�V�5�lR���U��p�����y��E����M±%�f����qW���~�f/�@�W~���Bs��8��R����?�`�1P��{0��H-YjK$.
���4�����-�H����M�d�ʂ���ez[�кe�-]��\ΣE�-�߬�~_�DY����e���D5�4�d�D���}w̱�S[�)?h�>�E���`R�5�ҏ�쫵�X��I#��z��X���L�����Q�'W<5�f'�Zr�Α��`p�PfY݇�.�u�4��¡q������hop3(�y(���4�r�&mcd#s4zR-̀� e��./�FIԍ<��?����$&���2�N��`����E剱6��;��\u���zd�ژ�_,�g$gV��v�0;�M(_BEm��C��l��/
<67�xN6�Mˑ�d[�=��˶�H}��|c�b{��RL����������5�o�U�
'G�'\ɚx�҃o��"Ţ�TO��-��'��ى���Ɯ g���MJ8:��%+��_3H��R:sH�	��BO_�o�^3��-ͽ¬}�39�������S~�ɺ�(l��%�$a`����
1`^���**K՝�B����Y%c<��Ε�J5�+�_�9��Ӄ�E�"�(�z����ɶ����N�.���=�|ۇ���]4�H��|H�#�c�B�a:U��!H���XN��g���(�?���-�_��q!ڮ�²�Y�Xϥ}#��yR�3���C��H�`>��Ft=O�=�?���r��&}$� ,x��	W�SUr�̄4�K;_Ψe��vj��H���XD9�[��+'a�E���N���������=8��e�^B��=I����uI���L�Ƞ&{ȹ����+�7H�fD�o���%ٿ�WH�h��B�G,�� iL]�^�U�$��0yD�\zDsH��E�L�h��������:���-GR�0J����v��V|�%>`g7���+�R���~����gs���8��{���O�5.��Tډ
�jgs��;Έ�1��Z�/4�E\��}G���c(pJh�IG�eȇ���B��
�"3�/Q/�����|~e%��BHJ�e��a���t8qSkVg���O�Vn�7�f�6hK�ݎnHD�����{��:�\��a9�M��9����DM{��5u�C�;!��s��~L�d�)�)�E�Kh��c6\@��b?��4��cX��2{'��p�AyRw���3s�8����d\W0�te/�������a�'�n�V���.�]q�h�H�4�,Ζ4�̎���]�v��a&�ojC��"%wN��Xj;d$s��d�yr�拕@t�n�[e�Q���PA3�|�/�XPfI9jͥ�z�4�6�!hoX�O�f�jH����5(�N؝5��{y���6 �)f$�wEr��q��u�R�o_���Ό�bs��RK�i�g��
��N+R<�ZY�~
�LE6��/4~��}�B�Zy��
�/�����F�g���� �>����p
��L~=��r�(`9�1�
*�i�j���fZ��by�{��GWV������$u���x@���U��Ŕ�B;/�_���`t'�f��yc/�Œ�y`�"r��9����`�H�
�_��v�YSP�U�A��9.�bڹA�� �jk�A]C�<=�Ld�Ƿ6���8s���o[ÏU:�E���F�5��2Sk�ف��hwÁ�혿b�Q��򟥰D�9+�.�t�_����A�W�r��r	�nğc8��CIo�����q&o�w7���� M?ռ9��a��N9�����#&NuS��Wg���vUUu��š�)����֢��y���<y�`�S�_�BL4s3�����vg�����l�O�P���N7���0�B]"�4|�����rt�8�@���(�<�4��ǂ�.�X�Pĵ�5�4�-�U�n���}�2��\�A���L��R�!Y�S��l�Q�0��>~i?��-��g�@�$J���į�~��a�Z	:lk�_�_�ᨙ�\�RRkGk� �T���$��4JsWv?�1�ϑS�g��"��σ�)����3���S��sr�s{cD0L?���毳����󣟰�8��[�������kIvY�G-vD;��m��d��+�Oߝ��Go���-��>|YS��J̘ʐ���� $�ȅ���cH���8,�&��{��a��LI�*��O��圢��������×!cq�{���޻�zK�.�I��Ԇ_�V�4�N-�R���یy��g���=�!�߈k���σ��i��1�=��]BT[ȸ
�(JR쁔���o����T>f2q�k��X��q�1X�F�&e	`���� I���K��dݢ;׼�P�v��������B��2�[r�@t�$�.��%ѳ��D��b�H�d�"h[��n1�p�
93.��а�a���)���`�A��7�X�r��/s<y���-��{��gy��m�� ����*��{GtV�g>���%"2�7a#x:䢜L���%'���NA����jNW��b��O��[/���!���٦u���Φ��mN�ݞgu���^Nt�.�d��ٳ�D��P��E(�� (I*f�c:Y�,�h.���w1����~¯�g��.A��Q�W�){9��pC��Σ:[�9`�^�������T����R7�F��f��C��-+
O�X�,���W,��(�"�ژ����X�}f�6�>-zV�c��B��/Q���ߞ1A+[(׉�MM���� Oo9�O��Tٰ�gj�Fg�P�/����L�W�yqx{}�"����,3N�|BdH\q�xUD�t#������*�4�}��om4+?I8�*�R��ZF�j��tz+9�Kdy����mH��
��P$+�d`9�~ǲ�j۱�QT�"5�ޙ��e�T��%�}����ҧĢ�Ogc��O�עFh�����>�=4I�BQ���tu�b��	�$Dȁ+��c6xt
\�� p�^��F��fd�<z�b�y�ޅj�U/��?���U�0��nMgA�8���LuNL�_����>g*��i���v~:[���R�Y���bu�]�U�yQw!c���m�u\��еm��7�F	�)�����!p����K�P��xߖ�1�R����c�Ϙ�N�$��]�l����sIƔL��fc��?��	�_���?���c�l
�0w7��M�-���S�#`~�k�l��s���Ư��c	�������JW@U�s����f�U�����H��t׬�t9�2L0M~�b�ڝ��w�8�z���u���j��6�&�	�9�u�����/��n]M�\�<���[V��&�Ns6ֹ*��P�y��Zh,ж��s=��T����u�>�O��sL]A���k�M�������&%aN�u��x�ї���9^EQ�7`ʎ8�?h�����Xa���_x�n�m?�&� ��5E3~BWR�H�7�,�	��B�"@�n�6�ҟ�~�9T���IB]	�>D$*S{6�P�K|8ћa�^��q*�UT)����:X���x��PB�����WBɸ-���+�'Sa��r�o�`�>��˷������J<�	�Ja�u�E�:/���5)��B�1<*(�-���l���f	�~�%z���[���Z��kEgʔ�u)&cY$��m��#��8^��ݳ߿��R:&�R��D<��IG-S�P �z7�=�C�Tx��O��g�q9Ɠ�%"f��B�Kκ��>��Il흀�������6%˝�~�<���+2 5?K���y������KI `59l6I�9��ZM��̎�;[Y���X����Фd� ��50>��ʻ`��n������ۢ�/�m�����bEh�O��^�"��B��.��O��JoD�.�cN�e�g�G�J�-Xs�1!ϖ������.���.�ލS/=�Bkf�*�F�P�z�iqו}�M�ݫ5|J�9n�Å�n=�e�&o+t�>}$槴�GT"�o��� ��Ƈ~�E��P��\�J���K̛�Ԙw掭Ym���	B��|hR��5V�YN�q�Y�%�"������_8��&U��Jŧ�H����1a��Ym��-�]�)!��=i�	�������Y�� n �_-\%��Cp�;�-0���%��\��,���I�Mx�@[-jq��j��H�>�EXo9�y�v�2�I�^}�a6���5�m;䋷�%)F�i�ػP�=�T;2�L��6y��f`������9�kl<WOYj2��L��C�� HO���W8C�o���WF��aD�n�o���7����9 7䢰0��UpZ`���Q������^}�?�/n��QH���6�,�8�v��5�C�29�m�QYA�������ʢ��KH�4��rm�'ƺm��4b���҃�}R�8(n@g,��Ӷ<�"�$�F�59��miM^����=Z��U�ç��V������1�䥀�(MJ߭�r��VK ����l|������BSQr���7�(���c���2L�IℱN/]M�m#����W�J��B�ߟ��z�m��f�d�~;�G�3�X�@�P~4����tێ�8�V�Dad!.���x����ѯ�~���� O<NAn�Jpmw�@�wF̊=�vzAZ��b.����[#j��Ta�(��&Y�Ɇt=)Ȯ/�@���ëE�a���Rb�t��J��orW�tf���� ����#!����)[ؽ������9:jͫsMUa,i���V�0��{�'Z��� �2���p7e͎=��B U$D}"}\�ߛ�YV��̎�It����7�L���f�R�c9-q��גF�|Z�v��OǬ��� d��am�k��Y$�|�vK��f�Q��N!Z�[�)pPҀ��]1�&R&j����6�ǲ�[��(B��x��n����\Pzd��%�Ǖ��DL+?�&�o����EBm��!k�?l�iI@�eCA�hM�.�;�,�	�0�:�~J"-��OD�P}F�!f9_��x<��_�ϸ)��%��6t�g�b(A#SP�q�-�����-{cA�}��C"tp�̍���4�<C��1ZW��U�c5�J|���: M�A"�$��-�F���}�6�-�����ۡ�PB����/8hrQ�g�fРA9�྘�l�J4C�yNG�4Y�� �4��jsz����7:�t�a��(��,�6ֽ�uh��&��=`uj�6�￉؜f�mp��L��T!�g4b'~�M�S�Œe��5�������  �d<�DjG��DڤB��C�<Rw"Χc�Ϯ��Iȗ����%�y��[6f���ٸ
��ZQ$�s�J�
iܔ��� �ȼF+g�	|vN��>:���]kW��N{c��I��jՎZ��5��{����aJ����-4/'=�uAMm�^�A?����#[����צ�o-I��\K�K��-V���۷��a�n ���^O{��W@���ħ��-��6 �	�Y+�;XB��dA�r��K�L�$:_X��ied��t�5���Z��9��^E@�>Y�G���PӴ���ƷV$�<�3�H(�`��oI&�9���)�0;�� �-:4XQ�JJ���Q�5E����q�0���牂zy�mU~�c�9��}�r�l(���1�)Pg�'K�oa��O{�r��^�YkB&�
4#^}�;`E��l�#m|E`�9A��?e��c�v��,��\5․��y�A��N<�
��SB�\��R��G����^H ~rq�r�e��v��%�E�X�ŇTڜ����(�#�u�)�r�F�N�����||�C1�?�@�>\���Pu�s9��8cY\S{Y���In0���*Ja���@�$Bc�A 5Gj5.OI�`q7u�X=�5��:R$nK{=d�% #d�n̢�3c&!A	0���9�dt=�!P�	��o�J� Ϸ��L^d�����2 ���kD���jb�	@��ɤ�ؑ?��]ȇ�8Tޟ,j|6\�E��8�PY���>7��p��Z��B��d�ĩ�أ��e�0����M�(��r/�;���5#��m�$���SC�o��P��s�L��!���zf�1#�x� �(�
!v�pA+�������z��_��?п,�0`�)Ylu�zL
�A��G�<��MYEuR~�H�V$�� ����A����y��]���+e�q$d��q=tg��w��2�賞G�^���ǐ� �l�{v�=.X}Ǚn��h2�j#Y��Ŷ�'9v��QH�l�GKK�ji��+����7�(	��`��ٛ���"�w�G�͂��
?<;�
���'�{aԻ
j;��:҅d'33�@��D8�d��Oc*3KI��QD�����R|�˛Ȅ bȤ!�a=N���D�0��e4�͌�3s��NrB�
�\��f�0DL<yUp�Lx����m�ON
&a��������lrª�9/b�
�������DS��+�_8�e�4�!~�;D��b�����cj3!���P��Ӳr5�����
�����]�AK�ܾ����w�l�_~=��%�Ө� �I-��+l�G��7�b�=�C���q
����k��[��2
Y���&@pw�M�uT����26�ɿ����L<�["`��e��7�Ϝ�K�� V�3t4�l��
�^`��k�^�e���0*N��a�E����i��-}zoQ��I�F�����vZj�v�}��;b`oy��߬cu�u �>���CO�ѵT	���0u�+.{Ӹ�a���ߴ)�ge=½),v���tE(�-�C�
n��L��ş�4�L��#��%$�T���/qS�K'�,�ֱ�23q枠�^�F
>M��&�=v��Z�Nt�Ԕelv�(2�TNx�.��7D��nz\]���Hip�Y�r�%��_(���w6�#9/a���Qw�K2�,5u�nzY��/eԪkb��4�����6�6!�bp(����GF�}hR��P�6C�)s�����j�3�P�J�_h�U�S�s聂w:���0`�fDO���~�D�}�+��+-,���C���	>\�v�� ۏf�&2n�{�Y�6����C��RT��bș5�.�+�M)�sr�F�j��t�&4��� ^߈��B��Y�Vr0aD�͵�����"��p��5��̶�:mW�Ur�����
�3t�bQڌ2�F��H��xJ:����}�)����&��������+A4z�,[�P;�Pe1��a��b�J�}y62�{ V��¥��K�O״r������0�ԠA�*C���j��4�Kc���hqkH���:�?�m�E3��%�(�c��+]�o�!h��n�M��xD��g�B��`#�-
���Ϛ���j��+���Jnj���c{M炈n����\�cw1�H�%��2���G��2@G�md2��O��%�d�z���L�8�ooh�y�"��W3�Im� .˺_���Z���^<&':^��������B��ߥ�W�i�rQo�n�j��^�-1��7dB.�L��}%Ζ�.�6X��)��Y8?|Gٛ��yZ����t�m�ͻН�ls�	��/���r��/)$_��y���=��-.����=FA=��:��J������� �����CS�����w�:��6����o�z�n�h��!�t��3l��l;�}���������of��v���t��	�E9ʞ��ZĲӄ<�]�\�8r`31Nq���H��O�d׃�\|���!�Z�QR1��� oN�]���dG�h���$Pr�AA� 	��;qI�]ؽ���&���F��Z��)zt����RU5�nm�Eɪi[�:�KF�,�0<ǾP�{�v�_
ss�(?�BC9�E�pdz:x�e��	�*���A�H*j<0���	Z+���8(�I� ڌ0��E�d��keK�^˪^��n�:7L�\�/��R����u���{�HYv����Y�Z{���g�b�ȕ{�Tb��׽͠gE@�|9	��?x��)�7,O%g�)��}��h�`�Q��.��1��+�}��{W�d� YDy*�ġ#�#tb�&+��F��w1V��6�& %ɢ���ޞ�טl�� �]��1��� 1_����
(ft�X�ܯ��KΛ���cfP#�,N5%�9iF���[l@;WH���y
��K��H�y��v���<�ں��6���4�����{^U�e���������zp�#�%�v�-ed0M3)�S�Snb[��g��Zm�6ޱ/=V����s#CS�a�]��~�j-���t�}�:�v���*{���x��xN�_���a
:]���GO���?�ѭSqv�'������O���ڛqh���o���Yo)c�,El��8��U��d
����]�͙�6b�Gy�d:�sU�;�e��1j`c2Gߪm[�j�#p�+�Ɇ�DK�Pg��/��/������}^�����L�+����I}�p�S���4l�E���c=��D}��:8��Qg����	��[�;��y�CB-��%�5�0�pV��d��84a�툃���2:�r�k��N0U�?@�B�]a^�	?5���=�7���{m�-F�y,��WH�ά�)�� l��L��J�#�YJ~B�a�v�G��9�@5N?�@!�\*��z�ĐOĿʦ�<�*{hI��+��8��h�Y)��]�ۧ��dO�3ӳ�+���4tsXW�ȉ7"Kz�d�Rx�h׋dx���A���,(r��h���������Հ5���]���e9_��_u�!�I\���
���2��x�Corj��=On��?�u�+	�k�*�`�U�ې�o{��Xn�j�1�*#�o�����y� �n��BUF��<{�5i���fg� �)�g�G<�/i�^�)|!E�r�q��%��cb0��yqr�6�Z�j�+r�N��p͍���zbm+�R*�@��1<7 ���&~B�a�����fGX�/�
O�U������ޒ�p��i�$�-U6�~,&�D^���X1a��74�}Z�:G�e�z��~���J�8E80{Ί�K��K.4{N�͌�f�d����v��g���eu[����J�j&�ȁ?�P���ݜfj���5�h�G
�A!�!�v 7�/�5!X\�T�����v�&�"�ͨ�=���QI��3q��j��� OI�a;!C����R� �����r�P���J�1��^�M�qm�$ײ7y���e�#�$�fM����"#��Rqc�j��������3R�DY9L��%%#�x�¹�v������}a��ȗh|�t��3�?��JC�\`�Yuw�jW���U��/��an��6u��Q[M���R��f�o�8H�K�5.��~�Ql�t��jXo+���=c7��t	�Ϲ�ng��7d�b�7��~ty!-j>ux�>ϸ��H �b�&��%�`w�fV�(5��#�9����;]�!�L���͒��+����^o|=��i0��$\������֪�~�)���JŖ4��Rc�i� �>��U�*������7�m	:�95sW�.d0��5k�w?Ke�!���H�'.�j�@��$�[m؃=B֜z�������V=�`����k�9b�g�W�T��� ��xl�p(p�tB�&O?v=Gެ�2O���w�EJ�~/�\R�^�=�`z�3:	��p��Ž�B=�K�i����ĩf��������y[��kg�v$+<������{RH�&��y�G��e+ �/'��wR�6t�ʻ�Y��ؙ\��9u�6�:���XI�a���o7k��ڪ����'׳a��.�^��B���O&�����Кw��51�H�$*)|�O�������(�̑*��Ƽ�5�𩂟�d���-ڡpl^'�}*�����"R<n��Y䯎yV�+�F�xQ�G��Y�&������t�^�҆�0��^�PR����P�7��1�Yg �2�����8G��,������(Ƕ{��Ʈ��= ���,�W�Re�EG�+`��ZP��O:��ZBzj�?#����~_Mnu����垝Kބ������m��TĤY��J��cdTd�2����R2��{��-n-Z;�8�3__�~&����S�^y����8w���?���~{j����	#��L��s���3_��; d������P��@N��\�����5��ޥL��.�Q���!���a��[�:+��j��=@��AL�`ʐ�`� �U)�����cyq"�.ي=��VP٥���3��#�E�3J�}E>ړ%?L[�/ڒ��1����n��!��i�:�jq���glv�B��؟N�*:��6� �h#���O�.}@�����#�"/˖��1�.��p��D͂n`вj�!@��ںR���ծ�| ��RP#�*w��Y�����X�؆�ހ�x8���0Ή�1i�T���|"�ptKBY֚$������w[�|A#�ѳs>H�gX�$�%��4:�~Q�~�������)؜������J�r���>����Ct���XNF��F�2�,��(v��Z���]l�O�ʬ�����5���v��Ӕ�F[�ztr4�f~�$b;�b�	�v�S����e�@���ߤ��x�*w��PBC|�������]��2�̅��A����x��KX0a�u8-FhH���Ё�a"m�Y�]ȶ�[qI�<������y�f����&����~��!f�~�f��$���R�%.![�kCV���P)x�n,�B��S�����,�.�W����L�5���%��4��D�7��v���u�ݻ"X��'�i��f!��i����VĝK@5���a%����l���3
9�]�p�]�&�x�B��3/�����r��nsB�}V�E;W���>HB�g�H�T	�]�9T��h����F���1ѝX1��3�Ed	=ջ�ޏx��@m���3�ɳ<X�ֆ�K��'�Bw�{�h�b\����λ �N��6�s}Y H��)�!��y��z>�G9jkz5� ;1_^P!��YC� T�4W�/�Z�7!v\�Rի��y��ڷ�p����>2�f��hu�œ��Щ�9���D��sS����@[[��_k�f-2)�XM�}��Î��}U��xw��3�YN�\&H\��4���I���2}���G�g	'�O���J���$�l�D��x�T��X�^�8�ŭU:2�^
��>3�����w�⏋JH��_�k7��f� Frk-~Ŭ����^�d ��i_{�+M�FǬ���WA���jN̢�3t۞J�:�j���eY���?��sQ!�uWۨ�4 � %�o�H�h?��EP�'_�7�ѝ��r�x{����B+#��C�7�u}����O+����W��Iu�?e
�	_�׸�L�koD{�mH�D�A���@{*ڭ��4f�dq��@�%�G�+e��C�����9����9^��zJ��*Dc��@6dei�j��@�{�V߃�#�!�g���֚�Ȕ����~�G���L�z��3�}#e�<�V\n4>�\,Q��Ml�e�y5�4^����G���ť���;g��|KW��zy�rn� ��M����`��Zj���J�ɀ����"4��N�Yc`qF�T��b��C?1�� R�����s>z(����LR�'�Z:f7�:�[ذh(���@P[�@ dt���Jd�ƙD��)���Y�Fp� ��=`���-R�JF��HWrY=�%jl��H��\%q���tY��TDPƺm����K�K���U}uLV�㪪�(��'�����<�����k�t���	��dTo� j#�����끊��~0�%���5�D��6-NR�nQN^Ϗy��\[�t��PVC �BnDXS5�x:� T�h��v��@�#XZ89?|,��4 s�:[�����)���Ubip�����TO� :5א�/.��]u�_y�G_J��d���V���W�|�Ȣ�O�ɣ�:#K��8׶E�S�2���r��ҍN��U�G,�[܀Б��= O#�"m�sl�|�k)��@��O!�����!��2�[i2��^�8�l=���j�%f>j���ƣ��yI������8<��vnO�a���d��`00��p"�.�7#�=,C�P��DJ�<{��äg��8��C�^��Rkb��%!�y�!<!+N�2[γnU����2��ѣ���:]�<���V�n�i�J8!AQP���~By��<�mh�=��Pa�M���@��⇓�"��Չ;K�����)&~#�'��"��ђ�n��",}s��;��2�Sʢ_u3xm�p@Nn���8b�CQ�9cn�X��IB|�Bw"9,Cbt[@�U[2�C��V��.��\)�抋�U*���2��3�iB�s�x"�/x��m,a���Z�|���:�k��?h�ȴ�I{8h2L f<N��(���`m��Ց�F�w�����W��OX��R��'O!�ږ�}��npS|/�t��H~�����DEc�k|X��*����57����ϲ���ˍ
��R��(���/s�u/���h�?�Xk�+����2j��W���(��0�R��U��lKi�6�i�;�M%h��s�����'����!�d��P����x�0d���
��Ǧ>)Ȗ�\B����`�޽���Bi���7�Te\��**u�-�FF�9@�E�"ȥ+�`#Iw��;�D��Ǆ�w���V���CV��)�q�9�V��D�H��:�%�����dD��@�W�Kg]�h���a�!4����In�b�`����*���ڶ8yw$,�K�4ù�
X��L����*��J�)����J�㬬2��d����rm�4pkuP2$�V%��lƨ\d��OwIo�k�#�ڴI����(ua���0fq���� X�\ۤ��?���cI{bEo^Ի�6'DSov�n��VR5(��O����3�K�����o�FN
Mɻ��<f��^2��l2���q�U��F��G}�'?�4�Q�[��r	yFL3��0���8�|4�^c���IH{�z��\��B����1 @�q�-"�����CSLǈAA�3�����~�C���U�b�c\�{�I+�	�B���eO6:V�@�3`�������`a1��Mn�i�릙1԰ys�+�ҫw_��X��M��1PC���:���*S��(�J����T������\7>��e.�V��ϭ����3U�
z;ʼ%\95-�ͨ'd���+E)���<�_p�n�H��}I�ɰʘ=|���x�.A�[�7B�`�^z�ZD��^r�'ڣ���r˂�W$��*���5��CiVFX��cHb+ߔ�K�{3T��rШŧ�t�,R@Ifk��<ͭ=�Z�룩�vx�m&U�u>���c���K��;�����k	��'�#��y��Pv
�Z��&5���1�U]�Em�GoQ�� ���7ղ4�����;���mК�%,�R��BC��c]όJ-8�B��}�A�x�N�)d:����〧?6�Y+фX��=w�!甜���xs�����JǛc|�ɸ��"�ơ��!���j�@ݘ�s��W���������SǱ�]�� �G������zUNuY�a$��Gpp]W�z��!�\q��!+������(T�3�r���[�^�"-�U>'�V��A�TJ��B�E���=#�ބ�k�p�o�҆����2.�zV�	��6�2|�;!��$�Zp=�i��;���6�rN���q^ �����'���T�D���[V@Bhקr��n�ޕڋ�զh��haV^�M�Ei��t2c�x���Q���x]���i�<O��/��5�]��{�D���J1���[�<�>E5�|���11)M}�ƈ_�e��c�]�%��N�;£�Q��#�Y���O0M%�e���4����R82t��coC��$|������,g��s�����S{䩔�}�-��>"����%`���]D����!T��l���q����)r�[�A̐�}<���� bW���8���Ba��+ƀ^�6�oU�M��ZtB�r;Roю�ӻڞ�ʈT��$h��-J���k�꛻ڦ�!���.?� ˦��g��������z��ەn\q��r�4E4k~��=���R<�ߍj�ͮ�ki�ǣ�Z�^��g������JR!�I������q�qحiRb�_{9dd�F���\�������){�Uط� #1�`.�]��"Ԋk�<���` ����c�8W~�腾$����' �%�(�-�`�)S��L&�JXV��͐c���!ZF��t$F��_�RЛT̲��\��f]��S/�y�V��Xh
j6�S���Ťz&E߻��8�?N^(��/&Q�![�gV��S��p�_�ӽX�����;�t���.	��eP��G��U�󫕄�KX���!�.� �� �!i�=a'2�G�GI�[�i]FY�����GiS5�~�
Ԓ䁅u����x_����IHj��y�8�]���kB���chc \��L'Q߸�h�qB����l��0��*�t���M��	]jS�`�Q(�0B����EE���U*J�59�|\6LGYy'�&�
��C�S�'먶���D��/~�A�vf����Qͬ��>f��+r��J-�v��#��Y�`�n���a�M-�Io�%3���3wAH���x�tvh�e���tYl�Q�����Y5�ϙ_�^�����t7�"F�f@���|�цUP(��b/)Ċw�ZAiNk>�M��$5	H���<$�N|��0^�ʏϴ�v'"�>�ɋ�j�Ԯ�2�?]ա}er�=�U�M��z�(��%�n!��X;�{%�9���B�D~ԫ69����A!�����L��+WxV��,��"���[�8ɜ��"��)�;�Y�hT+p;�#�����u���(��O}9	%���ڂm�$��P�5)̡\6���#��i�����˝͛�M�TCV�_���&�u�����B�``��6`�L�C���ܦ�z�;�Ț-�4���/�����r�O��������x��*�cLn�r���f?�!�%3=�qB�)o���@l_[(�Y�k|	%�RKP����J�7I�s��?I�
Jcjo���e�iF�]�;��l��t��t��j���h�\�{��o�J{8�zf��r�����\8S�K�>J8�|�ZF�������챊hf;wD�j*XTz�wD�/����n2���F(ˬw���C�$D旟�$"P�3ZGfυ�ɇy���0L'1<��'�c{�'��Jr�ȗ�� �&�A��"¼��ZJ�dE}S���E�����d�a���X�C<�L�a�r:g�5f��������b0��G��j��Z�07�|a�M��U�XW��U��9�>��G�֊>�����ߧb��:�?ts1/��OI��(�Vf��h�ŚQ>9TPKr#4�K�.����gb}D������I��_�N��7��w��i����6�=��Q�ǖbl�m�t��<��I�p�\4�N�"ŭ�rs:��6�XQ�TTs���"FA%���@�����Z���m��_�F�rT4?�1��� z��^7�lZ�+�߭�f�A{R䱚�(Ѯ��9Dee��bsQD�<Ϥ�-����z3i�p�oE���G>P�� p��/����t�ſ�}���|N�2L-�\�z-#�"�!<4�X���uA�p���$ܪ��K�XŨ�C�@J�4�o��J�m���,C�z�/t�#����0�޳fU�$z�<֦�[۰)�[&��7�C��~f*c�!���������1��s6�ʧ1y���8��Q�� 6"��.{6���)X7"7�ưO�V�B�,K�H�J:@�廳�A�U`�h�uu��&�R�\s� ZM���[_��xHZS�\k�����d��48\H]�W4irY�����|d,�ě��MNGB�v�h��]�t�el�D)�Y�9 ȑ�ܞ�dJl�U 8���,�4�r�:[-�t�ф�ӹwY YB�������D�Z�}b]i�!� z:�శg�C&���m0�T���{v�ڋ �Dlz��<�q��#'D8�ú��j�q2[��Y
/����'@N��8��P�P�����+CgI�I���C��~����) ���`�z�$w|�$ԉޣY]�t�:b葼����5�?��5/�GS��w�淔�~'E֖���n\��N
7�4��=@D��f�_ə���Z��`H)��@/��z�V����<����ٳ�����Z�� ���9���n!�YŒ�_����0W�!�_h��M&wŏ�=,�`*�l�0���l1�*�+�y@�)�Ð�q	�l�OV�0`"[y���RS�'vN�X�@���|F�k���m���.uL@�͠�^�S�m�*���'���v*�̼Qā���+(F=
�I��Py�;S�Q�q����L�vǝQ�D)B��atL�1NxL�Ǽ��CH���1��re��s�Q}6��ߓIV�їL��v��󱍯N��>��@.�,�g�C�ܟ�=��IbP�z�)W���`�v���� �B��.���"#}���٢]�YO�tfX�"�@����]���v��q#@LE��Yo=m�"�j�������Z8�Ԍ���\�k���:?�<{��-₞�ff�䑥�0+RG��U�_T]P�u<�����yTj��~\.�ܒ�x	��|jR~� JP�q�܋~C�bǂtn��.�u�;�t�mmy�����)��V|����������+��խf���}I�(�j>��(z=�Z�H��T0��vdW���G�gڷ�'���38�g�
��P@���r�)�c�T�`���>�������[�����Y%�]a(%�E��	�*�
�d��,��Q4\���<9i�,HF�F�%�׻���#%Ә��
+s,�9h��|uN�
V���_D�����l�4�M��a҆�[�nP��>zB�"2�]��b~.��T�@0��RbsF�.4oA��]��*0��`�B��h)x�0-��	�?f_��O��L�U	�*�X}��Ip�CK"1�Ǧ��t��y��ԧ��+zl{�0�r��8��j�b}P�5YyƤ�F���ޑm/��& W�|&c$~�> ��t3�4>a ̀������[!�����UF��ۚ�F��G3Bqm�X�I�R����/���|��η���),�l�HF�ӳU�K�@�R�	�O�F�o_�XNӔq�-q��V�Rv�M9�e����3������{�]��S?���o�Ē��^DR��OMdd�D|7V���T�\���J.=ߵS`+��@�<s��B�I��D�XC�bЫ��-��,���p�$	�_�	���Nxg�yw[k!,�1��0"�԰�&�{��� ��x�@$p�P����,�+k�l��9��c��w�C��zZ�oÿ���.����}�"�erT5L$?��� ����*I�̧��[Q��҅���ā���'�<�('���݃��K��R�h�SKH��&��&�X����%TT
�s����LJ��i����K�[{X%�Z�=hl��\���Qs*�8&�p�k�2�$G2{'@���P�z'�=L*�Y0WkV�L7��\e�_�$3@��ُ������G�Х���0D�I��M�Ya_�J;u��u�b1�O<��=�����}�+�`������i��/��+�C
ܺ뿖bN;���)��p��I�i ��&�n��ǴJǛ����oK�����"'"���)�}�4x�/��c����q�,�(S���R�$���8�Bt��QԨ�1�^�B"��C��?028h��l�b�g�ϔ]��Q�k+�A���z%��++������*�Ӝig�?kNC�DR�A�냒��d=Æ`�ri�"X%� �4�� �l�n�n���s`[�5�X����f̠-|���Y�w��o koFuʔ�8�s0��ď��C�.hgB��4s��躜� H<F� 1C\<��7��εf� l�x�&�K�؀')"Efg�3 �l��ؒ�a��&R��I9*A�!��]4��
�1�f%㵰�r���l�pY��~'Q��k����z�����?:\ %�D���Gсk�`�,�d7[�Z8�n�p@]��qc�Sϱ�\[�2U�.Ǧ����w �f��F��qh���_w�����.G/�M~F���*5#�ݴ��w�-:�wU��ŕ4��SDे_����g����䆸�f!�A���L`��.<���~�t��ST��1Y�8F�#�T���صw�~M����f�[�a/ M�۷�{椆�/��n��-��������L���TZҚ=5��_8n���`{p�ik�
�/��L�9䐼It۽4�9��P��&��K�s#��t!2P�"ѥ@*��8d!ce�H���{9��<T��љ��|Z(���v�&���W�
�d�~���pgV�'O�� @�*���ږw4_��޾�::�y��b�ϹU%���Uc��㵤Γ1p�$�s�g�#����R;^����DO$H�*�	���g�|R4<s���g\��s�|{.B��\Re�xLQY;�W�[V�}p�A�7J��].�Bu��^�#hr}��6H'��~�]�`i�;�J�:����Et��I?���D�ѽ�y��M����i�:Q�/Hd�9�-��i�x�nM�*�����_�{�:�!#A�߄��F����+��pؗ��c��I��m�t��㶜�'F�j�l�^�j؎n�unF�+��?�NB��]�#��l��QILd�f�3��Қ=��3�E��|3���?���������Q���C�Y[��`�/��_[�2�u4 �6(ՙ6Ⱦ�⑿��"K������|n�m$�jz.��Om{ٷ ��,�Fְ����R��9"~�>�$	��W�ng,yB��ɉ�[��O-y�X�.�A!�?*N��m�t}^*ܠ�}�;�3�6�� ��\�Ċ3�B�ݡG$�B��*+D]*$�붬�^<]�� z=����7&���g4�#:�=K�:Iϟ����H�:�w�~�<���	�W�_Hz9)�����UD�8_�M�d��~�?@#�2���E�h���O��Pul�ݍ���j���>:3���t�{6���3d���EC�2��KL�yL�{D���>�\��1vӋ�~���-XBv�8��Z;g��s��(���)>�M���QG3���h�t�0LD��1��`��cz��4��hY.dK�/�3G��e�_OV���9����Q~E�s���T�ܑh�:�+�e���0YrNs]Z��o1�ŏQS�EA������|��7��E(if�׮lNƧ�߷���NΕ�.������a��g�U�ʠ��I�v��I D~��Q<}�OY(4kg*�]I�a}J�f���_���LbL=�o`Oi����ݖ]E{k =v�+z;�o:H��Y� ���;��g&�^AD(���@"��^�lN��E��~S�����[E���~m�2U��I���T�Q#U`P����
~R�4���jz��V7m0$���_5���YlYF�Kc��]�W�d��#K,�$�L��F��i�h�g��L���WRE&GT�����l�ѥ�F�#7����ވ����Q����0�/�:m��բ,0��>�+7N�!�j<�X�L�$�����w���������Ca��_�i�d��ãG�R�/w�+~T~:e~��=�y�2nl;5�Ҽ ���|�� �A�����y����i'����@e�!cj�V�����	f
Z��������L��%��������oN�A��F���"P��:d�=�X?䩭���β�Gn�8�v?6��C�Z��|���IL�.�|f��eK�?'"�ٽ4�!��ק�4�zu!8i��p�@��d��U���DjI'�_����j� ��BJe^N�J�Fs� P�$��a^��i��䲕��)�$�Ik�Q��8����	�����t>���}T4 s��ʷz��&�޾˂m(
���	Yu}�w�a�=�WGsfL��c��5O��B�v���)��N�������y��Ο��3:��E���7 �[=�յ�=+�p\��U͈�J,�rh���!����KR�?��h�l�̈�aCԌ�a�Ʒ�$�	��]����r�%��?���&�8�+,`�g���+x�.hU�����lN����>�$��c1qsG���d���Wc2�C4z�������-v��&1E�r�蘨-���)�Bi���$y�h��x�z�e�#�ǩ���R~Hqn�(�m���ǚ��W�r��O-�\��7$�}Sg)D�,xm[�7D���$V��	�
'���uV�W�9R����V��,yu��$}8-���fT����|Ct��!�ӝ�;&��1E�tV[��	�'��"6�3�M���	�2�f�F�g�.e�M�r��A-<�Bb1+ZG?�'.��u�a
���*��KA�,�$���,"HFg�>�R�E'�uzt��x��ٹ�������;2����rNs�)��hW��+��50�	�=3juz�/�mى�0@Ù߫ �HNs�J��<U�њ�t�����bF�,h��Td�e;�n�+�qo:k%�m��G���v��[�1g��"�BLm��
��8X��7u�t����Kb����|g�X���/zP
 V%Ѕ��]�.Xa1��H���E�i7{(����l8n�	&T��1�h�0$J�,H�@ޙ�m�ou��%�VG�GJ<C���0"���c�ª�I��F��@�t岈f�k����h��j�?Ԩ�y/T����v&��ui�?�{���Y�f�K��W%�)�m��9ؿM��Sf��������p��@)yDB�o��0�לa��T��h>�]C똁%�4�G�t?q5_�/�n���)Q�e	�^c�e���J���X���������� 	��Nq
�,��n����V��ܿ@a������i߀m�`�<b}�￥x��d\������EԘj`��l���p�Pb�^��C�J��g�yO�騆������귐�]����/�e���p���vF��·�[&�EKJ�Ǫ��� Y��&g��Km��3�K����|���"n��hi(-�h��JIۂ����AW���-�b�w|ė~ۄy���_�oث��N��,�?q0�o�R�rw
8�<�-{���o�A,Џ
�z;���������G�q��P8zvT;��X�v�|>�8�Ź�GE�ϣ�(��w%.dq��4,��g�caӯ���!�xXc)y6�8��b�i���s� �ݞ����;I��g�s�&��yR_|���(A�t�U�n'rVh�}7-�EØ8s������tLdK�nȏ�Ρo�e.<��3�!��c���o��'�6DYѷ�����Tyh5!��e�!�j�NӃ+���oA93E�0�1䯱���kpo�Y�t�����Z�u>O��=�ٰ̄����)��z����+܉R�� ������z�L��,eҺj�8�_�r�|��ت��@{G�PkQ��1���ecD�Y�F��H6$���8��	MA�oΔ�_c��d/�� �m�J̺��Sg�w.pb��n����j�^'$\p��ո�Wo���6(��~��L�p�k퉓0N���m
_�hx
�o9p��y���o�ɱ[�bوU�o��y%A�8���i�򟄞H��-�f���`s�d^�6�'�Z��ƶqV���r�[)`���0� �M�/ak�naNĽ�3��Z��SJ.�k��4��Z����^�H`�)r������5�	An��!o��@JÖ��R�dRz�i=%��)���J�MN���h��MG���%X�,�&���*2��7k�Km��,���,�B����[��TT����VRG xE@'�=�P�E��{��|����6�bj�M���-�
��<=��f�w&D�>�lK�A܅~'�KK��c��N���MU��e|������D�����7Շ!j���ַ�>u.�R�V�L^r���0zG-�Wc�"#h�kj.Y5\��J��R53���u1I�+�D/��*�4NOd���P�O/����Vѳ���\��� ��/�ՙqe��Ǩ,��])Jv����O�"��d(˘>y�fp��{��e�!�ȡ�h��TL7��#sc	�.����?���=3ت:�{ev�����������A��8���3
�A�Vp�c���]�R�+����9�B6�>�dj�z�9��m�׍��L3K��A�g�G	��bDY�iE^�v��X::�����w�;D��$�H��,��P.#A�#yE>U��
ϭ���ʡ�-e��vڤp��gs���Ky�v�R~H�����q�T� z��:vR{��r���gb���n�͝�
��>-M�}(��wZ7��)QiV�B�|g�ux;.�_:r�"U1ȳ	��R���)s���j�}��;��A{���o����{y��j�z��Q|�;/�(E��@g�°r1�J���<��7Z�o�/������vƻ`ua!�)����M��7Mw"�Nnv�א��\6����AH���8�9�	��]�(G�؅&����>�����rĭ�f%�S�������V�ǳ��+�J�6�M���1����X�X勞�6��&�r�({�g�@";u}��q��DV��Meи�����r#@q=bc�E� n��e�l"�T��*�Y�E���k��W�M�8|ɰ���F��#c����1�>�n��[3�v��T�OW�`����s�D��P{�x��������`���3أ�B���>3�.��
��g��G�c��t�����v㺜�I���Ry!���[kbW/���&��w(yG,�G��X��F�����B�T��!�/э��پ*�+��F���ݘ�-;�Ӱۀ���]�}����V����;���ڑ(E��HA��l�}�'�,Er�5p3.<���Q�NH�����C�X��گG��n�6_`Ddp�w�ɮ��{D�	Pņ���յ1�ͥ^�O�^�N��D �U���:�d�G��X�b�¡Yڵ�I�����ߍ���B6�b[Cq��A��y(�����V|� ���!�c\&Ҽ0�'Փ�Q�Afͧ���㭥 w�#.a��]�!�F}Qb�ni63��)�1O<?*�n���.(�[p�c�5����H(��|\��,�5ye�P+v?�7E��)�-�n���Ͷ
퐢2Q�*< ��
��Tt5�G]IMo�6���t�"��|(o��e�H�!L���_�b�,>��Ŵ�~m��8�=;��-��L��1�"Ò-������wo%-n�4�B��ņ��j:���Zʱ��b�KӁP��	Yn\O����P?�8����t!ڲ6�y�����#a֥��?��@�����0�w�B6���& ��Rp���E_���@��>�C{���?�I(3��r�	�hw`�q���_ar�i�K���[���.O$��1f��m��#��?�ݒ�&o�YvX]6�9�v�_����څ���kN��17Ԇ�ß�j_�@��S2�̂�[�B�?z�m�S���O'����U(0=�pԼ�.��F�U ��B��UZ]j�دuOY��\鵫�I�i�d<����+D|��'�lI���UR���ub�86�O��E�p�}�J�e���#�΀B�up��f?�7TDI=2G��.8�;��쒪�~�M�踲��./�0��\|�m�/�{W�����>�Ёr����w������U���n���4g<�8�P�Y�4`�Y[�o���b����@|d�c��zF��:�챻Gq���cG���#sR!-苣�v����`9jVjR�S���&�3����3l�!X��hߏ�0� A,�w�w�?BC���qk���T�U�ׄ���J`>Q� n4��)ʟf%�	=�D�
�뿊��i�Z%�b3��ƫIs6Es�w�aZ�����k<?�"��Nͤ�b�H� �h���P)�m�j_+��&Ekߌ
̊o�p7�|� ΀qB��K�<`��ȊXI�*ve6-xr���M��������j���[\S[%����p��d����E-��ٯ�U0�0U}ͨ!1ԛ�b�w�@�H�9��+��ƚf'��W>r�bB�`Mb�w�TC7��ј?$y�/��"M�|e��|��O0f2I��J�z���V�>�q���I#���J3�W��2L�j�W�޹�	�	y�;RẴdWQ�1!B4Y~6�����#���b� U|����8�})ժ(��Z�������X�q}��u�P5l֔Wb��W�C�?�a��It��m|�
�>�k�1�w(͂�ʩ�z�y0���>����O�����pL<Q�kt�T?Qs���?%�5򱻁ħ���]���X͈��;_�����Fl��U��������%�|�koS;�|K���{�}_�	�mv�1�.�5躿����Vԯ������ȉ�O��W�QO!��sY&��0����[j�#�E��k�z  ]��Z�) �������r%����D|[��n��&�t%d�H��0/��p����c�SY*�
�-;���Y��	��}!b��X�1������ ���p��ov7Rʉ�K�nk�ż�2~_{�sZ���[s>�M�h#����;��s���_Df�[�i,dR����sx9�Q_L� � s�	��u�6�+���Yh�\�f-��V��9ga �tp�q�|��>YX*`P�?b�u�R��f�?��(�P�=����6�p�`bO�h�;��*MT 3�� q����o����;zB�f�y���'��(�`��m$Q�]�@A{��D�WE+Ǌ���1�0�� L�@��.��+6�k݃�~�����_�;�Rg<3���[m��Fo��*���}t���^`ԟ)�&QN#vþEi7>��D��̣�L��W�\�.��|����C��@��K~]m�n�~����x��=�B="Ҫ�d��D��W��͙.\0 �z��B��͚��K�����Ĵ�ؖR,B�27iҬ���B���d�%41����0�--��d�b�F�6E~���22�5[Bv�?En#u��z�ݹh,��Q�J7�E%���%C4������vE��Z8��S)l������x,0yEEJ���Z:�@ٰ���I7^�ˠ�_a��M�M4�h����Ep��jh��<:�H==4�?B~��*���J�:�=} �c�r�[��	���H�r�8uߤ�΂	P���"	�e;(��6��aVGu{YFణ�����r��u����0=T���\���p��<C��@oV⟨���]�T��wdxĵ� v�1��r�� �E�hf�$��9l�o�P�CQ%?�F���z���z���;~�bm�1��\���U?i���x�m���}rV��G��{D��*��%N}�Ă4)�>6 f�bc��F��~��H��H�+Ӱ${U!�l�T����g`�]�YS����_��lIQ����$?�*D_��'�l��L�Q��s�����9�O�t٭,.�S�0Z����n��\���;�a��(c����-�-�?�͟���Ǒ��ð��.�Y�%�O@���R��4v?����-�#��	T���c'$G�&@�{�A^X����I�F6S�Yq��~Z� �1Mtͨ�ׅk#BcVi�P%l���[|s�N� �jݑb@� RO*�y�D,s�Az��a�P�ԧ�b�X�'�q_D����^�vg2���K4� �z�'{6nx)m���@��;VN�8��D"�G�'	�x���Ar�W������U
�}N@BѓM�Q�ݾf��e�f�p51#3j��h��Mt��,�
�ƴ���j��_1�/?��.9IYJy ��:X�_'U�D��N�����S���7A�2y�m�b�E+�J�d����\Ҧ����6K��i���	�}��(�˰cV��G*���Ն��c���Nr���Ѧ�kΐÄ޲6��R����,�Z����`&���Qn��H�ü�l�j���k�E��R��vC�^�,��=�$��u�JQ^2���#���������7`���%�j�=�JZ�h]V�FW��Q��+��"���t��ʭEL�5n(�V�5�1ϙ&��55!�qY%���#�e���KT� b!)�EU�3��}�j�����t^3��ժ�z>��> �)P.'�K�r��R׮� hUq����;rY�MM�HQL��Ќ7�w(7�t�l��]�R���uJ17o*�&�{%xvI�-r����4uC;�D-`�*�D�[	U���&m8��J������&��Oq��ۆ��H��Uo��Xzh�Zù�ÑM]�I����+�4��>7i��s�����]���$nO�jȣ�=Ѱ����������b���4���s}˶���������V���,�����1] 3m��O��k$$OLv	'�k�5��m�`��dzە�qL���KzH7d�YӚg"J�7$z�,���VN�4Ճ��g0D]����Sq���zl���s l���L�z˰w)}�,��c��A�9J�K���j�=�Ro	�p��O�	}�S�C�r�3t0���{9�3ZFJ�xy�2N���.���E)٩1`&�ː1",�����9���9mյi"L*�!�<8�)i��O��'Mi��B������~�Qͤ@
�0���aEi�%С�* ��N[��C���8�Gi's�Y��z�e���HX��5k{�k�����x��z�� �[0(���<��탨8���-�6�,����-���e�7�3m&�O#nr��c�Ke.a�
�cZ(4��:����`=0�}q�Ø�NR̫`Z*S���X��P�>s3:�^��P���I�����*��_P�I�E�W�m�ED��]��2(X"��ƕ��)5c��?���b-b�2vߝ�y�H���������\�s��J_<A!d7�h�p��xn�V��Á�̄k�[��e�1/T��� ��G��4�=��0φ�P�n.��L���	��E�/�hn�����D�Km"O���*P�?t�Q5����ZBN�z���}��d��W\�ٗ||GB�gIwS���v�c)����i�4oL�,�t� ����4̊����G��%���6c8z�չ�EEa���W8����Ϗ��{.S��V4=&0�m]���uRC��]=���IRǮ��g�D���l����#6������0�id�a!�>�FS�Z㽚��x�}
����
��==�X~J��S`F���C5l�9Jt�Ϸ�0Ah���Q�!4{���������pR:D%1�M���<��G���^r

u�8Sc����Orde'�$��[?�Gca�wm��zH��[ۙv�u��?!��<�}�*��$w����"��vV���њʍi��.}�NF蝿<���$��H�Z#A��u�ya~�**kX�
N�|��[�QHjF0�r�q�Gٰ��+�5;��)��s�eH��Jv�B��pe6v�/8�%]�o\��/r��	&E�IB����>;σ��TW,o��q���f�"zH`zN�3�:���(dsݻ��u�>~�ž���)wK�����+��z�H���E�'M�4��c�
a@ڀWq{�,�Qxtq%բ��Y
w6
�4�]f�w��5L��΍��0C�p�$)���\;��P�����9/�3�0	3���N����ЋrG>CytcT��b�LjC&
���Cgcm�����Y����"����Ѫ�Ę��1���ˈ<O�����0U��9�jI/�S�)�j�1OSӘU�jƦ�.�R�Ua@<��^������O��V�Q��e���I�9
��B�3��)&z�d��V��V	���xIp�/9n��+C[����3� �'dV�þuOi�m]�-����ț��O�m��� !�I}#yg�4��}��H���/��Z'�H�Ž�=��:N 5��5E��n%z�>}F^?E�|��FE�N��,����TE����m_S����Ҫ�Q2Ɓ��1� ������h~�����Q)�Me$�֔�*x�QфsB�����1pگtKS�Э�;��M)#������7UvT�!�T�.����,{蚭��`�_�|�j�<��ր���&�n����5���癢�n��gBj��x�,��%}�<w��Q!oưLW:�!�������lW�V��G�{�S������t�D��rx�7�/%�^(ȅ�h�G��xo�Q�9
�|�� ��i�1i���ݠ��f��vT�p������{
�}�?�Yu]`g�n���)�\����jOO�Ǩi��Ph��׃�<�+�l�����V?�|��K�������X��	A�F8�y�;��z�
h�݊����z�����|!��")E����~���<k�$���q���,�Hs>[�W���2�8On�B�$�@�T����C�;@
�%j�5H�Vŀe����Ϥ��'s��m�(V��~�^�Q�J���qپ�o���▍�|k��E�"e�!©��P8�<�9.:B'|ؿ��X���{ԟ)���[�d1�@&���.���a�pC�C-�\�z�s����Sb��.��m)˔53��1C���-� 8�V������&�2[���>�+�,�^)G�Fq�N�?} }C�y���Y~1���!�f�z�\�`Ի��z��2�� ���P85�yn�%r��"�����$���B�,�+M������6�1��pl��,D��S��$'��xx�O�W�V�V�,H�B�t��<�n�q�p��.^Op�h��o�L{��lKlD��s�&Ci]�9��4�4����p����:�Lk
�!��c ���$�wc�F+�������V����Z3������e[���I|&�2��?��X���Q6X
N3�Jm��n�kh3E�C������֐�:���9o�:/w��w?�Z��E������&,.6{�Uk��4�:�	��n
w����Fa8����p�j|�AP]�t�]�]�ݘp���ݚ�&��tV��Y�=���vS���_�ϚY�
�ȸ�$���5��y�,np|L�:�yY��	�$@��f����e������W�Cg+�^^�ǀ��ĪEw=�IƐ퀩"y��u�בv��&���q]
,��!�.��J��{G�t"�u���T���i)V���"U}��<��2G�E¸�[��S���rSuL�Z���>�W����� ���s���c���7͉�ݴ�w.�C��ү�X1$�lt�E��f�U�XB��T��P7b�)��e���S���+kQ[���]�[T��0 ���H
,�?)�)>�dC��0�ΰ���9�D�+}��e����:�|���xr`.]�3�Pd�J�B�!���=7�h�4J��Qj#x����c��c�N�4�um��V��*�t$����jYl�}�AQD�]��B�֩f�3.�>�����������S�O���}�K`۹B��_Q-�(s�U����Խ"`5���AV�ܫ��7v��-�Ax� �H�(�C��G2l�Nk532d������LV�7qd��N�a�Kc]�v��Mt���bX�p�?\e;%�I]��%�G3���L�|JUI��(�x~���z�--?ӔC&#DNF�G�u�r������a����g�����;/���t���k��-^��������	�õ�o�{V�z��T��+n���B��)b/a�'���!�% M�pӵ?C�ƕ�/XYIU�M�yj��~ȯI2�w����Ue�6�b��%����X����(�zڌ 3|}!�q����9��I�Z�<@0��q�nT�R�5�l�AE[�����ep�4j%h�����mڑn1�2�����,�0��N��
{��F�頷/-[J���n��xIu��bk�}�rJv�a��$lە6���dE��V��&��_�V0��G�O)lHY̾&�M:�E_��q ����jc^�V�S����>�\U©w&����z�IM2�JUo���i�����YA{���O�7�����{+\���~��3b�!�Z^��1��-����艚N��a�ǭ�-I�Z���^�����PM��6	��9��󛮮��``�}�Oӆt${`���N�_�ה���y��Vk���1*�1d�ˋ'� ��J}�P3))<����#��g����J�WL�WW�W�/LX��6��5��*XΗh(�~�3�R"{ i�blWV(A+��m�@{��A�s}�F��������A�ԗ�\��t�C�3܋�u��E!]~��E�����O�iZ��+)�蕺M+:q7P�aORM��&"/��W�O�������ͬ�%-�5�3�g���dbMr�Ar2O�i�_^�N?��xQ��̰(�ͻΏ�83-�ۡX��3�dt��k�TA��s&m��\��?�<���n%f��c��u��Ѧx��#��$j}K�B}�"N�;,u�5Ԇ�p�`1x�.^K��Ml�j�B_���l��^.��j�>167D�SUS�V��,ZJ۶lxW�����ܛ� �/��T)Ey��L�(0�t�P`9�g�e}����nj޵|T2<*��n�\��l���L�g�H��}mf4�3P��p�L,���₰�y�k^U;�K�/����A}���CH��5꭯A�SY�v��1�\�!ޮRb�ӬJ�����)��:��� �Μ�y�l">�8�Y����ws����ೋG���e�,�ZT)����
Il#t���ᦹoo��Ѹie��q=�w+��\�r���}D��s׷S��b����A
����e���[��M��9���b\ܵ�z�t�:~��K)��6��9R2kh��Q��3@y�%3��cl/�rSc�m�F]7C	}'�*�Ľ͆J���'���D̚��|�V��c�O� �J�RZ�ؼ���;!���j��#pǕi.�#*�Z'ҒYݦ�S�C�l�>&x�Ӿւ@�)i��3K%͚��4���,@:��q�G9;�Ot��T��F�W��yɄ����3�����O��uK�H7��>gďK�-D"��Y���w�*خp�S�X�V�\��l�I��x�Ҽ��3A�M�O�U��f�qv��_�=uT��vO���M��{g{D+'Pe��P� [z�?�pn��P�������2�߇1Ъi	��Sh�У�bk8���)�9�Qvh[���{����/����F8`qͭ�����F�}|I�CT0�&ђm<�O9�D�ԕ�8��I�����
�����N�����"`W�~���ᶧxn"�R��Ӛ/!��>	"�~�����b�����i_�:G���'�S+[j3�ٯ�CN�%��Uq}�(������^���b��+d1��w�04��~?ބ�u���˖����C�ƾ��=���c���w�9�"��f7���E�ǟ$�	�r��~|92a���!j0��k/+%���$|9�xc`Ia4A!���/jbM�lFr��'�q��c<�`0�Kij�|V��yy��j^�gc,�ZP���Q/PAkh���X�. Ɋ��.Mϕ���WB�[�d�,�iR�	�J$�J�_��Z���fV�|N+�Z�w�	.��9�Wz�kr��&���um+�[����VLu��Cj���5Ĉw(�݌�&Me������փ��_����et~b��,/�@��)��Ԓ9)e���s�)KV0�a���$�^���R_Ѫ*��Sv�Qej��fZ�E�X�U��yh�ʖbj�����;8��L���^/��s��%0!̈DU�_c=�]u
��>�����C�FR�����uʘ=�&�,9m��P�GBgAf{��6IvUo?��о�^U������ƶY�&������f�Zo�[��P�,�O�3�	��[�Z~F-dY?�lB�@���C����䈜��#ǖ�[uW
妶���:���J��Q���sR0V�.����u��1u���JG�|P�� �
�����*�-�C��+�&kW�·������ɹ�Yx��)������vM��<7k�Y���t{0�^j���sB>p/ ���b�����K��[*�zpW��b�Y"b5;��Sގ�J!�h@x.�[�ڢg��"�i|N�n��|k5���X$������=�]�$薿��	�?V��Ϋ��%�>!?�.>�д�*���d����Q��:J�{��ۋ8��HB�A��<@V�g�u� �5�P#������}'l�b (�SfAް�'��HB
p�iJe����<*�ʹ	��:��001��"M4��$�/��?���ϣ�J5:��a�C+��Y�1��?�|�?Uٮ>�Ъ�o�\`�zˡݥL9��

�@��}R�	�{�/�f_U�M]�YU^o�%\�%5,�|�Ⱥ��ɋ~JY����zJUg�Q���4RJY�Y'���J�Ld�+�_Ζ�Y��� ]��n��h�A��z�w�W�s���^�F/Ćx�/�6ET��R���w���8�Xhdy�qg��ڞ���a�s��ژ�:���qq}%5F)�fn������?<��`e���4;-���	$���_�,�/����ZC�S�`ك3��XKqW_���x�MED����C�c���r��'�<�&+�ln�7�Mk���[�k�Ku��!��9��~-�4��ud�G���)��C ����eE�B:�o�����S�T��EC/�:[ɚ����=��dc�1(��0��xu���/��!�1C�2����㪪.|-yF%F B��ȅϡ#�wC��Uu��0l�U��w ���k�e=���%K�jb��G@*ȗ9�%�2���E>&�8������n?OH�XJA\oU��^�������p_�C��%K�a��֓:7_$N�B�y�?��g�EoC�U@�a���m1>@��xB �M<m�f�|�vBh���O�����Dǂ�y�oWM�����*���{����ml2ǖ���V��u�����d���O���F�w����5�\��_)^�]9{��=���~��U�1Vy;X$��j�م���C�����ڊ�t�65�xy��X�؊�ô�4��G]Ǵe}�'1�F�|�9���CO/s�E��!]���q�?�\R��=,2��fP�#����[Z�>	��'�% 6��ѐ�f�b%�sr�8'����x�g���a:�F�w+�`H�G��64�LCPL��#��.�P~n�+GQK��\�>�����0��-O5��8��*�b2o�e�&� '��t/�Ďg4���+f��n�ʲ�����3��˭Se�(�~:;�ְ�P�ҫ�#�;��+���&�hN��/Dx	�Y������g�I���	���R�g?n�S��?fzKVJ&F���`���^m�f �%K_��
�U����V�5���)������%�8ʼ2'��y�;��l:���D���W�P�ec@I
j蛋��wr�D ���\d�F_��3�|n<"^\���Y0�%	x��X2Gzi�<;e����&�l@_�Ne�G'
�Iv�ds��ުY���"�Xأġ�����ٺ�G3�L�	�PG�=/�t���-@�0b�$�!}�d3!~����ύ&�e#��V
IEٶLT?����~�2��+ʍC�	�]��Q�@n;�N�J��T=���%g�^�*���`�t�~�ى�;	`-��!�l�4���<M�s�G�O4F��A�r&��P5<��l&q ��>Vϳ�*�y�T�8��w:��Ě�_�I`��n�Р�	�lc�V)�.}���Lz�i��P9�nX'z���}���r=��|���3���wR��OX����	$�Gz�h��HI���@R��^)�.I?�y�2	��u6����ILk/y�Y�<R��]����Jq��4��~�r?\�Z�_Xd�ym����i�YІȼ��W�p"B���\p����X���apf�:6�I�#@����o�F�D�b��|���v��Mv%ׇj2�y��Ǣ'd#��I��m{��uHq0���)����cNw�<�(2:	��h���IXډ���-��9��~ʂ:�x8D-�&@�$�}��6Ϲo�@!��q��*�s���&J	?�F���%8m��٨C)Qa> 1�9J��y�d�k2@f��6����ePa&8I�i��
�>~��k�MG:q}��uĬ�F���X~�6��Y��#/�9+XMm�����PՏ��5ˇ)��ɾ_H�s�Ac,���t�����Mq�r�~�w1�o�L7����:,v6b���\m-�]khr}zM��6�5�<�yZr�&j��w�� �m���� *�d��c}��g�1Hⷤ�U��ѩO����l���W�"����''}������
��]5���5���!Dh�:V������#�`�T�وVU�$a�{�^�>0���t��ƀ�
�<�I l��5��F�A����R�f�!dŹ6�B*s�������1n7��sp#�7���>Ǯ�>Pu�NS,p������7����b
P�<bA�x�Dy;���>[�Q��v���:Rc�c�i�{sVnc��c����e��Ul2�|���TɈF��	�+�q!P�6T�i�f���U�����;��(^G�v.-M�Yn�5���p��)���2,��� ���f�,�:�~������:j9W�@�ZS���"�?�܆��8<a���*�
���"�Y�1o�&�a���ޟ8�X`h�f�I*:��ub7:$�η��U�b��F��e2��¸ =f��e�t&���ё;Q*�/�nL�B%�ֵ9ڼXLCEK��*�F�d�P�VU6t�U	��)��Fs�A>
��7��(n����	4Iq	׮�UZ����-��0qv�7BaP�}ɟ�,�41�뷁��%u�����,���M���)M30�Ty[���i�t�}��w�wk�kK�Yg%����o�"o_����h�!lQȥ�{�L�I`߸;*��ZG�#�oO�[h%�aG��!o��X����~��P�oJPo$��ȼ�Bk��^[::�����u:�[ �Dؗ�F�Z��A�n��Tm쭚����p�l��a/�`��볗��M����\����"��t�X(����$ϢN'|E��P����9M���P[�D�&��v	�+����c��6L;��[�¤���4�{�%Z֏�ʪ
Zb�x�¯�3�Ѓ5[c0�r�_�j
c��n�wp��*��9l��2��%]���J�|S�ぃ���^j�$�x�Yvv��LR������u�lT'��#�PK��bH��ឆ�;�=8��X�{4���������=��QMhv q�l�_�1���mD ��z_�&�~�{��.��6���1����v��H������Ğ�[�q�P*���i,ֵHp��D�V'��@N�g3��]еuF	����p�C���Ci�ݙ��j1��ͷ���F�L����8 ��zL]!�<�@��5��Ь�沀:��ؚ�U�L��q58��V��i����E����`r��OݐBJ7�S������ȋFppGH�oB�U�d���;�[��-���7����l!�ȽQ�ou�%����� sg�.`QRS��N�$�E�glZ�y��ư�\��R	��2ȥ�{(s��5B&����¤�ZB�?�V�)EWV�`���ّ��Zh�}���d���8���K�������u�R�o8��O�I��#���Vs��ަ�}լ_@��q(E`}�4���a\���K�@C%L5�5�[Ɏ5��!�V�&��1@��}��ݡ��� ����\���8�PuCc�ٸ�<8-�������~XsfjJ��N�����tn1/@2���Z���!��?��W<�h��Z�SV�c���uY��̉hT�������Qix#ۚR_�i�L���g?�����b�A�@e��'�	�IQдR�����W��`�6>��X�
L=΋�C���[�F�;%~��DvA�z� ^�@<3�I�s����
��E�+�8��PM~���na�����������	sn/��Zz�j$��2�)O���7*Q*{Dh�����:0����!/�Ex��E�m1,�i�5��{�8 ����d[�+Dhkc�Ml(�I>��Yi��ULY��V�ٰ��ox�Vr>��0�{ξ��|S�XyW@'~j��d��ۘ}�Z颉�#�2q,+����T�*ޯ�M�8�X;ű�J�ťX#�ɃR��l��+�4!:P�kw��S�]8_��n|��m�#��I�����3c�~�����;|*0]RD��&$)bu%**`��̏Y������\�,y��r���?�	G�z�/�z\!�7sE�B��� 5n��9�? q2�k�<)�t� 6l�/.�G+�)��%��L�(�����9���3>O4R$�s<���l\����,�\٭U��%��0���1���j������K��絑������l�����N�O|��?���wy��ߤdgd)���D]I�ɿ��6;5��[��qo ��$\[#JF�l�I�m�_�H����R�c�U$����񄔕s:�sE�L�[s6���O2��%My�d�.o�;񌥣$u4k�j�V^�R,!�ì5�BU%�q2��
Y�ʠY�Yi���s\�/B��WK��(�j�U��[��I�-駨�4I��"�p9H
PL���.�J��f��A��v�T'{�r���1�k��rW���0�}9���(�ćBJ���X����t�cW{�Zu�/k�5��!��/єѕ<���16��2>!۫����wa�T9��?RfP�pP(d�	ۢP}�D
2�6@1��ߗ��֑�r��k�J�XrNi5|���a�n�J{;�:|Q�?xt�w[?nօ��k���lF��~l'ӫ�S�	���
9X�~����=PR�H����@qP{� �_W�7�֭��PM''�9�'iSJE	i����m�$l&��1P�ǭ�q\�z@)��Z�6���bd�FE9�]�c�%=�9M��	B&3"��z�3���k��Hq��zA\���>��a��Z��c�%$��)��]���O��l��zF�TYԄ`�ĺ]�a�?Q�:t�t!@�C��Oq�������xd�pD�6������q��D�-N�a%�0q������d����Ѻ;">ݷ��b8ae�m�!��(�t����;B;�M��
���fZKj�ImS��vC��\F����
����D"f끾�t���� �S�ٹδx�l}��A�q��>p.���n����ׁG$��t`��M��?��!�Š	����W�n+��"f�x_�WH������ll8�q��Q��������90���[�����\#+���ז�Ɋ��P
\}��d������P���RYe���<~U��4ӀԽ�O�L�r��&)Á\���;�Jq����*�r��&�����������Pzw�<2��I��7���Yۋ���CS���)��Z�6)��\���|T�_��>�t֗�*�u-�Ό���x&C�A�A��"Yq��	%�+��`�|`�1`�Č�9�n�sy*�H�e��}à�ҵ��2Bm��]rސ M�]A��½���`���$٘�|)��Y ��~�p�M����$�"�G(��A�Rz��@�Y�MP	Ϳ�5��p�^P��R!���ܿ� ��� h� !@���p�4�=o����$�rI��Åy�.�F��$���I��i�mΪ�;�����Y����=�P*�2����QJ���(B�)0��K|���9n)������RK�hEw.l`�EC%t���d��]%r�7���G�(�<�U��"�7�� � 3¡�l�͛W�I���͉�g+B�$��XN�~m���R��ߌډ�`����1���u�f.m^�" ����#`�y^� e��HN�*�H��`{/���L�E���I̈́H�x��u_-=;p2xf�����Y��P�,�H�;y�h,�6���}��,*m Jd#�j�x�R63�Շ�����^JD7m^)������<d.���:3��ozb�U��1z��Ԏ��_d�����o'�5�{m��>K�wM��OQ�^�A�b�Kɭ~����4�Yѻ`������!�nj7�$�B���&�u���#�=;{E-��K|ra���EdO_6'�$ ����Շ���?Y$�e��9"G �łD���}#���z:$	_����)ҽC	,�vQ���X������+γ�)	�n@>$j��^���-J|�aL�k{�W�j9�h� �NhN8>Fr�J���L�XcTߗ��7�b�J����N�_��cB��e�f�>�X5��֍#?��7��[M�F�*����rJ�'pR��ͤi*dI�O/���:���Tku<���O��˨�:�lC�^�&4.!�k�;�]��O;<M�D�����R�I�l�o��Ᏽ4r�fP��4��o?�U�#��\��}��]ρu�\n�F&oL��u�/j�}�&`ߞ�|�KC�n���72ݵ�|����`���UF�
[T�4m��+>B�g���s��l|���eO?c.�@�]��>�_�8�<hO�5���Ju*L3	N&���������9R�,s7���X�:��t���*�����zٓ�qx�7d�yu���~~�N�)^������Q	�����962���L�X?�'�$��3����<o� �sV̑�ڥ��3���ʖ�}��c=]�ڔI�B �~����&�-�U �k��P���d���	3�c�����XP-8N*Q���<m\d�&�	2��3�}�6e"���Hr���880i(��(Y�Ī]h0�]�����>�79�X��	h��(����L
�_���ۧ,2������y��������w���uΚ����?�NdvA�)r���bc�����h��A�h��K�>MX���U)qd{�y����jХ�-�+_�|���U�`�pl�@5Hk�!k�z\m���q��n�J�a���S�+��*�i�7��EN%>�W4�����w�'�z~�0VC ��ѣg�sE�,��4�ӎqa���R�[�b?Tz}\d��@Z��[TB|�27=X?٢��a��t=7��^�R����U�R���y��a["�I9K���M1�{;婻��h|�S������א4S����6ْ�m#��QG����~Kg��:�>�;��|��:6<{c��Z����q�Rq�3��/�_��Λ0m�>ݗ����� �=uf=�g���θ,=�5�d�?ڸ#\��/a����]*���]�@ߕha�E^����(�bo�%�jN>0o���^�\4fDW�L �ɐb��+A}}�O��x�e����2��{c��ȡ�\�.��N���n�?o�sy �'WpŰb�@eF�ʻ����i�=;��B��՚�:%�D�O���q�'��a$-5\=fX�H��XB��s,l�;�ĵ>���0O���8r�y%8�8�{j�����o5uJĔe"�Q��OX�D+�?1�D����d�m�L's��84M��*����:��w�$���ᦛ�د�.G�{�8V�[�!C����)z�Ad&ӗ�/�L�V���IF�X�=Zz&d��X������$�r.]��DC�F6�=�*�YƳ��W�l��u��-}����V�uk�䑣r�O��W�6���{�)�Ѩ6�"�� �q�a��V?��/X�4Z˘�F4�4RQge���ޗ02^µtdR6�`:���	n�^m��,��L,3���N��y�&�z dS�p�vA���z)Q4��/��;�j4����#GGd)�8V��Z�{�ܽW�ZX�����P�m��{0ؖ(�eϝ�E_(�i�MO#�I�������f���T��@O���3 �&ŏ�7tx+��ǐ^5����C��kª�3�PF]�r E�\D�0N��l�+4d�:$a>�RT�:�;FX�=nG��IDi�����P��c�=]{���~Zg� �3U1$M�\�'�nYg����xa���ϢR.a��F���qO�j���g�~��V�K�[�Do�w2�ԑ�9�,�c}�ڃ�O��TT��	�mM�0�n�r"G����UCƾ=�YCܢ�F髽�~C��78�y2���t]�C�#êX�3Mf\�a�!�E�a�,_F۸L����A�v>L�<c�'V��Ӟ��>R�伉���Y#��Y9	)[*�-��g]T�o�H_��f 6hgLXBKT��xp�Z�x��fa���ݗI�����>�5 �jݾ 2N�ӎ�Gl�Awֶؚ_޼6�n1���+�0O�!�1����������L��v?k�k����@��Фॷ�>�*\�l������/��Q�.̅K��������P��+�7��O�|_������V��hl坯����b��}���cnT���c3h�~�n�[%u�9V�Tpt��u�e�@V�kz툄�LR�����$����0U�F��l�G%�:՝��`m�0%$�'r*�ʒ�A}�}�_8���b�T�v�d~�`����	m�w�s�ݽs]�Kx��a~�^F� ��}/z��ٺ.X�ǉM+���+U$�	$�顺>i+K�#��y�qD��h�?��ڭ�KJ���h%>�':�z��l���"��)L�#ט�4xy��;�?0$�q��7lf$�jL"S�s����x�WF���o�3d����
�:,l.��Oq�Id�Bn��},�Y?(�����}Y��y-´1�L����)L�h<�n�nt*|t�c�䠯ĸ�8�`�!����3TAf����Ynb�f�MR�1�kj<?�C�:WF)7���!;ֲ=ź˗��]���_੅�|�}o&���ؠ5_�3,�åӃ�/��#��� A)�%{a}8�{��]�[�wl�cܬ���w����L���l3]|Q�;����LE�[�ɸ��Blx����LO����⣾!��[ ���>��$��L�~���_�}	y��\*ސϟzt�@$�b���N��g]`��n�cƻ:����D���67�=���y.&�4�<�ʇ���PTO������[���?�ㅷ�8eYNw�������3�y<d�M�B�Z���i�.T����C`ǓkP?Y1���\�;�ե�`�Lu�ه��l�)�[�gO�*K�FkA�k�T����Q ,�2b �o�� ���J��J�l�����V�)�B2����P�%�^�j��,;ao6�k^M��]V������)P1~�|!
��&(�m
�6����~�ĸi�}n*�8;��:l<s&o,�:�r��h��q}��޼����˘$��%G?��ì���p ���Pڞ2�k$�N��jCf����q!!w}~��\����Z�X�z��g���j�n\�����
dM���_m�߻�'_��^djOp��hcb��W�Щ��7湯K#�db�ů "[G���o3�"����3}�93��m�� L��"�6w�<=�F���Bl�f �,���N�����b�{!���u�j9 t���F�]!�V�OI�� Y���O+h;���w�-�W�)k���E����u6��m
�w�dzg�?�30q}1Ʈ-p5�/l���;.襧���I�����8N�"Vc?Cٶj[��+d�� n:CM�յ)z8�Z���:L�-@��R�☬����M����PW� ���'����R� ϱ�L�.��2KF��p�6�+�Ӳ9��-�_1�@e�۹������<tz�5��m�0=���`����-.5㺩e���,�Vw鮱��.������i�I����	����i�N����̃÷=��?�ׇH�ݯe� U5_4��݊�5�jPR�m�^����`raG�YyTAbql�;������U������� ���7J����#���/�g`��H�Y���㘯'��8G�!{��P9*�7���ų��ق��'��jM`�e5�|�74����18dr���'+�8j#��,�t�6*'���Bh��s5�1�Z�����BA�ز�!�\&ٻj2hPE��,���0�*TQ�,�7ǡ,��,�*����g����7$���:,t�f��VB�Ĉ:.�G����_�ӝ\jp-�H3_��\�e�]tql����&E7�K�>�6�cs{��疃ݖ��^�*��X��ka<�)�o��H��+���@>{9g���P��h����J��c��B�N���]�ҹ$�%P��m<aE�S��)�����Aa5���h!���1W���]D��v��\�!�vET��1���� u&� `��w���c端�jMn .n����2�,0�?6f��Mj��W�	�n`ڀ�����z��W{jhx�I*sm����xّ҈,��ݠ��[�d8�Ck���|ݼ��Za�'V���x�f��[�t�3�hxA%�M�18>o�0��[ ڋ7/��ѷ�D[ X����u�?y�س�#o�&8����	o1��mp.e�?N��~e�*
�����b7�)����ۿ/���^F���ϬQ�$�k\?3����~�dTpK}ZHDXT���*��}���vlw��<�#g''zu�Y��i'w��]�s��.�'/]��IM�|�#3�� =<
�|M*r�O\C#��z�ߴ��9 ����������o���IX6H@��<Dna���Ǘf���z]�1l��.��H�c:�?���DO-^d�3�"��$K�'JH��~��Cw|Y��tKUZ�G\n�Ԩg����U�T�G\j�<cFl�s��9����l��<)f)�$��ȸ.[xJ�(���,�#�RL�U�S� B
�j6� ��� �y�G�zL�|�� ژ�p�n��\�Ci�:j5Z�3� ``!��xX�?mx
J�"^y���~iT��M��v���k�'V�@N�(��6�UX!-���c���O5^�(A|�"�4ߕ#7�%�������
��Qs���9A�B�V62<�%Bw	� ��*W��� �J��۝�?���1�o��oft�����LCv̻ ZiKi������CP�p��=��p�+(WS�hܕ�B)g	����w]X�.=!�@?p�����N�s��z;޹3�-��������E�z���:�D���,�r:���4X���bT���m��Ʉ�ߧy�=����Ob�)�|ixIn�ζ1X�]�'ߩm��eէ�g��D���ۗ"JE�1��&[��0�N�#6(.��hY�Iqwf���k�ʣ�,�t���i�I�-��Z�~
�Y֒?�||*j�{�i�'�G�LEX�����<�xcSF�&�M���7W��X����\B�VZ���uO\b@/e3>ߕ�=:e$�?E�%o�p۸�R_�ѸFsG��ɉ�|3�!BWBp�p��������U�aV��'�ƴj0��?�j�}��0��D%�Tt�<=xέYR��|ƽ�=%��hݪ1��@!�x��}�驟���T�8$�4qK�+�9?��k�g��uGI�.���<u�o�eξ*�C!�Y��'T�5#��xv|\ވ�,�bx{��Y>�a�B��^�?L��*5�hҬ4����3j�|"�tx���ٳ�ۇ@ɂ���E`aZm�E+��?��H͂�x(�zj6�N����Ն+�y2�v���d�o�ܸ���j,/�k�0��$cJmZ��g��N"������*�u�̈i�I�����jT%�p�]��VR���I������@mI��t�V�̈'Z�(G!�9�T$�����_���M��A>9p<h7�Bh�d;�ꦐ�n)q�p9Xo U����Z��8�/y����Eٿ������qM<f�#��o����# �`\}93c������(��l�
o�����CÁ�r�6tN����5��m0�(b���m����=L���� �x�TV���Nm����C��3�nv�Z���ޢL
~��z'�����;�gh땕��k{ı>bG��}�Bc��~����i/���ݹ>��MQZ�����g`�9Մ**;�bѺ�nd2�O����;�7�X�Z�� ��'Jiջe\�f]?�����i�4�[�ٮ��B�x4��x0���Ԭȓ��zx��1�b��MV*OGT. PQ.��U�q9��>+S∈����4���β��1)��������7���I�������͟##'�+d��ٍ�'% 0�G$���M�%��"�[��T�(%����a|<�!%��-�e�,
����g/L��o�H�H}��Ca^_�[[g�{0:���iC��c&�3C��%���毡el�Y ���\@z.!���*ɫo�6P�msA<ZV}?~�K\���A��:Keop&�?��Ĳˤ�Uߩ��z�2�uU�U*�pԯ�! �}�g$���!�6��oc���BX��[vi�=�����52�d�2��*�I�=9"u�ih���&��E��vb�@(��(^���xK`8{D��N��b�M�)a��X� �[$��P��؍`"���m(�SE���!-�SY-
�W�|��2u�~�ԋ$+���x�['�y�|>̯.�?Q���;B��P:��̅����<b��cş�G+E��~�곓�j�ā+s��*"gZ3S�Z�`�����&U?A-��o�Z�Yj�MR1��v�O�K[J���z�G��s���::$c���9kO!��@�޵� ܆�#Pa��%5��j����J�1�K�+�o'l5e!���#( �/�|^J�f�iNa��L�����ʍ�F���� =�^�d
�f�[QXMӇ����A[��^ɝ#�s���H��!@��s)��Ι��2zx%W��׶1ܦ��;� �/�{'�Vx��OY6��U���	ni�r:r�GJħԅ�I��vO* LZ�BN��+���.*+����CF$N��:��`F��g(���g�N�@���P7t�`$��l-h"KB��+i}�+T�[âC�`���ƫ������F�9�<�X�~u��Tz��\�p���$5�բp/�D�QH�l�i=�) 8�����ZU���9 ���Q��w�^g�U�-r��7 k���CjQa��`x�TS���`	'<d�^Հ�y'FԮ�bh\o~ϐRC����y�%��D⣁�-"�O���v9^Kj"0�:=_�](+����O]�m
�� A������Iu�Y1����X�umu�W��(������$@E�����4�_�t�-/.�2BB&(�vO�?gۭ�
<����Y���7j{@��#.1hh��M��K�Y�sYԺN�f�DP,ym\��|>�DH�|�{\-h('#G�i��T���}g�n±���H�q�6�[C9EC�@��:\�������j��A|�ly��Z��s�&r �J�~60��T�dP�Pli E��-��):��	��?[����1�C[�
�cE�j��զ�l��D��q@�DH�����EW�����)t(%�)ń�q���a��9�A��	"$� �e��2ćoo+�WЩ���y/n2;���4)k�
s��Ek'����B�/ud)e�^�OouW��Mu��:����uS���t�ų��E
�d�҅�����.���+h��cB�&x��%��Y72|�c���;���Dq����2%�+L��F���/�J�������R������YDe1bp���6�4у^�Cp�f�<;�ʚ���y^�^H�g=JA�Զ�-f�hq�Y>�L?������_�)������Ӎ9�����&˨�9�R����֜<����z��BMVʰm���x�nkZxC0�ාndo���ٹ>���6�3���pp��m� w���J���t�6�u `���e�m�0�5�Bq{��q=o��۝A�+��J ��F�	!��9z:�7B�%=�QWR`�-�՜+C��]��ˑS��F�Fd��2Y[r����v�\�j]#3�I�rFn[���0c���Nq�,�𨀕b�D�I 5����ߧg,��)Zр�J��QKY�L�$9�YR�B{��qd[��==��l껨�;'6(Wֳ��N�FYF�lw4[( hV�(q8���Cݝ�HU�ݣ��]ݕ��]���,��.y����^?�W����z!>�M���Ҽ�7ˢj��F+7>q܍ɼ��[8/��W��*b��UopwJu�	;0V�>���E����N'�w��Y�_���P5Z�:�2�&YY���6�9�s��7��p=ս��?�巩|gu�
���A
"�$�V���ȴ�I����8�A�Q��:�Î	�P�-Ϗa�1�����`����fx�i�N�G\%MƄ���zUt�S��ަPjQv�'*��
.y�F��Ty1�b��
~=����OS�N������M�=5S� �����A�"�xhFQ�C���'��=�H�
K��J�Q�j��B��c����_L�(_ֲ�|'�ȴ���l����.���tk�#�3�H��X����@��"=_��?�C|r�{;\�
�|a̘��Y�x;��OL[�@�o}w������-�������^��D�a{VKxP�������-29�n�h�]: �z	��*n! ��,X�o����� �n��C�ޖ{�C`�������	�l|�}����p�w
V���6�zn�d^4b���H�&�s"M�P�Nh[p�;���f�R �&��O��oe�j��p^�xkn��C�Th�k�%u�����巢��&3��bʹ�� ϒ%��"�\�3�X�n�l�ռ�cC���O,9lgLQ�ڔ�HG����T��I,�<���N�F��g<�i�?mf��K�+��Y��T���^�Y�1S�����y��A_PEڿ�&H��ך��bs
~ljE�o��C�RV܏)� ��.5�ʭ�Ŷ����֪�p��	�����\w��]��8�N^m9�co^?A��:=V�WFz�������������+��\�*�N_�M#ˏJ��$L˫x����En���C��8�&���Yխ���Ȱ�lf�fK�f}r�d�������8�±~[�W[���O�j��s+�ǘ���'�d�A�	�u�e91�v�J�� ��)�� ȡ�̧=��L���ؖ�%�fj>p��\\�j,��g�B��#:��g�[�;^c�zr�V�w<ߋB�ǆ��〬�In/�ޤ�'�@��w�<A�A�/��٥����,[@]��dSe·.�=�!�d���e= A���g6!.� ]Z����u��N��wק�-�؏�:{��axL���VB��V���0�߇O��P�38|I��-29��?ۍ�O�ip �]Ac�`��ZIj^�6]�����8��ʴ���ƟY�[�� ��0�0�fx&�5s6Q�X�/�ƒ?��G�j�<��eH;��C�<*Β���i�U�ŷ��H9g�:pm��л��J��dt�T��w$�F�)�����0h_��_�&\��1�c0�["m���#}Ѱ���Zs+�Bi���p5[�Mo�'�>�"��
0�� |�/��ֈ�q[Q'� �B��x�T�]����m��)�?��S3*Q�Q�ґ,�;�"�Pk2d�T��|"�֛i�ݲ�6a=�[	}�����˟�U��v�'���c�M����q>(`��7-X�b6ϭy�*�6���Hڎ~�&m�}�����ov(��g ������x-�`/�]��g��@��;K��=�_il�* 8�������
�����_:b<���;�B�8�a�3��}����߀�>��cS���~�jfCCX�Id� �k/�f��dː���`J�T��b�ۦ߫8ϫH�,��n����	7OB�r��s^� îF��2]�sH+���m��BIa�|

���	��x.�6M�D�Laj����p˅��R��Ҧ��A��y,iB����gC����P�#+����E!_����Pؠ~�}1�;~a:�qRՠ��ʈ|�q`G�M���L��*�[͉�-`����̷̔F�y^B�Y��b5FILc4�` �Pઌg�7�fW���G��c��0h�Q�4Ҋ���_v�c�&?���t6�[�����J��u�"b���>q|�Ӊ��#��Apl�tm��{�FBK�4^1�@;�űl���A>�ى8'�AŎ�O���9�J�I��6�EE� �INc:��H3�bʙ&2��`_��E��Ě*w��y�zLn���-����������V�Q���x��6�5>b����fkc3Z⑀E��*�EuF�Nc�-48��p&�RlV~IJ�.J����,T�9��Ϫ)q)��{��,c.�Ol8�U�$��$BW|H65�Y���}F	z^���%
`�g��p|+ˍ�|��A�\�<ĝ0��_%���-ze>&i���n��F*��$δ�5Ĭ���%6��8āׯI�o�hx�ĲV���?�G��k��yq��M�-��UCk��p@R,�;�=�z2�W��22.\֖f_M
_B�i�ǆd=_�e�R��eMT �Ҿ�s��t��8Ѿ��/n�|Œ$��(��,�����TQ��:m���p=�9ݙ��x ��D��8I�<����j���
}{M�~8������mNw�I�.d����}P�fzyUG�H�٘�1ѫ��[�m�70�}�j�"���n'�(?���5j�<w���r�:#ZL(�(]ԈS�U�t��������Z'{�{����=`���o��;OQ�UZ>�:����2�����&\t�]�䮎p��{W��.������ʑ���������ˤ��a�'[�o�]N��M����椄�*�_M��8�sg4�u��/��3�Ȍ����X��j<G�ۣG�'C"g J�%|�'0|ݠ��s��>d9D?�`k��������E4���@+�ïq���9�W�^`���׾�ͿMJ�V3�O0M��T y�~��]*�M��,�'���9����I��%���f͒Eaހ��u�..5rtO���`P����W��S�w�+d
,!�4;8 ���E�{p�!I����G'�6�<�V���%���-��uǦ��^�0 ڜ\�_���?�K��F}`��v N�po���:�@*�EA�����b�k3L��F��3�U�Ͷ��@���Mi(�������/�����)���k]�Er�Z^�GС�Yx�D���Gr�,�{"�Ɲ3�|5e�21���:�I�y��Kp��1;�QI;87~D|���i�ڳ��~t����gݖ��E<!u��+[�x3+?}L��>����$�ݟ"�<�13�{��������H��xkw/\/u��ݠFjQ��<w��$���h�M����C�k�FX��,4��p:��*���ȓS�Z"��X��˥�r�a8��w0Q#E�t~����Ӗ�IFt��o�F%��'L���i��kvu���,t��#������
��2ܤ��Ds��=-��3q!^1�럥q ڍ�h�B:�~��M�S;�j>�q�j�ߦ4li�r�z�K�ͫ�W�{=���r�a�k�W��2���`���Tp=����ثSe����r��I�6����?��}@��>ZX:�QW�,�p���p�/�
1x��ݘ����H�3�E�p�1 |S�&��Fϩ�<�~+^����E�~5gb�1ȝ�d|7��Z�lF�U�(�&��>>���p���6_��p/Jw���W{��R�L+ߎA�5��)��*��ҝ�R�ڜ'�j��%J�Bv���R�O)��Y�@/��[�n\��ʥ�e���=��;{�)%L�%'f�=�_	Zr
��"��'GT��Le��3K�hi'�a^�Ӈ�fL�E�)��8���M>��^����u���cl{�R�7˥+���� k3��ݰ¸��l?,VC��6��Aܦ�䚰J*z��p-�@9F��Bg`����V^�A��)�E�.&�$�c�׿���U�x���m;�1�J��9ɣ�SL�TN�-��'2��U'~�O�*����qL��o��_2�_�6����2��l��,�w��m�c�����KhF��˜K�Hs������8�9{;���0�@:���y!�m�]��+T�'�F���j��UՖx�Ͻ�=2F�d��
B��,$��"�9�1�a�߾�����?��d���jw����"�UQv�cR�u�lyVɵ�����Yd�I�����3]k��t>t`@Fˡ�La*����U$j�{-�糞$߳�8PN�p�^�䢛�Hi���D|�w��lp�t|��v��ƭ��&��m��o6�o�X��������k$M�j��ncE$�`���nB��7�ה��@�GP�QK�.��%���!F���J)rrf����6R
�0J�Oh��5gu���L�O�Fg��iz%*�{~�� X�i5���J���;�/ҏ"���>� D+��|v�,	ץ�b��3�[�C�:�"�"m"Կ�T����{>Lu�HZ�c��p/�?Q%j���	��E_��@�j�M �U�I���'M��l�2,����g�~w]�����}��V��,�ZܐN	D�9��(5'z�Dt%����v��{��~�4�8.<��q[$i+�h$�o)Ҥ���^}��y�w�ʪG|}��}�8�3�]c&�&��9o��N���	2��z�EAE��T�	C��>�US=N�(C�"%����t�h��3��#Q�	^4�D+��6ż�c�1�9�cA�.):��#�o��`���/�}���^3��@i �2j�__�voq��֢�+����+�\n
f\��e�WK�d��������op��e��z�I%��b�U]�n׏U�w�������s���a�+����N����b�j��V����	�w��w)^���.�k'�:��#Z�M�p�)�л'j$�T6��@kt[�d7-��Kg��qN�;��$Y�d����s)���*����8��f\��h��4�[���b�ʶ%$��e�-���f�
8���q@�V��%�В�_�F;RA�� tJ�ςu�\=�3�S`\)~���)����5�G�XPK�޳]�X�����.�\�E�%��҃���qU
�]������w/I�4Ig�u�d�8������F�2�{���a�=�d�?�6�}]�T�eZ҆th���ϩSѮ�� ,�l#��Y>K�ݏ����5�����G�<�֐���sK�~�
�	/�'{�2;nc�R��X�4�.(����"�?�\o�[#3���*�*\x��w��*�0r�/�Up�����ߚ���A�h�G ���[��z�v�@e��f�j�ex'`)0a*,�%�N��Q�B��A8��W0�\-7}us���H����6y4�f�$O?���{�X�8B��5�*ia2�'P%L�k�UߚM,t/#S'hvV��^X��=��+�'Kփ<�#� �2���n�j0-��䉬��}�#y�=�	�r u��`�)��!�i��(����hRx�ᨇ���Dr�|�\�%�G	ƕ�c�.�ګ~v�+v��Ѵ���@�����s�2z/�ru���f9�,��g()�xc�9���9)p��
�6=l���U����!z�9��{�.8#�* �*�����B���1`�2!`Lo!�o�'dh���vN8]Q�!�
&��n��H��C�M9��Ki�)�J]Џ3若鈪��G,ä=�����u膀��sGYy��,ӦЫS�8?jb�_┱�W�+C�?Λ%OÂ>��u��/�~`���- W�(��I������c#ڶ���9��I�X��ޅG�bJ���K9�_����B������>�Z]U��&�h�ӌ\�y��e��ʻ���;�� `k�þ�~��Ź�ar�3��x� P�XI����<��D,^)�8�`�m�7.��������>RB�[X)rH<sp&�d���~�� �Q�>)�"�� �ê�|���e��'1�f���~�]ҽ�E�*8ǻ��&)�n�C)N�և�����8�q�
���!=�i�yp�D�}�`C�;v�^�Y�mL� ��&�	��bf@(��TV�]S��Ҧ��E��l��b(.D4���:S����`L(���������]�F�)í�UM1� Z��[�]qQ�i��MX8iy��BM\&��_�M��A���i�@�נ<���OD~
s&O�p�sU�h����}�C+_��`@��z���%�<̫Z�6@�
@i��)�Xg�x.�!�+0�������Af预�u+�ӌ���$��������7��!�_�k���3P���*�Q@�Ly��M��.}yDK$�J<2�wu�$�`�%���hr�5ڛs���$�0p��6,�V�	^��K�h<���P ��C�/�S~��t+��$�V}q�M5�Ұ5O�۹(/���k����G%�&��A#�]���>�M�O�%�Q̄�F�6�q�j��),���Ey]Gn���ܤ큮a�	py�֎�êvJRO��*�>v۝7sܢ79z��UǶ >� �[��<�f��&wwM������tD-s�KB�������nE�Q03�f��v���3�/W X��pCW<{U[�D�2j�4�٘ff7��������
���=�E(�
�lXI�uH���{)ҕ����OR�B,�Y
I��e�謥J[8Uㆢ�Oǿi�Hz��5��E�[���;Q�=i
 !55������7��#����H�;�^lkI��d{����@�g�Y��F|B��1j�^r-��Z�)���}O&�*�Ζ�g�@U� �i��q��ϸE��v<�\1��B�TĆ����ꨩ�,���"��� �����Ǝ}�
\�����!���^/���:4v Z�IFB�k0��l�ji\�bQ�l%a�r����=�	�jd��R�V$E}+`�:{@���5�Tp�h,�4ۚ���$/����IV��'��Rˀ>y�L�!�Bl�ݖ�i'�
j�!3����}ʊY4h��*Bk��ϼ,9J����k�#�� ��5�NP�ϭ2X}d4�2�U����j�-�W��T���
�>�\��JI���$�#�8��aWF?v����l�M�������qFrҨ�2v@pE���]����%p`�m�q
 #O�d�^��U6VD�3<�f�9��עiB�i�0Y�J\�Љ��|x��#��H�ǟ�MŁ,�N.�س�E�����'� 6�>��'�ےp��������k�cG�xk�6^����xv����B�N?���crAz�"/q��y���cMZ9Sw��G>���쳂S
�?U����rY#2
#K��"�v�H}�Y�
x�����`;]�I�/Z�
��I���T@����v��lB�a���]�s[~ZȠ7"�l^;���?FU�[

NYB��p�[A&sE\ �r�S���׿��j�����O�Q�z�E���jr@4���(�غt�����$2��j�QzP%�w���}�'�0/�V�N���i���iQ=�g��9�`���M���V���9Ȉv��y� �Z�9�P��g�oFTA��:�E�@E[�+�ܝ��𤔪M��K��U��<)Ʃ��qqX3�y$L8�yK�5��:{���P�5w�O΍-w]8��+�b4�4��P��\D>��u���w6k��g���ɖ�H&���Uz��Ę-
�t<�������&���m=>��T��|+?�?�<Ǳ4N��o��L���_[�=Â�(*z�?>f���-�G�T�!�
��#�Ц�Ӡ"�Wy��/��v&�ju��v�*k}����o����h��y��_` �L��d��^��|~�x�~���n��fP5f�D�y��/d#��.k����3]&�&��f�$..�������]P�?�C?3������Ě����9�q��~Z�qH>�������n5\�9�v�*O�r�\�s��	�D�!]kF�	�=l�t������i`+���Ǎ�y��u ̱��G3q�$L�
��\��d:����lwW� &���|6J����ٹ��|}K��f�:��2-ޔ�*�%�h6����s �`�����;p���g`�Z,��N���lNlYpʄ�U�����<����+��	�8����o�9`�^Τ6��n�D��YI��T�j�
�mH��p9�
���4/�y0��(IoY�Ê��Ǝ�m���w�]q����m�֊r�$�R$c6(a��0�$cW9�f�8�6J"-�W�a�"ƞ?�)�\	���Yb$�F9�y��ƕ�+�r���^=�K�Gc������z"%�B�I(�:O�̬���
bXTS.�})c5��F����0d0Q�vW	�w�Ѐ������iFq��Ȳ��v`������2Ě��x�+4)S9F�u3&���l�@��/ƈ7��Ի�ߊy�rB>��2#c��������u���^�I�!���G�3�8�hң"�;��Ո�3P	��TC�W�$�2a�ZLb8�ܣ����z����H�+��וּ�1W���ۺ��%�v)3�KP�zi�d���RЋA\G� �m�܅󿙣z�aI�����u!sK�Z�t�:���4�<�(g�J�mgwڱj�jpb�K������4낕�%I����a�7y(�9l���le��E�M�>�f��=D�R��:;������øZ�^x|X,hޗ~�3�]�@�3:�'_R�.��
��͔�6<�%���P�������'f��N����:��U���������ߴ漛�5ǌ�!D4 >לE�67DDb�mlCL���X�7%q����HҲ��yW�{D�2V\�?��ϭ�?���4a@�Y�=���L�8#"�1�r�G?��J �*I��i��	�-�l�\"}��۹M;�N&�8  r�U4m��w�$�;�*��0:,�oVN���Pg������0aˢR����]�<8z�S�ܼ�a\`0S�k�MQ��c����4�3��K2��WU�#�A��<Z�o��{��5�ڳP�\c��U�A�v�i<A/�:�S;L�H��'3�5�}T	f��#��Γ&2���, ����խsÂ����L>��d��˼u����?���8��b��^��w':,���Qӫd/��*��[����NTb\_�0M��QU+G�N���6i��2.s�Ɔ�[-���\m��-���:������%y�2f��Go+Q��!��Ghꑭ��t @��1b���,��52���>�1�F<����[ݸe���5��G��0i��]��q�ܝ@f�V�%t������gtK���,l�+pG>]��	���(@�j�ocLamY���4�~.�v�O����]q��[y�F��o�y����F�q �t�zZ�{�Z���Uʹ"׎�962R��׼^��^sb��1R�����_gS���8����qM���T��-�Z�@��7;4��asw��jK��D�� �/UGx���1(Hz灒���{пP΂A�,���Y=�J��z�26�X38����$.��}|��m�U���Y��r�t��o��o;(�R��{�%�����ims5�#x���rg��S\q/�0�k֓Sīʹ��(�\��f?`��b3���$9��{�LF�F���$��y��f&^���ȣ0�Q�B{��LC(���:^O-�[p��ܶ �4q�7Ȗ�����x<|s-�tLa��d�]o���)����|�X��a�QɃ�͈1<3��d�łR�I0�gb:{�hƛ�v9����8���P�%�g�J�4���#������{Ǘ*L5�rǮˤ�@�H����04J�&�Է�����ѯ�1�������F�[	L'Z�3Y��TNh�����4��^��$"����+GQ�by�=�[�i�=2'ˌ�����k?f���	�]a%��_�Q%*��ȳ!⾹��:�$h͇���GdFK��[�ok����d�x���*����:5C�f��v���tn&���l�@��{ w8��5`fH�.��e��?�0l��Bw�2���0t'��?�\���N��q1���;�j��ZT|��!"�*S�i`j��7aP������Z�S%_z�c�_(j�⟀�(�7 =�����ό浘��&����gύ�?Y1\���u4݀��=�I�������h�Yw&��R@M��EE�:�����Hj�2AiSk����}��SY�vG�%X����z��,���f��W\�����lc��ټ�ԧ˳ �5��߰��v�F���#>�ar�F�DN��5���q�գ&��}b��ˀ���#���V=5sQBq����Ш�Ψ[�ׯ4&��^��i!Q�`�d�{5�Lm�h<�S��'1����a�����m[ZL��G�*3�1P����c����Z������\C����C������ZZ6%�*��).9�N����L��ӷ�#�R�1�Z�_�" �*��xJZ8I�<՞g,�I�JߜE���t���X�誑>�&��M�|��;_t��w�WN�FM��}҉+K]���e)���Ve�X꣙}W����FND��h���-� -M᧎�9JP�'���V�X�p>�9K�Ғ�3j�!��F�}�i�<5*=�T�a���v!Xj�d�Y���$)��@��y��妐��~�vy��!lI;~x�T�uL���'U�^���	�6��m�l[��'��Ǉ���\q���Q �4h�7&k�қ/�YF7�l_ u	�+}����!o�P�5`t�z�S������:��eΏ<]�1v,Jӏ�훼�WǱ#٥)�H�T_yh�F�Kh�I��лUm�Lw���0��7,��&����UI\�sD�x@�|ź����>םt򡁮7�O}ϐ��;ǡ) 9[�@gB��(V�Bd�g���T�ݤH�Tk�	��Z| M�
�dPN���������n��߆1_`�+_�eû!O0U�1��������k�q�3�@b�Vr��e�+�I��լ�S��ͥ	v4�|�3�dn�K|�?�p*�����*8�*��oVV�&ܼJh��խT�0�F���Ll`l��]��ߏX�C�R�0�h��=r���*�~w7��2�Ox)}-e��!.��8	 �1���yz�8�o�\"�5��U/��a����.G=�vP�S�`�O<��t,7�	���z�. ���g�Y{���a�!K3s����2�t`�vG(�	B�]��E�@�׬[Li �k	�lzw0m���Cʪ���;�4mg&�ip�L8�?�����ju�E"5�����M�=D5m��k���PH�X����>���	��sc%uvb�-�3�%ȬC}T���H��r��*WưQ.��X�W���ɫ�Y͚�+ݺ���f�sr=���Ud��v�@���`�k�XHpY�ёtC>9�G��vbh����C�o]��M��)hu��Ԑ�&�;��Gm��6j�e8h��T�П�7Y�����SJ�}G�jaKT�������a�x��+�k͢H���5b���h�rmh�bګ�zq� �e�jn 	`����|2y?oA>�%1$����=��Ѷ�����G �k��@�(���)I[�\fV��8]G���#(2�JT+e��KV�H4g��L��G����t�N���?(a{ ��m��|�1��ץ<v�'^ti{�}�lk=wF� �$j����W{���]����2���T�#b���P�r��ׂ�g�;x�`��8���県�X)S�u��yNsC`
7�7n���y��\'��ġ�7�F�٫E�&�igɬK���|��<���8d�q]U`V��pqY���7��nl�k�y�W��4|ŀ����!�Ə�4�B�kF��8�����n�_��,&I��.�i�!a/���,{�I&��E8	��.,j�:_�eg�3h�p��s;�&��dG��6c˱���}���Ŋ?>I1�9V���D�����/ë�!�{�g�z�;��U�߮vG7�|J�7P�U¿Uó}3V�y�����>�a9J��)}>� A�oz�<��U�J(?{�
Qp`�ZQ"j	Ru��B�ݵ�����>p����	|_껨�-������`A�k1�����e0rr�f�9�w����3 �W'N�рîd��)94�ȰO��ԙ��9��f٦c)�:�dA��~�;���>�O�6�:|�6� .q�L�sc���<���eՏ�}lO$
�//�v�E\�}$��1n�I%���MR�q~I��P�n��E��k1�s;����G\$�זY�l�wf�k�;�L#\/hM49�L��8��7�}[�$����\w?���	l�2��)�Y��c�^��&��Y���Ma�]�X�e�C�YAu��/y�[(`�ߗ��T�O��Y�d�@Q����"�ԓ-�u�oV	�u�9A�7)#������l	�EB�6sܞ�h���J/�Y��g&W�.ͧdl��R���@�TC���5Hi`iD*��O�^��O	S� ���"�?#9b�/��d��]��vEi��4��Y�@�a�H���0�	���Ā����/9��Ym�_/��QIQW�����F�R	�T9̱�漰�_�V׿���e���f�,�Kz�T����;Ǳ)�GX]��d�}���!�g���޷�����8c����6��΋�%��1|����0cg	8΍����jl,���D#�_��;�d#V�ε�b<[��)�<;띌JǵW.ۡ�;��w�	:���8��څK�8�]��}��jKS�(v�lz�u֫pܽń�����}B�@\fC�B\���Y�a�	���u�8_4㶶t�V��$�t��@CSV����D9����-�Gi���a!ʒI:B̠����*g���I�wQ���ګ�C"�)��&�w8�f���eju�Lh��%m�[d�x4���E0#��%�	H.����ь!�}���.���~X�����OQ;��܀Y��vq�!�ԉ���-���`��D��v/:��� �ƑPɌ��;���H�7�
��Yi�\����#]�6UW�)a�5
�!���y!�٬+��oȢ�����^�ō�x�B*��C>]wMmFԚa�\U�ʩ[�?iv��(Y8���b�x<>�[��I���>kZ�a��h�Z���s9���u�� �"����n��_���+���B��o�8o
Ջ�w�M�婽��Z�;���ݖR�����*%@���C���"��1��ש�΂/�:e7G�Kr������3���޵�8#w���$;��3/���[]�p��-�1,�ឧ����rp4"��2�Y�X^�w�I����f
����o���d:��c&�B�1R�{���*�skI�ԚֲQ����@��iʷ�V�aC��y���E21�qvQ�$p�I�@b�[v��(��4X!�� 
�x
*>�'�T߿xE܊m��3�#Q�{#��+M��*�ŗ�+P�l�Ӊ����u��s2��N�ړK2�A�>�*�_#d�	ʹQ6/��j���  ����k�u[�c�� zp��i&�o�ɝ
m)����[8���_;�H�[�:�� �p���.�w���Q�f���;��Y��9�
�:]��O�$]�T=E!�,����H�9��*=H�����s)�
�h��GR2��n� E�_M_���Vs����kr����8Z�nM	�Y> t#W,�����U�q�-��\j�?���ʊ�� !��7���IMٟڔ܅��ŭ�'��{�axH�W��jH�����ɀ�-���Y�����˫��)m��=���o�����:�"�.!����t���1���fF���Z?��`�	��6���C���瘵��4�{������-3�$<p�x���.���F����q%���V��{ L�8f(r(�p����yZ��A ���;w�P� BU���<�0��l�ytӜU-�9���T�����و���ז��B�B{NF���01*ȉ��j��m��d�ߝ���%�En���E�ށ��l��9�U_�e�������l<�0iYB��:�蛐��֡�G�]��6�JJ���ld�k>:���	^[��AEɥɨ�yJ��C,�0X���Vw��a�4or��-�
"��C�hز*�^3�@V%s��ܜ�/O�x����5�\-�=o�x��m����QP��I�װכŜ*|�"g�:������ul���P�,�T�z)�f/5�l�>{G
@7��|0=4���Ҡ5o4FPotZ��N+��/��dm�@��DE~���[��hk��3�T�/׭�C4�ɤ��:�g��@\@�	�e�}�+.O�5y��t����ƫ�,-�h��*�n��i�/��w� En���D�V9�D�1Z�ak�m���%�{hm��T�7�c�+�`O2���+nu�����JW�k�&�F`j�69�]�g��M�ހ�G<��{�zP���+����=�%$/<H}u#�-]��J�v�f�7��4c��l?6��ֲ�M�'n��|(\��LF��7�~�� ���UB[�U�ɼ��H�V�O��>��N�����n-���w��-��'l���[�WR�
j�m��s�7�4x~V�i�7�u���ȘX\q�������%Z���]���d�%n�3���E�����-*��V�t�ϔ���W�Q_EM# L�~I��l�T���LAxX�"ʼ��OCFc��o�p����F~!�㢀B{��Y���^��� ����2[�/�k����D�N��x��E@�� �qd�eȟ��-%)
cE��᏷�.Dh�I����G>�	2��g)���2��u�B)�Q�7���n�w|��!�g�i�P��U�!ϼ�}�� F�����N�����Źq��"��	DW��G��W�"��]�K#)D��|�`h�2vA���i��7�t�e���Ҋ���G�6K�q�n��|�/�Afw ��/�<���xz�Xw��� �Em6C�~է������n��T�R��a�'��\�'\�Z�6��߲�3el�[`��붿uE��i�Y.��Q&UF��^�jK�XJ2�%6M0�ƆY�n��}t!���:�mL��w�Y]j��}1�*^�2r~��[1?�+I�[u�u~��b��f�A�߳?���s(��2�ˡ��[3�|�A]�d&��'ũ �z�	6���QDY�%s-�_G�����c��x��q�qNw@x-��O�9.Ho�J���X��Sa׵!��c��.͡;��[�B�0�A��B�e��d2�o�����|)o���D�zϓ����]�5$bᵖ���{ �B ��w�Æ��ux� 1v�;ґ���Xj�!�7�2���ݚo�b6O�'�쥬�� wK�o�;�	�3�lN��PXy��,�!u�Ā�4*����h%n��������y]���g��Ƹ	E)����É�W�*�=E3�xd��'͹߂r��%=��l�.i���TSC�1�O���٬�6AS����I{B]���~a"�kU�[�3���RW�RB�Ε���M�s����R$׀O�����1��KM���&D�s��Yi��SVy�������|a}Ldƭ?/�70����:�I�d6<�f���k��:�rAN��l	��ؚ� u*U�r4l�9�5B��J��$}��}��[��V�Q�e~���&9���O0~���������G��̟��,4��v����b
���q=S����TD8��'R���q��?"�u���w����������գ�@TjH�j�1�a���c�}"�Q�o�*Hp�n'T����x��������u(eSnѡjF�%:�����r�|��L����A�3ьA�"Ql�'�T֓9����M{(�������<���l�/�f�	׋y����h<�u���`�GgwWu~���B���6���V�ƍ�#�� ����L��2&2Pѝ�9����4�j�ț��VF��
�������8U'^�$�ld
K��H�$g�w�CE��Af�,{݀��3�N�_�����ay`�<�:VjK��_�m��]j<���_��J�>�ƥ3�L�y	�e�oe��s�H�TU�;h]��
tҶ�K㌒��Me�����r�L�N�&r����(�"!t�3 M��� 8���bñ?�7:DC!��Lʹq��☃x>��C�<-�1�Ĭ;%��g�٢�Р�o�m [��;�/��L�A���ԕ�)�o�g_�Z3�Y��i[ܦ����_C�o�!���B(�`X�ys`��T���3�%��lɓ�.�����R�q~@�����@�}�|U���̐&8M�3������4���]5d�^���#�Mn4 !i�����0~&F�ܢ��z��Ͻ�J>����f����J^�HP��i�i�3�M�he�����"���;�
�ſ���$��S�|�Z�\�Z��J��e�A��Lt�3���G,�"n�8/1Z"��auy�CmW8��:I�#�|�x]�"c*f�����9i/���"n�����>� !��/A6�E���!|�MK	T���Vh�p��l�30��>]8��˰΍I�mn�u/�y;�9�����'�"-�{�f�-z�R��:��S�N�����usӁ�
?��'1k��s+��!�f�l����* ,���zD0�I|�N�*
��E�G���f��^�@�W�@�+H����F)�:H<���gH�!�,r�\�7oP�����pDݴ������\�8}��o`�g"���}�ӸH@8p��5W��c�̷���_H�"��}��d�ih0YhOV�7d/��}�Ī $����\�5��^~@�4wz�Q�\��+P|V |z꾝u��1�95��tER�H�;5u����Υ����ZP��Sb>P�! ���I��goz*0��31�Ά��#1?��%�����-O{�^�*�,I��e���+f�I�ɠ����s����({Xg��y^9�Ҡ��^w�X�~#���[���תP� �^��Y�y*�C"��4�0��vқ��Ü�RB�.��B�c-�W��h#�D�x����=g񔙏���,N[�������[�4X*Y��h�~�Wξ��{s���#�%Oi�о$���
{dw�˔ˎ�7�k��&�j\�_���FP�Zʜ��F8�p��c���Ͷ";�q�9`�7��W�r� B�|ie�D��9�~`naǿ��S}���W� �>��I)�Tg��@j8���Q��O"6��?�Z�����Mq�_bVV�9TXT,�ʼ��ij�-E��Ԉ�,P?���XEX�hh:�O0��d��
>nX�]Fˠ���APKZx"r>�-�GǶ@�Vm7̌|�@�f��m�c�F.�ag.�H��
��O�*��vp�F�s���!��@�H���7�pd"��<�[v	?��r��h%��BKC.����w��1M�hơ9h}��nz��U���$�9���F�//~v��V�h&�!;��gFv���������t��_/�����z��0���	����_a}�E����>�2�u�7�כ[D��t�"N�<�q�/ի��vZTb��h��)a�<�^�;	4��Ll7|(|M�T��wY�T6�"����^�h��%�r�����:�� ��Dz�&�8WhT���5}A�d4���o\d�M�~Y�"ɏL��7���.�;�hĊxu��9�@��c���
�i����@Y���Ŏ��8�2�ȩ��A�?͓f��u����z]���O����v�E�<�����yHb�u�#F���<�z�K2�S�Iy��̬��)C��-�$x�`R��|	��&������K���[˪
�se4{n��룳o�d���T�5+�Ք�����p�����n� Y�ϟI<8�gU�k�"Qh�	gY�gjh�H�r�b��S�c�p��5�n�nwmD�h� �L(��eQ�V����V��=_��R|��\����q�۔[��睤�����nl��.6A�%��Yh��R�j�.ce%�E����i0��3[��Q=M7hn ���z�`�5�\uwK�E�ဳ�L�+A��H�����Þ�UL]P�r<s����@��l�^�Ӳ)�5��ٽ����������a����*r��r���j����"%�>����r,P�"�����\T�D�H^����
+?vpd5�g�yo�-��޵��RT8��c�j�s�FC����>�ԛ�W^>�m�;X�՗J!��/���=D��&X�GA0ˡ�Y�$.H� ����,�Ӧ���=E�U0�:��'��/Z0��/ӳ�`\�E��K#�(H5uV`�� ,O谖gx����]�ɾ�Ğ���sl��+���Jp,]�p<�I?7��w�T�uD�qf�q��I�M�pe�P�Cr%�w2����-�e��������B�E��
"�#�g�����}�3������qh�3����+j�G�����������)C�h�&�GN���]�����Z�/�Eb;_��I�_ᦿS�!Qߟ���=��v��Nh3�F&@M��PM�^�ҟ4���[k�
��y�WG��δ�2tm�x����A�a��=�1�e�R"���%����.�ڂ���w�{5�|�icB1�����~�8�	�zyg��B�2#ߍ��� ���y���]��I��o'!�8J�W���0�)���IQ���8ݛ����D�4�$�d>��i��3k&I��ީ��k���բyV��b�͘�z��*!�Xp��=��FEA?β�UW'��3�����I�|>IHT>�։���JH��n�[`w���0cE3�9dK��'��ꇓ��9֖�_�w݄t6���Y�0E�3����f�=8h��T��WV��i �޲h���8�@ԫ�5����X%D���Fr��ІN6��R:m^�Z�q�?ʔ& ?٨�*<ק ��cf�~y�hT_o�u/zT�熯S$���m_�(���Ct��7�����������3����Va5�	�p��������Uؾ�:I_����ǳD[p����s�uf��USBŕ:F�9�	�7n��Ϋ<�e�N!F�~�H��:�
,
@��Y�wM���/)����>]�|R5%����Q�N�%Q�Z��u.Q(��Qm�dE\��U�,��0��>n���v�a�/�Ia��4�;c=��q�\)�i���V�)��=|慡{G�:|"�j~��V��-����럶+袏G�g_������0���o�P����4�>��K�G�=��0��W�Z-6c����RC8㨑\�X�2F�����B���f-�t��O t��y�QU� L+dG�E�n*P*����6�x�2=!��!
|=�F��n�l����c�������W�����xQK�d&h�9l0l.�Tp��g���.H��9e�v�st�@��a�$"8`��}��,Ù�{��9�}��u �ޞ�� �%�g�>!�+�%2�zbW@��켲����KЁ��ɘ�/{�`	����z��B����{��x4�R6A߾tV�a���C����i��Y�G����]Y<�ʍ��:!"�����4�����;CW7!54�R�Kg��H��|�LEy�c��R�X(�UK�a�k��Z��s$���{!5"��.N�ͽ�m�����|�ت/E2��'i�t��Z��zOڻR]3з�����޿����������g���u�M(2Z���1��@�q�Q�����݅#|��KY���CR���Ĕ��r���mqDƢ<i��,�=�^�Vla�����Q n��zPی��.1�'s-Q��儠�a���nW&� ��SÓ��۹�ܦc��:�#�Ѫ$��&I�#�#�NjiPTR���A�g�-���DA<�BqO&0���37%n�^�	[���N�
'���=��8�
_��¨(S�k׻��w���oO0�m���A��Z������j8�����'wi:Y�{`RI\�7U�ً��V?7�&37�(=g�,�09:Mo���3����F y�|I�h�3g��A����7yCInE�$9��DQ꼑��3h���8A�R�;��%%2D�Y�C �����y���J���M����ι�(��h����=�#�VM�fJ�����X1�<�T������f3~���b��Ҫ�&�X���`U�!��帵V1�Z	|`
Ei�(��Z����'��9�|����]��l��v���}X1�޷�p��gד��Gy�L��)������f�ܔ�!!%+s��V�8m7���vF��;H�L����)l�Q$O�i�
~}��錃k ��5�����/�悌����Є�=K�nX�;�~	�'[�)��j�W��o�ް)��bL��о5�޳]A��s�����Gؠ�Њf���K	�h6�Z��F�|��c��:�[�iwEu2h�ڒ5�3�^m�2�u&�-k�W��Z�i�/�0���󱓶���23��l��GƧ%���K{L�ϳ�&ohp\�ڤxXœ��1�dy����N�׆l`6�b�h�kJ����ǖ�é&���5;8U��mu��}��@�̑NE{�.RӢՑͰ�fr����L|����z"���؉���[��z���B�Â��6-�8Y�x�PCZ���]��`S �4�K�@�Wo�VW����4pS��XOE}�s'�AD;��ؖ0yթo}3��Q��~�Xꌇ<} �� �D߽
&ON7�L����N��P�C�A��8�W	��~�Z?�l?5K��H�3rə8�<ʭ��e<�����=%�y��E���ӹsE'�䘛����ྱ�bI�"����le��J���~��������l"m����pA0�
9�'�t\'G����6�#֮����;dSH(���:�Nz�o���G�� �Y\�O�د3�VC�C,��������f��S�:+qH>�u-�2+d����j��=ؘ՚?g����,�x�=�?Ӻ�0�ƻ����Srs�߶�i�u����l��Φ��L<����9������`b�V��ȣ��+�C2,5#O�x��ML/jDn��QS�����>�s3����� o���'�kc/�F{��}1����ӹ�E��Y���Mx�<���
8"�\��Mݢ[�4�/�.]��G7ul�Q�d���|��w�xԂ���t�ek��]>���$]�x)�ܠX���BO����?��������#�'�b���������{uS�Χm /�U�`y���$�*Iuh)D�G�MY�l����}n����<	X��w>���U���D� ��Msn�ɪ�� ��E��r�أ�j��5:�?�w�IE:JĖ;�%�òj�_�'��;��7C_��g�P!��6U��$q:���SL�VIDp1��ӡ��k̭�	���4�C�6��Ej#���ű�7z��"�<p�q���l�K���P�&�=3�I���y8r�YBu��U������]|?L���̽����e�c_^�u�&����9#i��)��̬��ᖳ�V�m����1���H�z�r\o����ΠB+���%��a����K`ω�*zR��\�K�ߥ���A!�
R+���$�j���#��b��P�f3E���ם�b[ï��l(Ж;�WF��9�7E�r���-����7���->
�^�f;c+�
g��@|��Yo
�b���g�H�V�A+<���t��6�m��۱�E��t�o	p�d$[uÅ�?�ְ��B�@k��N�t"ҭ&�c�*,��U}3�;�R7�>�f�+��!�:չ��?ٕ�c�%�h��������s.[3��+�L�a3�Z|?|I�T5�F6��Q�b: ?�A��^�L��d�.�����S�4I��R/H����V�xc�6O\��J@~�����{T�acX��\���Q��_���31?�a ����z�]8���D�iLK���?�wT���i)���ۓf���u���ΘB{KI�w �Q�{Z��DY��X�'�^`F	��G��c�k����t�[Y��A~�JF��b�İ��,E�v��h'�9�"ޓ	~A�|��l*֤����D{].��F�~n�f�����\;Z�G�����>[h����sܜ�p��M�/a#/�#��f��J�F��f�������܍�]M�Ͱ��t�h� �\E�Z�V|5�~X��dxeN��m�)����4��!D���0�d���1�5��H-3�R=���UW0�� f�z���=>;��.e�3�G�}ǫ3ay�T��\��-�<���6���[���:�U%4!��Niv�J8�.�_�6��ɘ��.b��2��h&e�j��(j�>#)����c�B�%�Pm�`�
�1mm��?�%qZ:qi`���yf�ZiJ��X��s��GrW�:뎫�#1���2�������
.넲����M^�����2#S�Z�M�`R�Bu Ló�����2۳�y~�Ov�L�)����@K�<�����%e�Zڍl�p!xm8�_�\4.D�����S�����
� (Gǔn `�ҳܝ�%�r�S�`�Sõ^![��a?УB�v௉���` h��B�\k��-���o0�^6��)rP��g��(��Z�=�RO�~�]�f�69�tb�a?�=�v)&N�f#���ͩ�iS���`�Y�Lcd�78��A���� �V����9����{֏�_�&�?Jˣ����x�8#&�TٌJ%��Z��Z��O4>�
����&l05�Ӷ�"Ox%O$�(��g�gEe�fQ64Ʋ����r��J�c*�j�Y� t(�}�B�#J�*����������%I����-���"dV}h�Ƅ.)���z�G ��B�+�1����AM~��GD&#!|�_����EŸ�C�J04�<0�)��u+�$\;��u�S��&�?��gk�a�d�VF�r>��td�$'C�@57�1y$�eQ,.�9�Č�rK|���`�K?�	��O+�|���&�:�Z�Y��WM����mF��w���[�5��`K���#�>G���G�rE�*y���aId򲘡��*����$����5����2%M| p�BS��+��cJ�l7Q͇P��[C��5��za������è~��ۻc�H2]�Yh�$x�C�A���N�o��Lt�;HI�������� �E
3�N�x��4W�e(�`��&�������S#>B�Ha�ŕa�����-N�&.U����O�ӂqx˩����-�z 6��Vt�xN!Tsv�dZ�5�x=ᘱ��>��ł�lD���4V��� 曾L��ю����8�� ���ߏO[o}�������t@6ȏ򺝈�m~�hk���ru�;g�5#M���p6⊱��x�2�Օ�5>�)<���E��i��r�<��v�k�A�H�?eBz/M���7�-h��o�Ek$�:�C���ݫ������w��f�Ϝ6�e�8E�<ڟ���E��PHԟ���:�W�
+���dF��p�*{����~��3��kPW[ 7�t|��r[�P4G~�`���2;�kI�@�>���%*�
� �#�N��f��4��$��iˡ��Η6P�Ci�\���@ܡ?�
�Y�@�<׮m
x�R�?�q��$M�i����ry�H�&!�Z1�`�$&D�a��b�bz���sT���z���(�͛���A��)�ǥ#�x;�
a�s>��S�'�(�{t��*T<��y%�h�Y�/:���'���kwL�H��$���������g�wZ[�$rY>L�ܤ��k�p����B���쐣�N�XV����M���GkfC�C�"5�v7�^�����=-+p��bRE_<�z�3�k��c�����|�A�L�Q��&'_uSM�\�����"����M�L �����ӥ�Lr��� ��Q>�X�M�p4u�C��A���G�2��`��3�Fz���pQ˧f3(���Q�T%��D�d.G�5��s�!H�A�����DZc�����VuFx.�-�D����t����)�i��� 2ݒ��Ѥ���+V�^�|�9^o~�������e6'`ZP����p�2�l��[��y��ti�m�W_����T��>'������4��:M�N�[f��47�๮�VF����N�W���[l����f,.��k2 &
���ˏ�>�ȷ�<t���д�E9i�s~�o�g���y
+(�k=C{����pڏ�j@�����R���Y~�p�V�8���)K�ʇQ"�uk�1ݸ�tE$��7G������Ή�����U�dbk���.@�B�U�Q�U��[�F�퍺�D��ٻ����fyK'c�]���VhgǺ�(j���h� ]���p+Wu�jNU�֡�^��$E�
�VA�:K�@�'������&�����xr�"6n"mJ������	;�3���"�o�[-P��&�S<^�IH�{��{�Bgv"s]EG�M�QLXG������,,^Q��؄3oz��DU)�B&\@t�7�0�k9AN}���l����-_�w���I�ً��s�5\� �p0��ڕ~v�)�j��ڸO�b<%����dG"�
�8K҅k�h�hf&ե��& 6~M�k�0������AN��;71e��!x3�~����>K"hVY���?-��npG�-9�����nS�7d��c�\�A�\"߫�WN��R������=�����D4�J*xÏ�	��C��Me
�7���ۺr��#oW�J��ٙ��)�G�K,xw�l;	�3������9��J��yp�X�g�v�,�����X�Yi$p�����D��lU}���Fj7ｦ�&��fk�ȶ�s�+]4~��67EC���̆����"��h]gya���Y
�Y�d%K��y-1hmy�Fe�r擆
B�����V/os����W|9t���?�-�1NS���j>�x
@����6���2�q"�^�J�,������-�����Me�D���S���s�,i{̺��&=U��1oD�g�I�������m4�_Q��c��X����[Xh��� V�j-�n��Yd�w)�ߖ�e�'��@��JyE�¬��jdG�ұL�v �H�h�g�wX����QR�������2uZ��e��!�B�l͹HyF��7s!�JO��+��Ƞf�i�Z4�����Zq�dC�х�1��F�OO�L} )�2������&��0����/L���- ��+�����i�"���Z1��P�� ��Ƽ��9<�`^��=�5�8ޚ�}l���k�1��S^������I��*���h�\ÌH}ф�r3d���o�p4���gx�9�3+FM%HY���gw3#tC�W8�a���`$�I�l-�N�"zW�	�[v�w�7�� 5�}�Z���O�\����[�}���-��w�=�N�]��e��Xnɐ
l)$�T�T/SHD/���z�i0�%�ќy^B�b��Ex58O�#q��Y���z�l�#]� <�p}R���ؔr�꒺�)�w��� ��pq0Y�GO�$����@��t����7,ūr�Z���Qi����� G
��W*]��	��e��:��h�|m�/5�﹟P��S�u�	dXz{\ �
9i�u=���(��m�h� ]0,_`k�R��[�>�������D87��a���鱽�!��9.5��}^U�k��Y��3�}[�d��Ϝ�?��x��ΎM����L1<�0c�)Uo�!S'Pk�yi�� �G�w`�ǿ�Z1�����{9���Q�FC/�fm�D���1~���;����*�����n��ב$�����Pș�cc=)�K��|��H�@|ݰ�<��Z�D���SIw�;.Vj]�.Y��;�Mb}Y��7
�����tiG���H���1�%GgcJ^�ytn��砘oL��t�eOn�$\*�����Z.De!K�Ir�o��'k��M�Rk�ӎ�c0�H��ظ�1P������m�{�&�c�(
��B�x����^1��&��zhˤ��I\���Sބ���C1}��}������	x��=��2�5�O��7����l������pT@��}�{�%EէN�e�lh�:+��i|�X��7xYÉO%܆����2"���]"�f������E)ms	�2
���7Wm���mҀ�쏛�����YړYk	�Jezm�� u���P ����Lc<,�U�g�;t�C��8Ř��CŚPq��J �p�>U	4ЦVH��y��	�y����C�0�й_~�QM�'e_���$�}�t� Z2��˹����"����q;��"ܕX
�t�KU�w��uOՕ���$}Yk�61~i�!,ז*� hK-���4h�{N3ŋs�z �S���c�6"�֝8���Pgu��6K��">���.�#�f�t:�����_�X��X 3�sq��lb=g�4���A"&{�W��<�8���*�h!ҷxe���%L-}s�_�MD��:s��w��W��fM[�����i�C���8zJ6����P\�x�Z�Ŷ,n��oC[X���ve���uS�4�p��:�$a�ȝ�o��g>���M3<:���Mj��-k5 �X5��q�����,��b:��-;!�?�)��P\3L�[4Z��N�o� ��Uc�W�k�"��?\�r%>Q�^�j@�4|�E���]h�2�y�;��q�^��v=B�_������;�R�H��$�PJ����U��z����}k~A#?@��C��zP��7����ڐ���+o�jX�R��<����[ɯQ��釳z�B URe�N\�&��f��2
��>��m>,/̅o^�q-s@p�Z@@�����U���M ����#	��Md�RQ��@�(�����ى�&����q}	���5'����][l�oX���Mm.{�@Gn���b$u�_@�'�t(��ºwKk�J��rꔊx��>)�s��� ���pp��+���zAO+��� ��7�n51�;����D#ȹ`dPj�-p�u�<[e�e�-��mK�S�m��5Ǝ6��O>�� �+����c勻O��?����J�f�us���O�؈Q����]��s f���>��r4ۄ����0�Lwq��_���ݡwS4^�W!��*�i�9�<��%UR�.�MQ�+�G{�u��i�﷊�Q	5�����9� �˱��/���U+��59h7o'ޫob԰}B�'��Pi�Q���C~�Ƅ&[(�YJ9p!$���S�Q�����g���pc�_W�'~�,�F�"R�}����q�*0A�lo�7A�7��]O�῁��셶c�w���D��CD?�ig�	��ÚAKk8�~�޼>�P�%8�k~�ˏd8��F�TՄ�Vy��|��n[/I]��1( ��q(kB�=���QE�}R�|'c�F�;S�@'��%&��(`td��u��2#~�ٙ����0�[�z	����Ȥ���g�S%�!����`�0�=c��\NE]�+��l!o�}��Xz	TdF!�p��z�(�h;��l{�D�ϓr��B6^V?<�e��h�f^
�RS�K7|���g��������Wrˢ��89��#�P�d��%�c�+t7�	�LӞ�9}�j)�rx0I{��@��}?d¾(�m��21��q��ÐKfcc�[�9Ì�y�9QxC�J������Ƭ��E��m��4)�rh���u7���O�[���/w�Ș�u!�!q�WP:�~��Z�楞+�C����M���N�>��^S�4�l��2��2s(�7�|r{�;>�8�F��κ*Ϙ�\+RG�E�k�#��n���=����r.����&7��F�c�����]����(���l,���\�vs/�����q�L��zz*2���I(߇��\7[�k	[�+�X#xp7E�b�C��+O'���ȋ܂�%�8����S��T��w���I��qG	9ZG}y�DR��*тب�cuS����}g��V��K����8
.��c��-e�q@N?	Ց��J��]7L���Gټ�
b�p��8%6=�ḱ���{�H�X�IAӗL5_y�"�oz���}S�=LEGT�IciB�}�[�~LY[��,��{A�\~�=W�d��4��]�����f5h�䰜��E4i\-�e�O`�楳9�w�h����8�:�-^SYcL���f����q��#�:��^U�{,��6����lȢ�w�s/�{]1 ��㍔�u�=��)'zSQ(�+���S�]���Ws�r/r��cm��%�,G��!>�>�g�T�ݜ��q�Y��њ ��(=�>�g�*�'� �7�N@N��b@��j�c�|7u�W�����\춦tΔn�}_.7��y�B���vt"�뼹W�և4}�)�w��PDY�ԝ����!���}�g�NF_g�&z�����؅��+�N�M]�ЌN�O�}}!f����"6���IM��gŧ��{���������l}"Hwa�h����̸���Xy�u�0��[���n:�wsuyZ�<��ﮪ��r8V����_�!��9�!K$ئ X�l]gDK������J׭5-B!�D������a���'����x�΁l��}��z���N���ֱޫ�;N���q�;{��i������ &��T��תd�����
�z%�N�!x&���L�g��Ӌ�MFRؖ>�ɏ0�=���N s���tE__֓ЛPԤ��F�B�e��s� +��*b��]q�V�A�����`�gz03/ˆ��`Bg:�``�4���R�Q��Q��E��QM(�����I�������n-��'���Q{i~�<	��]�Ȁ��S���Ti�� ����T���d�N1�i�u�ҩ++_vN ���|�)���U*,1fVe�./��U;V�T��k�����@3��_1'�cGWb��M(h(4�YT�m����±[�86w�o����O���D��jpQ���a��C}e��X� � �A�e�'�#*�q"�&	H���Bd�"j�����Ǥ��i�!Ԗ�an�/�M�(�d�|�9�Y��@�R���S�/q�m	�!��Ю4 1�Sa^p?U� �җ �;v]�j-�UyW�Y�ܑ]����VJ�����C���;$Zj�����:2*�
�"�Z7�-ܜ.0�Kv�\��Y��ߥZ3��o�Gth��k����3�O�wg�_ûf��;bJ��m��X���m`�0�,��m�x����qd r�O�
�aӾ������N��Q�U:�v��l���������Hg���ص�UL��\��ʴ��k,��7l��J�A�>�@����G=a6>:��o�[��y���2��wz��s��Ӎ�`/����|Ba�G���p�W��l-��:L
��B�zsZ�7�{5׻�IGv�+���?�G��(os� Cv>/�E�M~s��	����S|KZ�O���كd��` �,���!�p��ڬF��)���ƃ{�
�5y�[,#H:�p�m���(� }(�ф��f^��H-Q	<��'r�极�vV�1r��[Xj%��3�_�tlh� �Z�v�-�5.���B�j�@y���N~�V��$�����*̏mm����"�6^M6l���H�V1o��͊]�ȅ�^�d�iov�[J�崕Z?���N�@Y�o�&pJD�Ii����tT�_�s�G��%�Z�桪w�m(��\�P3��^���x/�ű��q`�ȡ"Њ1�X�f�?���e�&�,���Ŏ�����ع0z�/Hࡖ�������X8s�O A�l_���2�r�����6����(;U��FSJ�?L�����_�@���M�0?U-+�Nn�J1jd2t9
�Yf�'�$FHH�%2���MG�E�;!���I=NH��&�%}��|Y�U�����d�J\����3n)��X�B��/�3T��f"� �($�Mp	~>����4��{�Y������Хֶ�) �R�B�����a&	F,���T��j��D�r�d�@D(��gq��T���B`k��&��Вɂ���fJ�a�ϲb	!��e�}�7�"��+����S:�\kBɼ�L�H�{�
��G�G|N"�!����G�1�f�eF���-x�ز^G����2���� X�'x��K4��:�) D���%)�b�#��+Bl�4PkO�R��L��ZM��}��kżP&��Y�oz�%��o��E��%�|A�ã�E���à;'��{UaE�>  ���཯��U�b�
���ȉW�K�Y�Λ(Kr��k��D���S�r_��e��_n/xs����������@��@'c�ژ���}��0o�T7�V'���=��@ܓ*�v*F ��e0wQ=�H���>�,D�!�
�-⬩ܕ���l�+;oّm?��Q�+0]׎Q -o+��zM%���kLڤ�Uh�	zl�^\���Y�R�D�ON�j�������|��n|� R'<7��x���#�]!]"�����,��a�w�~��@��Eq�8^��2 1��'��,�D�-��r��U׬�S�@������p+N�|:l�'',Z�Fc���Wߎ�Vc�K4��l�)�4m�R���kb}"��]/Cl��LU�1WIk��~���!�Y��[�[~����������	�۝����4�R��E>5���P���z�G��G>��e1�y����>�dիP[�v�j�̡���pg��w"�T΁��/P8Ni�wף��9%K�=b��KۺS(�����L���1BR8W|3yQo��ɠݣ��4V3���K�*|�b-�F��Eɰ����EBKf2ɛ��P�	#���5�<��a���QlX��w� � �pZCw���=��?��(~�p-A�I�����Eo��{(����`�?�K�P*�u����$����Dl�]��^�(C��z�]k
}���m`i�P�����A�q횐��S��揳[ڠ�|Rx�Pw���H>��<�]L>��bYQ�����_P1�{e��J�ڮ�v�;mMב���:P�Ŭs���fW�xD��0���	�$�q�2��g}�X��^!������*���(l��Z�)�Wa����H)����{{S=׈B�j����n�ϵ�9��ك �_S�V ���\�m��"(*H"�Q{iQ�Ϡ��a���� �FT�t��|z\͍b�5`���*"[�j\N� -�����F����p��^�w�U�Ye����?�)�r�_�t�<*[���i�όW�u��w2�/?�!	H�O{P�������My��`h�'��"m��˪#�s�Ԥ�E�B*_2u���S���w�1�"���y����Y�o6��K6�7�2����1�D�T�z��W�9!��g&9{`=�;�'����g:�R�|�N~6��4)y���n݈�9��c)0���#F����!v	���/��Tk%�!�����W9����|���a������i�Y@E�����{W��LNQV�A5��3��>Ё�R��O�Ⱥ�^ا�jgSd��d���p���0�^^J�H����[�!�OC{T&ˑ�vZ��L;��)�n�� �����yv�L4��l��p�`r�^�Go�l�|yzi�͒$4¢�v�� �>���7�}*��d���Wfd  �
۫���_�E���5�A��u�D6}��lj�����$�ϡ��J�O �kr�Ao^D�i�A��y\�u��!e��;��)�z��Z\eorL%�Wy��4����K��!���.qj� �Ɨգ�jp��3�nR���ZfG\�}��"v��j���p��6�"��))����p>ZV�Sm '�@t��퓕y�W��Js1L2Sa$Os}:x�>�&��!Ϝ����ϟ�XZO���f>	�=�hqT����	Y�Ǧ�,�9hS`~W'ɕ{�F������w^�i黁$:e����rAo���=T7K��.m� ک�"��:�]��h�����艩
�2 ���L_sQ�P�`[ʛ`�2����3�!��u�r~K�ᘬ��e��h�d�Y��W3 ]#��Ɖ*��]���
PC���9�h����7�>��M��[D�[�2�I����w"�6r����� vN��8����Z*���c��ޤ��V�wo�͝�4!^��,�C��N�pK �kn����͞�_���(��Kr�R=��u�qõ��O+}cш�R�鄇����\;T�����m\��ꂒ�n<2�j�`��A5����%�����>,�T@>����˝�P�%�
	�ꪎk�9��^�(v�^�����G��^+��"��FXw
�?�5Dt�19��x��V`!�p��A�N�ne�@�'�7Yʌq�,i�����XO��$?�!�e)˷�H7��=}���º5�Q8��Z�^ H�z
=���1�.W[G5B �<]W>�[�ί��[�d�Y�J�d1Y��!GAf9ʚ�m���A-:��Yͬ�G��jz��e�=���r��ՖB
�椉��6#H��PWL�>��g����A��tHu2M�05�Q�X'k�-JIk+�3�]�L�G!5�~����6-O�lx����5��j��J|(�!�ER��n�7�L��C�n�
EX�3ig8~#.$��)�_(��뚞���оf^��ou9�/�����<�2��͓�T���k^���� �Z��S������7ÿ�����	\�5x��a�~[��A</ϣ���C�-n�{}�K��*
^6n����ނ�!IwT�)��H�e�H���\������aM5��c�v���'�C��c%���ȩ�s�$򱻸01P�}Q���Y&����п���r+�т�n���x ��Fŵ@
��T|�=#�
*�À��,a:��� �1�{�(�bK��W.G�����'~�"_��� p�	�p��E�����<&��#fh-/ؠ�d�^���������-].Ch�򼷣PZeYa����"#@�W��af��-�D������<�^m�d���Kg?�o�3���}�9C�=����тx��Y�
�i]��� :o�?�=�쓫
9�K�{A~i�t�
S������W	<��͆ 2�8�ٯ���'��|��N�Lz��KL�&�����0�u�<`�
���2iLiD1�s�6�p;: u34����-��Fd�-$�� :�^B?_yK����Yl��:5L���E3��5��ħ���0�Y=F���_+�ۄ��kcYܨT�_���ý�^S��������iӺ\�U�A|�Y?�~�����Ô�c�.I������g�� 3��{ͯ�������́�����5hr8�W��G��a��2sݾ1z^�:�u�Q>�ŝ�4�f:�8�g�$kS������	!����]m$~Hמ?<&6�2�R��\!Ns�,���i�vP�ÎX/���}w�(�{t#v���8��t��R� �J�X9q�I���)�>��j@��D� ׻�:)a�i\�:�j5 C|B/p�+m����b
V�oA�k�vGJ��Ȅ?��iƩ�aN"��MF��n���8�O�7��=���-�SM�fI�I�U�bk�����;6;�B^eƂ>����c�q.���9~��ؓ{�[<m��P���pʁ	�O_��(*,`k���;�_��{�����(GF�?o�ia� ��Iv!{��� t	7QN�0霘%�p�/����|)�#�l�}i������ ��|��:�`��_��������;$2�6�B�ǹp�F��Ƴ�|���m�!����#|C���W�-Ճ$!d⇰b���_
D���4$T�b�H��߇�ݞ�a�_���Em���9�bY(��g��oT��qo[��/� �f�o|�/Q;�{.���2�&�?[��'�M=P��\�����J����Q �=;M2T��H�o���wz(K�~�e�t��X�-HLP\r�x��|XNJ��x�LD��[��<B����$��Ņ`9��*��DUt[ *!v���#�P���`I���ݞ���lM���X/%����qF��o�:�XKѤIT*��)L\��_�����>{Ք}�ISϝ��iS�R�n딄ULr8n�
�M�x�xXtud��y�h`@��D�������]49�6�0��	�Y�wN�}�6�����.Y4e�Uf����W'&�?=-����K[p�u��G�}sN/<��ClA�HP�&�.�9�7�ޗ�����@b9�p��:l"`��ϓf2�}�U�Wwj�k��S^���a���
�� �n⩄
��pw�ԋj�#֥	�w�(��빾��a.9���!�>v���_����a=��M�] �|FM���1rY����CH��`�m�*4��co�E�˛�lʪ�����؆������Gx����{����:�G3�+K�D�z]�\�c��i���E��ɿ���dɮ��o���Sʸ��]���^ա���~�I�~%�\ҧ�an��y�ю`������Gcǎ�`����/3V"���:ِ'��G�����][/$���]f��@�FA�R�����T�.>�ͺD(�P�� �
+����ۖd�a�x\&�N��~�5Bm\LT��3\v�E�1pa�p_of|0ӏ�cC���bO��sj7�IR)��_�g���0�_��������=tkA,��s�l�I~+�%�}U��q.?QҹL������K� o��J��[)�S�:���Lϙ����3�!i���?F��y=��ج�*vU�n-�ᡜ�&.�;���q�ߓ���msAF^@��'(���=90~S� �w�N2�m�v���®q+$��7�����h���^v���I���0��*dYK�+>��G�W�����H�Ƚ8j� �����f+�!�X�w�%���lIWk��T�u6JKN �&y�������C�X��3~�_)z�rj��(��do��V)�U#�r��]���mC���	�jZ2|
�D*ʩvYv�I���6���E�vP���j�ȑ�����[�e�<W�X+C�.9�=r�\~LM���
Բ���9�{��gݴ:l �_��Q.ĕ��jS��ML�>u�ɽ�<�0���T���$��Ws��2W#C�B��kNiy��&���&#E������ h�H'Mr̤6��u��#�C�d���d`��	^�%.�j0����l��_-+�_@�,�����?��L<{�Yb	����+-��O�^Hf�d������ �qX�&���;��E��u��0ͳo8r��\/����|0�[���\�KM���
���.�����'�n��^�'�!}��I�{�������ucM9
��g�W�X�npS����0w������
T��@���L[� �l���u�����^Vs\S�4�Nq85�����i5\�Kx���~�i
f��nY|
��(�Z��h^�Q���A��\�H=���+�F����?��5V�o����l�@�o%WڰAX|���I���̀t�B������/l������L�N39k���U;U��B���T��)����Ǹ�{��c�o��%o�ަ���9m�Idl
t�%\��i_��v��B�`+�����N�A#�d2g���OF,m�f>�\����um��)�F�Zv�Vm�������NW�$�=�2GtC��$�V�if�2F����ƕ��'p��iK��̷��,
�%��Q:]���6�'�'�H�(�Ҙ�-�TB��1E=��,��%"B��ܿ�.�ep3�S��*��,w�oʹd�*Ӽi,�~�L���+d:��u!�C���������0�N�����c(J��m�(���2�ӣ#�n��%��iI��ږ�L��R��xd��Y�h��52:�h����!ϟ8��aI��!�d��7����n���W��P��4�"S[��Z\����a����8�����Ji7mKu>���߫�֮٘�оQW/�B�<��O�1�o����"N��˅y�"C��G�E�#�emϠ��˷Ѱ��a���^��T��}ZK��^�{�,"��|����E1����*Sڣ��^�h��������t�1Fp6��V�}O�FbF؋�M�R����4��:ѫ9��zo�l*AWUȹ��#l���0ݨh����L�%�pÇg�rV;�zM2u#�3�٘i3��!f/���m��?A, 	� Hd�a�r�k.�,��(��+�ǻ��RnW�**��w^��V�^A~sl���ʻk�!n��ݎ3N�>C�G���M��y[�æ:����F���􃑙#rI�D��bkن+�&g^"�Qͮ�q����ll�N�iE][��Gņ�� i� �rM���s*��a��f�j�&���^��[#�J��O+�j�&@�h��zDFw+M��bڊ0�/𒑦�ʁy.��9#�Ӧ2�g_zޢ_���l�BLگm�kCl��rĕA���X���ڙ�f
m�%�isє�Zg;f�@��~�#p/�(�¿��p��.^-c�4��{rA��UM�'���βr���E�f���6�	�>b$[����Q��m��~D�2c� 7T=h��p�V���:0���n��\�)�uj�PI��L�J�!���<.�[�'��=IH=�[r�8FO��_������J=D���wV��JM*�=�vO�ԭ`���\u`�@cq%�}�X������Ƕ1���v���̗6ԙ�����������s�շ�@�$2��0�3Rp~43�@�"�K�J֯�@N3�TU}q+3�m=������ R��3���-�x5��T�c��*�iw]�l7(�#��mq�G��m�?����f6jd���~���G�SVf��.���4� �b��c:E��ʉ���,s^���_�'�������T��B��Dj�����I��&%����hB�@����¡�b�Q�k����ũ��|�n����ep��2��*j<�NS���܂���Z���NB�5�:U�*������URf#�]⣻%It�U]���N}����O-��2DI8B�q�V�L��hƳ�������2��Q�æq{	����w�
��q����C�%����]��Y��ש��pxZvh7�g,lh���	:v(�C�*��w��z���
��j@�x�N9�I[]uA6{��e���5�gи�r*q�[��F�]Rl������Q�r�i���;�����.��]ZM�A(XY��66݃�Ll ���K�%a��0p�<�[+s�M>L��k���?�~�ܜJVu�+33p����+r���n�L��T ��^����0�:�`���l�o^�s	���cf�d"�	/�`$��b�����?�'�dS#Ǡs�~!h	b�h@�ܞ�g�g6��O@��zO�nӦ��r��ت������g%��B]3v��q��n@�#~Vz��q�$;'"�Li�?e� ���&��_r$�7��>�Fq$��*6/�&������NU���<MTs���[&�A�>��+�x���\�o�C����_L�}���q��f�NG2��@b���A�(��ޔ�b5Z6 K#$�����A2��:��"���&)҄*@���h�廙��m�ꆆ�3�v�t�^у��3��,����>�/�zv��m}A��$��'�D������=��b��G�&����Ed��\2���=|�`�Y殄��b��#����њc��YSV�ή�|f�mk���@Yr�TR�B�y��0��a~�6�D���K��1X��=!qi�娢�cd�b�L2g�(eɰ�<��QBy��S!s��?�; �2𯈩|4�UX�,7�	w���^W3s]GCOWUug�Wve�A��9���E��:Ǘ��֝��Er꾺�\��s������̈G�3�h�����C[ɔ�W"�/*���^,���ڥ]?T5��o��t'��&L�Fx�Z�	��ȥtϛ�t,� jm��0g6�w�+n�t�91����6*NCo��TQ�G��Û����\�U��i2@��sy'ʍCSS� ���f�xA�^-]hhr������(�8���7�sɍK=c��U��9�������t���ͣ�c� �ڬ��h�.���z$��EkO ^L�,\��f����A�,�GXtd�O�Ƕs�!��=Ə�C@�<���ԕ���NmL�p����L�q2nm�zK��3��(؛�Yae�W��O>0z�Y���݈��/�CjeSFg���='/$�{� m��:�`᪫�qQg�K�*+T(��*F�#�.� �g�7�,J�I1ck��R7�� �����ʜ櫈�@��{���Y�j:RJ�
s3�'���1�	�ȟ}�aC&7�ӕLPy)$"�ٟ�"E���(��wamI	�0�,�`��j�ϟH�<��(��y��S���,�X��fpw&�*�L%�j�("��W��$4'�~i�A���J�)x X� m<z���VU�N�]�v6+�y2[tj�Db�)�H�J�\T����sG�7��s�=H����1��2�^���8W�;�n��4u�N~Kh�J���Z�wr�,RB��̉wj;���ڽ�����F�X+6�\�q{�1�/��
&E�P�z�i� �Hy�:v��6i����D�޵_&e�Zf�����i9�KhA��t�_w��m��!c�T��m���]쁣��q
D���P4��"�'>���)�)֣��:���3����&�.԰�h�y�vs9bg��*��ib��: ��g��TX�[�)\���p;�s<9D����M���|LN?S�j����fN�4���	���\�M���=$�c��B}�m
�&�1��Dѭe�4"^�A��$��Es��gy��鮤�"��΁i���<�쉁�ub=-`~c��(�4gC5�@#V���E�T�"�5��􏄧��Ō6�.o�(k�k��^���!�o3��fhG�K�|\^5$a<�l�ݲ-ڠW�/��<&����;E��D�����)�}D%��͊����s[&�HS���q�n~���#�iu��z��D0I�ŕ�ĳ S�ևX%���P�@0�� xj-z� ���]����a�RCb�&����!����t��s��# �[�H�ww�+zwa�y'v3{�����W�?���&�v5������+����%(�6�������5HS@��_�B��H����m�݇�}n�dټA+%Q>����rM+�Qt�F�>�)H�d�Fm���)>��hX�O�x 9s��A��gM29�/H�4ϥ1 �k��1��6��I�gVQ(-Ȏy 17iXUKgю��}��#�9zj�(Fz�5���g���}�y�:<�9�7�X/ɭ�l�3�t�j`�8�#����7o� W-��6�X:�O�l_L���Q��}О���jQ�T���CR�Qޅ���Q���I0�U���ȣ�D��N	�~ p\����¿װϠ�u��+�n���B�W�5�a�8XCt���D�׽FV���@�3�����6���ڞ�2�C�C��̀b�pE
�~R��O�}�o���0i�K҆�L�(Y��r�:���$I+��*�g�p����2<�V�;�E}���Q~�ܒgjq��h�u7ԜR��(�J�� �<�8G���(7��X���L>�a��s�j��V�B&�,{;_Y��^��	�g�c��|2p�|�\]޶~>@5�4�i3.��+��c�� ̛��4����� kh� �5���2�wu�I�S.yv&��_G_F��꼑A�k��ʏEKw/F �VD�S�b3{�-��ž0��c�^�Yi�z��|��������3��"��g����5����ք��W3Mkgl�g� �����:%`��݉p�B�u�_��>2y�?�J�3��mf�c�
]l��G��7N�]`��M�<�<=X���&�;�9Ͳ�32RS�o�¼�d����]srt%�W.���3/�8>8$��{G��.���G�/]Y���~M�a�Dn��a��g��� ��(�i�tN��� (�]C������~H��o 8]��^�����n�����tY��v5��uY4��J�VA$F�M�#���l5�"���N0�D�q�e��u���x�%��N�$�K���[It�>�ҏ�gT�I�z��G���m��(���Y2%�!+0�b�1���63(qʹ�@.�b��K�r����$ɱ>����ۀ�围���V���7s)ל�i�+f��vp�^�zU}@��:��}m��$�V�֝O"����%� ��+��!�N��:���@Đ<8@�DcE^-�C��e���_r3�Љ��Om�Ղ��(;7�Kc����+��`�����[��ip.�mn�iz�����|�v�ȃ�F�q܆kɫOA��<�� u����(��m*��C�R`/44:�%�J��� �ފ�����ٔ!�I's�M���p��1����������5�F��r,�G��2��7�������ǑA?�r�*��?r�P܅�G�L	����{W�,ڰ��|=Ofk�ǿ���W�,��22%=,���Z�욫�mԜu��k�-zZ{s7��A�'��V/��櫢)pw@��Qs��0��LU��N�R�Ƒ��2��0W�����@��g���3^W1ظT[��U���>+4��;qI�9.��}�U��7�sőf��$_����uq�,*�������J�� ����{�6�G��U8#B���Y�.�dJG��̛&�cl��������#Uw�YE&̆��f&	H��$=d�i��^�8���Q@V�#�'/'�D>�i�����/aq!J[p]�^�����\��E.1���ɳ��\�8ֶ:�!���/���TN"���$i)�
�:IKĬ�6BB����l`��^Ug�_IV���y�h�Ε��f�k��{"g�O�}�}ts�D=�E����h��F�:ޖV����k z"�����-Ś�u�)\|���_�޼���/�8���]�E��1��i�?��t2����v��(�$v����,� =:���N�B��a��^QWI�ouC�rKg�
��CŚ�`�r^;`���d^ \�ŗ̨¦2����Ǖ̊���D�N-�yn��ܕ慬.�d�14sU>�Hs<�b0�1�����2�fhF��u.�	�Y?�}��i�FS����� +]��Cp{VVW�iݫ|&f���2�蒽��z'�{�J�X�U1�@~���6o�K���.�?��p% $Ƿ?���DE5Y7�S���OU3n���wQ�Rc}�G����<&LN0u!H����������_֥�M�/�e�xhc�y��v�RZ�];y���EtyxI��E���ԣ��f!*i2�$�FW��c	<�k�#s�fY�%��xpKkT�����H�����Tn�� f��Ѵq\z��F���i�Yõ}b�!�,�����0�N�]�'<�,�A9l�)EX��g$�]5�6��Z�X�I����O�(T{B)6�W��+U���XRA�`Qv���ī����
:�kO\�W�14؟G��:�L��*4YfJ��r;�h=�C�Bhg��v��O;ɯ���"�M�@Bu�=L�+�1�\����a����P5�B�����F�T Ow�j�9Dr�q�e@]G=/s1�ð|Z	� �4u������)2���Yͭ�r#��3 ����E-Э����	�M)%��l����s��i�Z݊.bv���d�d����O��<��[���|����_�"�2��c�+����a4�	�#���&�|�ʢ�u`���ˉ� P�NrAY�(':��h3Rc��8C�M+�954�\}j������9� 5� 	(��U�'<Ç��[j��*�tlU./ҙ��d��UG@��(��D��*���Q�j#6F�@u(��Ts5t@�Lf�N	r���v�Z�����������I�:	��iiHjy�.Qr��h@���	�!t6�����p+�fzE���VJ��_�|=3d����Y��ǕY��3��ӆ��^2���u%�H���H�@R2���8W�D�6nt��?:	�p�R%{kj7��,"�a8�-���cn��A�4�*E�\�S�o�����x����%��^�'{<���ʵ�!������n�bBJ��j3o 9����=NZ��eG�ߢ�=�����eG]=s}�.������s��z�*O����7���h�)!~j7�'�]@M?�\��J��-$�q�ήsf�At!��p�͞:�g���x��k餭������ڄDBS.؛VWY��#�
�}�rB��o�5Q�&ovh�0�d��珊S���K*e�dHE����2F7->�㌛5DV�vgo���5�?�,��+�^K�C0g"ZAY�����p��K�i��7��U�)-N'Lt� [��Z�e�vivp�+"�UE{8�1`�`lg1ɠ+9똿I�P�^~��� {	y�	����_.٫3�W����x"'*u�7?$�L}�� �"����xm����p�ǊI�X�J�غ�Gg8"5����6���,D�u�ۚ�Gq=7�R��9�2��Z���n�Oj�T�$]U��KǺ��E���W�V�N�j�4F�-[N~UU�ن��B��ֽ�uN4M.�BOY��8�A��t}75$�P7�#�7���7�LVf��V>#�&t����S1�S����=���wg�9�{@�.l\?**��).�Q϶d0˸�r�m��e�s��~�lY�7.���6
�V_�`B�zC��dlFh�G��Ӕ�BW����El�u �/;."$�A��2�.��?�
��T���0H���C�ҜU��\�l|�����)�L?��d�b�{����Pye�0M������r���Ҟ�E�0��87�����ti�U���O͖�y@���/4+c�5�1�s/��bJ����KA��`RM(�;
�'`�+1t�*D(����#?�aZ��r�T%<n˲Z�?�yy��!R}��O'�%�	�|�r40�p:o��A'��F'��[�C��0���4{�)q����آ�v#�T#�U�/�7�%,_�M;��2Df�OG�L�Y6��(!���C("i�'��4<(��ڈvNXB$����N����C`]K<m
�w�E��y���q���"��T2]������r�*���n:�!��Lin{FzdR��rrm��(�E\�s��W���J�1e�go��b;�����y?z�~��w˄W���Lȧ�f�;��U��?�[�M.�z�#l+;�u�;9���7w�n���]����&������\�'�(��W�2�)�;��K�������D�^4�9	���P��^��l�[�8�����bo%>虣u�Z|����}�}�Lw��̾��z�b����u��d
PF`z����Z�x��B)K�{�}`�9U�����S�x����uȣA�Q�/ �_�)���h���W����ó�x�~��y�> �-O\&��F���` �t}��	X��P��/��Z:�s��Ēg��+��|+�}��\� ���C(U��:�0�F�+ĩ�Oe��E��!x	@<8[:d����,����SGY`k��z���9O�C�͜���(�!(Z5�BYRj��L���)@EZ�8���F�I	��_Y��l�=��M�PtP�)���B�r�.� M��7����TN�SI�8�g]�aC�$׎���
���6��4�J�xK��~����Ơۮ[?kL%d�D�P vd�8�֦���&X�$u�������u���ԑb,�A��
��$�{@y0Eހ�I"EV3\栆�G�P���q�AMTu���|[i�b���(KWtF@�h���x+��5Ⱥ���f�[��8��ܥ�!xМ�\Wy��U�KJ�P�4%eu��G^�l��n��D�Y&��g_�L��Ձj��n��i��<����s���u�H�H��$t��ܧ��������:K�/@��\���)|4��Q���]��q��)����"by�KYڭZ}B�l�V��0Z�^TED�0y���7ļ ��l�x���rb`.b����lo�m(�����s�Q�����OR���	���O�|:�3��N_��L�UڪQ�����j�uEu�W�Mpj����fkRB��Ͷ��i� ��P�BJ�6�H$�x�h��37�T(���㑨�������c��F^��wT�\��IL� V|ޣ��P4?In�Ք�$��Ad��f�zqw�$���A����0*�`�a����hw�c�Q�ߒ2����P ��Z�wn��*y���4�W@�f�Sܢ0����JX�ɭ��!����?E��E��������A�N�ew>!?.�x�_%&]?}��T���$�_h����Z��mK��'�y��;mu{�Et�4��$rJjQ���ym0��'�s��~��B�+gT���~|�f^b�I.���-^_��q��.B�+�]�7,Yf�J���o�� )�'yP��92be����e���.�����機��̈́��[t~[R���z��ۭ�l��h<�msd���"0�&P�D��ѷ��ܾ�v�WKX� -�q�)σ}	�b3>�>p!�3�pg#k��K��ƒ�-�@�l�s�d�:�\ҕO��G4�cn����7m����G������B�^A�.1����*�Ǭ�n�ԙ�n��9P��mcG�D�la'a�C@���<�����^��e���䮩���=ڿ� A#���4w��38�R H ��\�U�~��c�	Eг8��wN��iƷCz�ᇎ[zҾ>~�3Z?�R���L:- � )>M�H�v E�G�
V�7���H\��ZJ�AW'�~�f���C���!F�����Mg���`#�V���y�b"K�YrI?ş�+�ǩ.���JY�Eg��eW�ə;ٚ�.r7"T����#�M��Z6?!���۷R��f����N�����b���{�B��wt�"��m̰���6�뿜�}��}�v6�*q��d(�dU
>�/m����#���L6���n�] #3����U�݊�b�զ��D�|�ʎ� �)QCZn����]��Ea5>��F~La��\�σ�?��/g���UD�P����0��=c��0bjwp����Z(3'8�_X�ӹ���A��n_��Qy8��$�-bԓ�.�h����@��<��0e�G)���;f�V2X,��91�M8�k絨������$�ǔ�1�9���"�d(���E ��'E�
 ��My�U[�Ϝ�Rҩ�ؘɕ:_�ab��p�kx�dD�P�n���3۹CKnv���A.�d���V��	q�s��Nx-_?4�?��M��\a�h��	d7�$
��$��E�tz�sa���t'��0�&ߐ��hS��y�EEp6���&$��w��g���ᜐ �Ьc����Y��IX�ɣg V��BͿdMk
{��k+Js��D�ǥO���8�&͑��K��#�c������J��v�� ��⬈h$�TM�RcgS1A��y��*��}���*�S�d9h������H�!��NY���x9��:&��y�zk7VDtԻ���u&��b�
�cUv�˔.kl��A�
O�����7�hV��
�nT�v��Fk�׎��{�$��"R,@���.�� yX׶�"�i�V��� �,p�A�a�e`����U<t����j��F�1�Xa�|��rN�K�nY@�I��ld��(m���7��F�K�
����E/0/XY��K�����kӘ�Jy��\��{�d~�1�XqW�(1�ѣ͏aN�֏8� �j�>�_�1N��#���bb@"�ӡI�u�O��� �E�R���!~�'�n�EV*aū,v�v�8/��5��k�?��Y�@�)Y�n{R9YGm���0��� ���S�}#6�/���x��XoC��R��K~��9����f�
&��
pGC��e$���ۄ1���?���{\#Ϯ�k݅yL>J �v�Q���f���Z�B�VP�c<���5�O>��q�.폙9�;�'�I�5u�üxwPU#�k�w��Ra+�������ߴ������
�6�G@N�$����VX�q?|����%9
���/~�?\%�rO,̺�{Vw�d���CPȃ/����0��~sg�/���E��U�5}_���m�U��=W�����K�dz���3@_^�Z�V�2䊻ٓȃ��<(��s|cF1b��=����v ��seJj��mX��]'��g"�i��U:RS�e�m��룜��B�tk���M-���e���*���[�l\"b���bRվR&�u��P��p.�08t���c�MɸM���>�j��u��߄IѴ�F�����r�5vwB�>K�wjL@��hZ����N�z"�1��ՙY��n�a�}V���4Û��jeȶ���+���=vG����+���h�Oo>�vNM�	�E�0��xL�<{	�B���1(U%�ď%��`����
|Μ�TjB̆ON�3=�h[�(Qj:-�q�1�NG�>�ѳ���޺���"�V����{����9��ϸn��c��c��!k-�MոO�,��Y�c��T){�T+���+j��h*�
S9<SӤR�f&Ј4���(q����!��?L���GB+�VB4.?�F��x�R���2���$�����<��=����49��y�y��JquC�aYݴ1��SHɈX*���˴��
v}�E�묶�Zty��#D�H'��m�ǃ����D|yB���>��?�����X'U�{6�J$��D�*M�L��0u�!]Lފ�B�S�0l�5VZ�ct����A���ߕ���J򲢏8�m6�!/��RQ�.���d�䲴��T�	�{g|+Y�l�!h�t��BP�>�x�F`h3��ã����� ���"uWwI� ����M�{V8GK�q�:������lv��R_v5�c�s>�[1��������IF?��|:t�}W�钻ʻ�bz܊W<j Z����DD�Є���i���/�f�-uh�u4�&hm�|P2X�O�7�T���]� lzh`������mE�z]�o5�uѹ�S�����-t2��D�g@��Ӓ�H-��w�*m�Th����9�M��YƟv�Q�Dm����"!�eq�	N���A��$g�GB$����a�\���~�H��۵{Ha�`�!΍��6���9��ر�����!G�g�<!�>wE��z����1�jMe��F���?�btH;|�1d~���eȧ9ђ$m	�[ٯ�?���͗_�������E���K~�q$��ۃ�;9�%�t;5��
��plo{�љ�����s .��X��	�e;J�^�ƙ���䛮�Ϟ$��c
;�;!��}";X�������%���Z��m��^�K�7��w������˪�ՖՂҰ�/ӿJӐp[J;<Z77e\��Xת��ƕ�G☵kD�'���7y������x�2�����<��	)�'�b�-��}�.�+Ř2J�T-
5�����rl�y�Nߤd�Ñ��Z;?_�0�}I� oL�������L�6�Y�WB樚O+�D�4.rp���
(GX���d��pA.b5������.;��T��^j����?�jIմ�ّ�2�$A���7�jA����~�_�9j��v\�����R��93{�c��~��Y
�'�<y����&�J���r�c�<ύ:�� wH�~�Ma���ާ�ZPl�űǒ+Ew` "�Q*-_E����d��Q�P��f��.�W�C}���g�&i����x��~��x��>5#��� @H+m���I���"���vWI�]ݔmJ�W�8@�����U
jp�x.R��~��ʔ�-�5k�p�l&����U(�Xx��ת���:������Z@�<Xh��T��M�o+����M��zz���7I#+`>����4��D4�U>�L���%V�(%�7�/ʖmF8 �S��U�yOޕ�jH��״�X
m՛���|�7+$[�6��w�U�7KI�C��ܗY؀�q�f���4?�f���2����b�o���5��{���e9V��h_p��H�K���Z�,K:�҅ZQ��x�Pg�6 ��A	���qj�a����Y��x�s��l����~f�񊌙7Vs�C�@5G&��wđb~�~$7��Y%ۨ;�j����P(���6�z��"D�M��G��ںL��ro3QO���T���@�N��.z_� &�T!@��;��χ(O���j�:��W)��u~ 4��iS4�>���A�	ǈ��_q��!a4V��h��Rj�2$N�[a���h����Ӭ��� $����ۗ�ژ{KY� ��*ų�j7�?�$h������!s��	�a��oA"2��������b��g�`J	��^�:*�ӝez> �rv�h��#�w��#$�q2yЏԴ�enN��A�Jk�JY�2�W+�0�pt���9*�!9XN�/�����H���j�,�cSwS���[� ���dI�x��p��3(��O�|�VvQ�S���9�5�A���Cf� Xdo�p�z&�f�팍RS �L�l���*Ή��*���H7@l
��:�̶�����>B`�N��#�ߣ��B����ɒ��Sc-"�r9�9HB쾹�Dk��V�{�0bi�渴z�D��3̚"�j 
==�X�Oy>����N���{�Ԫn����ʃu9��1�5v�Z�P���{���Z�� ZmZ݈��ˉg�ŝ��/Uk{��ݡX �\���i3?�wt�J��p7�p糗� BD�����VybP�����ʏi��=̊X1��;yv>����4[;E�@�כ0n�';�6�熈��?�i����t+U���Q�����ȯ�#}�
)8\�$eNe�W���GQZ�:��Y;�n�z(E�'�mCI��+��1�(ŏD�C-9�&�rs����EV�P$(k1�@);�����>L����TU�
�M ��9Һaz:O��TM/� �ꨰ�����$*�KP��<����E�����P5�xf37^�X���;�����n��<�F9�r��=�	මٙ���Z��<{H!O�`e�� �Ui���=�{!�r�D�^6w��^�A��i�I��
��7	O`��г�[���s�����7�K�w�n�0�ߡ��ã��_�'�����z����7�B��a�'��j��3O��m�F����pm-�z�`��f��P}����1-1�r���#i0rVy��ʪ�W�v8�1}��x��@��m�sc˾1�r�P�{۠I���^nw���mrx#�%ږ������m얱Y�t�[�����ZDm擑S**&7"�[⩌����V���D��À�(�83E�Ց��hW�(֟T��d�*�4�B	0S�e򫳭M���PjN6, ��s��T#$����qz,A7R���s�x9@�Wd"�#�d��͵��EoI�,h��
���+�[5����Z�^2'�ߓ�Q�>����j��.�<M_?$���M���f-��N-�����h� -6<�h�z{Xdg0(d6�M�ӤD}��턫ɫy�<:۞N�?hs[y�&�����l�Q���f�W����}5�Y�$��=?�9�'���:d5ƴ�_�S����?q��u%�o�B��q�QDKSB5L��u�É�|�J�*������\�G�`�M@�L���SZ�6)���pm�?U�*;(���]�B�Y��h�D��L_�_��[=%�����P����l5)�pۚE���DQA����(Kk@�6uJ�<7?2�x��%}<�=��w�-tC�I�� R���2��8Ko�SV���L*�t6�X��z�ܱ�{&k���7�����'��AL
�=3�bR��<�Հ����r�3%A8ԜË�e�ccV�c���s'����N�R��6)�4-<�P=�m�q��n��2v�=��<�K>�$�7T�P��6�$��騥R��0�>�2=�
rǇ:�-���kb&�y�ͳ@]V,)�����?����Ѥ9�Tq�`s���I$��e<m8�&9RZ瑱�i؜[.�<���9}�F{�z��:�-�E{n�ߜ�V�D�j
��|yu�*������������xH�x��D\��N>C`sE3S�k�k Bz"�\ {u�3(����"�u��.������n㫐�m�a�k�s����|��U��� �X�1���x	��ǒ�E�U6�A�E�Ɍ��<���i�w��z����-{���U��H� �o蓠�坁����A��8e1M�|(���� Ű���ݵ_�k��!������`4b;�{��O#���Y�+��t	W�$y�L���$�`	�ꦓ��VIN���Sе �~�#t��_��W��vQJ�"��gUD`�}� Y���W��<��3���Q#Q}g��Jꏯ$����X�xF�d�[�۫�^]z�A�[s�ӿ����>*��B�K��.OOl���Xb_S�L�f����N��!S�%ݵ6�u�q��{۽�d�^�P!�8�I(��0k�{�J�ձ	������̦s�(,բi%�GBR3��>��RC�NE�E�����iL��͌�i�=�F:ꖄT�l�dN	;E�2��VM@�I�y��T�T��h�U���7�~�+ɵ��,����U9;�y����$�Z�6�(X�.�n���3��סa����6:!MG�N�m�K���JZl&X$��a-����Ă�m~��8C��U�*����ז�Q���.,�!u&�gP�����먵��
���م����]r����}?���xC!3'�e�ȋT� 1$��t�ىH�|N]�@Ht"enG�`�`EȠVX�d�mf�2u�~I��״�8_�P駿�4��(�$���m7���0I��	k�Ѷ92��MmPH��"+H��a��h=���	3�E"#}�`���R|vK�)�Tq&b����}���}]Q�([�����{o�"�	�3ے�!M>��2N6D0�{�)�H����9@LA V�/d���rl�<_V��*�&��D=�����<�l����p��������L2^.rF�YUd6�Ri,�>%QyuN��Q���;��~d���j�Z{��Ȃ��v�߀@N.߯�����C�:���e��8�O���`E�BHYN����jN3oW�/��/4����J>�3�=#b�,cܢ�L��a�:^��AjBC��Z��/,��-���f��$X�
5:�ͅ"�9��ؙA�Q�~Ѕ�VgՐ�O/F���� r~4j$���gH��
.L�b.��\��#/9��gd�H21	�~�AZI��]n��.��.�'k�]�G?�\�kU��ݲ��[��Y��!���,e�0G����ŏ뮠�R���ݖ�����9q4$�Fl\+�1�vE����d�$��{"y��l%�����y�!A�Q')*���"zbpKkC�T�� �%��v9��&44A�2(�cUu��TV:�N�,?�xN��r�z�#�Z�jmdd�v���J��m�*Ċ��"�k��b]V�:�芪��2mx}˟G`-}o<��N������l�A�B34/A��50(�.8,��Ž��*Tt7�]�ȳ�3�&���{�����`�kM"����*b��:�29mq���,�f{ہ�FAp�D"�D2��p��e#9x
rh)�`��g�[Z?�3���l�[���	��*���o�D=�Z�YB)�q(��q�<�e� ���x�Ѿ4�+�&�ImB��x�R2���c��Ԫ����K���q�A�n*Z;u0���gYt�hJ�*:���)W�&Q��?�)p�uhB�`)<//�B�Ge�O�ybmx�>�F~��E9��{�B�M]4Ho!�cYXڻ8u|�T699�J�e[D@\�'*��_`N5�6�%,gK���T��sH���`Sl��+��6e�ԫ�p4�nw�z}@gb�?�(������~�[���F�tJ�5�����o^���6'>d��Z�g���Ǵ<��YxH p�2�e�؛z$^J9ٹ+��T��;r'M��٪/*ƀ�NԜ�������AC���M��,Ʊ�_4�N5$6�IB��;;�IJ{�T�n�D����l��87�;H�RȾ��T�cn��>U4�9��~�Y�db�"�L��ݟS%����+�T<��H�d�O��E��b=r�_�T��v5>��ɡ�Ki�	;�rd07w�)���<%��FF/"T��	H��/��Ֆ.��D�\�#U�kЗ��5���K��s�@��7)�c3ZW�*k#�T�J�r���fd��y��`�a���y"x����AF]�lhN�C"�$I]%P���?��|�nee����jJz����r���l�~��ם�Zp�(��مptG��x#q������G&�fJ���ɬ�Yu��Ĺ�b!�!#�"�l��A�'��fW�9�|�f���:�SyQ�_�1�q�w�]�����̈́-3�� yڤ/���.r`^�]���PD��U�o����#4�F����L��jß-��>�ҕ/�q$�GI'�1dV�F�][�~�c��*�NM�x��e�s1�d��Q`7�H���SqA��z���e�"Q�ͥ�V}*"��dR���?LQ��>��pE����J�x���ʚ�~�&k䣫R���5.SI��}���ԘHMߚ�\�e)N���D_�ߒ�ıEP��æ� ���SP�b�;|�@�����̨A>�y<U��B�����;�a$M����\2�}��O��)��,O4��3�]���*�I���b����V7�\Ѡ���G1�ͽ���Z�G��5:
%�$wr`�+M�In�jb��ٹ_EP�l��a��� ��2ev�Śwh4��p|y$�t�n�(�������dzX��\3�qԭ	V;OLA��n�(�U�e��/�=  ��[�N�( �ɥr�����=%d����]OR�Qo%/$"(m�w.�ך�!!��C�J�iCY����x/���1}g*��W�,sO�t��mȁS����Vr�/�H)f�M<�jz	O�����o��с�66�:������	Ͱ�+X��+ Y���y��#GM�iyb�?r����8'�lB���@�y�z�gfE�u��۪"��_��Ʊj�It��j
�;���m!8�'����f�������0-)�#�|��>��+|Na �,�����ϊ�mN�iV�i�(��������~�����U������� eC�qqN��E	�m�*͆�Hqz����XcFY�gz�Ͳ6��;��K\m���B7W�u�޽�Jq��߅�8�x��S	+���n2�#��BF��(2��`��R}'/����3\�2`!�%�0���q�?��o���f~���M<)az�2�|�{5KA[�zeE7��ɢ$BQm�j��g�b��Ͷ�����C�Vsk�H�Ė,���/�+>�xW��i MC���(���2]�A9�_��m+,|[���r�Z�O�^��){W�"I8�HL<e�E�{.�j1�z0�JfX]�xS��
A�V�S) qx��Q���E,��L�îtu�y����̜$
��s��U'��x��[��BC�uI��Z����:�7.��;�*�_ �1�S���6K�\�����5�/=nW�T���1�xTrF���}���B�ZA!��*Q?o��c>5�&1v�"���x���v>����!k�Ȃp�1��Y�s+��[�1��c���.rEN^t�i&H�[��b ��?�qwB8�7��'gTߋ�!���Ц�B������v�IH���}zR�����=�y��a�齆*ّ��<��h]�)�������L��M�B9ܨ��5@� �b9rL��~XJ{�uA��ʽ4��7�=4�ԽZ�ݹjP�|&�B)��g�N5�s�3+F^;�GhC`��Ǽ�f�@�F����S�a�����fS:�^�KުsC��S@�txw�8Sj�,��2A]«;�e۴���v%��I6�vk�R
q&�&:Վl��a�몯R�t~V�6Y���$d��T�%��o���Jt�K���?��Ґ�Lҩ�g���mcv���q?�Zp��l�$?���J�̆���`�0���RJ�e�G��E��r5��P�+<;�|���c K�)�ˀ�'�kI\��W����bM��a�{P{N�:o�e��Z:^� $�.��M��׵�������Hz;|��VŨ��gm%_�r@I�g��!aO�1�~�<77�&iYj��锔��qT���v4\�p�.�$�<(��n��F���n8����s��&�2��7�)�Y�G��$��Β��Z>�[x��>�ē��U+6�Y\݊O��S��;�xB�0C^Q���c5t,k3�Si�)S��ꊏ�����m+��bc�&ʠ��!���
j�����*ϒ���\y��Ⴙ�|0"U�+���/�kpb������K�e1�J^m����1E(p�����{~z��l�D��WJ�>5�!���i������(!fJ�dJ�E�@�9]o���)�2]�K5���$�w4�v�������D��92���̦<o�Yb���p������0��m��I�X��P��b��ܽ$�S�{g�3�_�G�ک�`d^�4{�=��*��x�d~QS���ڞ���k$Z�'Bx�^�
HV���B�52����zib�,:bؾ�s_~*o����B./YDՍ��:vX/���VE �}�{�����\��kE3G����?��
�Y�>9m,C[Mo��s(�A?q��V�_&�����^��<ʙ�3^Σ;7���ɛ7�i�n�x�0�]���o�;�<�D��ʬ��̖�7z� �-o��gɀ����AS>Y�n��Ԓ)� ��FI�u���){(�鍿KLyo��k�qs<Y+�u����n0#H�n��_Q1��9���F}Pp���*���y��+���+�=��
J�*)ו�����m�ޞF�����@�5�-�LHfV1p60G�[�fG>l0���-|���׺����(�Y���ME�f�`ȓ>��G���
%�R�k䒙�/5ˡ��=��g	c�O��ƣB,'I�`���J���OЏ�ʸ�R�����n$4�to��D�����&\�N=��&�S�LByO^��@�v�D�cV����-p��������� ��̆�H������ҧov6��q	�����w��-���i�=L]�\<�g�˼qls�^�8��Y߮3���c�"���R�u0��ϾFH8>�L7)�D4�x��E��ϚW#�[�I������!�_o&��#g�r�����E�Q�L�4z'd����l]� ����g:T����둾/�9��{=�Ǔ4+q��Y*�;�.VV��~�۩Iܸe�h)J��s���50��'&@�9SdCv�R��w[��c;ϧFD�26�R��7�u����$��Db�>�1���"*�k���8�Lܸ�D��---��g4/��+�&�ǹDș�}&�ȏ��6g$.a֜u(N2�`�~̸�{���&�'���5�ұ)��<I\�*�S�B$S�1��f�nɏfG3�3ޛ��^�۽��S��n�T��3,��zn܂0�ҁ�b!{�r/v�+��˩�5���֧��V���`����4�"���y�@�t�m$Z��M[J؋�7ρ��L2��l�-F�y��N	����a�m-�P�NZ�?_<w=B�k'�@�R��j��:]�Uf�Q���r�pg��9#��M��e�t9�p�0;���<Z��;) �?]'��6V��=���F�p�&��px���Ӽ�R���j]lC?�W�$u�
�>�j������v@��F̧_�M2H��hry>�fۈ���o�ofMSja��Oۖ��m��)���[�]I�t��rj��cp^���+Z�90�8�aZR��*��?��FGM�	`ߑN�A��yu�l�C񹳭7P����-F���Y��������=X2ӿ&Ǣ�?�}��F�En�X�dP�u��W���Z;ˁ�cK`�+*����14����ՠw[s!&K`7��C:M���W3U��A�\A�e3�V��	����;���~�H	lr�����o��jן�^���(�1��デ$�� Ȭ�:`��f��V��H���e����'x5��z���h��y�Oe���jٝCm��%��l>V���d�ע����*�R�9�Zg��=��Ub�������˔��k�Z']�Ǉy��G�5�����5�����n\5a�J�i$ ��@�� �M�]k��rJe�W��y�BZL
l�>[=bǬ1��A�pL�~�W�W@�{ԣjZw]?pJC�
�c(�s/�
8'U��~��	���O�z2�cϷ"?U�@�h�%5�*� �ݜtq�tN�#ݡW e���ܚ����=�Տ��^
 ��+^�=�}��y����e��ZR�7�ڋ��n>0���!���(�֕�|����Ļ��x�[�Quڂ���O/A:���?r�*�q�U�J]�>�*ު_��ɮ�e�Q�8 �kb�������H�P]V��B�v��D����а5TWq_�O7������l���dj�����$�+��z杴�*)c{Vq_��İ�2;$�گ��>]��H�$�1.����Ys�@3�Ӭ��fGpjB3�NA0S�Jt�H!kx�έ3�a�Iy���\������v��"�\M[z�P�x�2��d�|����<��G�*o1��KfWԵ��Ku_�yk���4L
ZÉ���<�X�4��x�EJ����?��#!_ �PX� %�*��!s��T�6�f��ط��I��,�i�5���.|>��K�&� ���qB̹�"��y�"r�`����c
�B��yv��=|7�&�YRM����dzT���{(/�'q컼Z�6��H��z�Jx�v���@<��~g�Y�8��W'�Y����$�� ��Ь�4��Bu{,�D�(��0yEV<[E��V
cZ���K�ϛ�
����j���j��]fB�f	�oT��(����1�L�trW.���8"
��.���F�J��d�0^7��;����
��(vVm:*���3ߴȍ�
�4~$c�u��QT�g��さ�Ju���"�c`��Uy�{x�����'@������cη�̽Z��� �V_�ݪ��QVE���d���\�*y;q����z�R ����S��ݜ���ػ��i��������@f�M*r�+(�kU��DN��rK�F"a��-��]���Ƕd�[�8��l[נ�d{ �ݶ"#F��r(��$x�O+a5��nH�E9��F����[b�1/W�z����@���K�qfb����Z>��q�����Dl��6,{��x\�0L��Vx�����զ�Pr��q��?jz3"�Hr�W���2S���3S���Ø�>���L���dx�'A��j�UB������'Lv�����tE+��%�K�%���ɐ��~퐛'A����ZDW 
����UX ���\j)�d~ �`ٍ�PA ��sqM���k��ű� � �t9�~4��~�n�a���hn�9uA��Ʃm2���z~�3�N�y�O�9�B���E%@���^�j���dApw��z�Ѿ�v �p͹��WY�Q�ܘ;X�AIym�n��	�p�n�/�3�U�u?K�<�ϓG�o/yO�����3OaW�B/��`C���G�Y��D��4��XaU��4����^�*B�O���cX��S�a��B��j�� ��>=����G�ZZ���L�9ol1��~C���C�����:m5L��yUE�Py��x�P�u++`o8Ԩ9�c�J��kG��n�*�ꮧ���4�N�U�I�`�K̯��ՊPqT��c]B�豾��i����L㷁�d�ďx�p4�+�f�J�n�;��I�81>�8lS�������L�߰d$��]"�N���je3K."f|&{�o�β|_���x�5��	�8P�	C�R߶\�,�[M{)����%'"q�<�ȶ���֓��I�bk���j�K�!j!����|�8 �U�F{�?Z���ŹA�"��@'�'@�j��p�YI��<Z_�\�Z�bO�DS�F<���}�� ~���˵�BC\��K̋���"Ѧ[y�Ur�������w<w\�&V,� ǧ���<J���t�x%�H��M����)i��5w�x�Ğ�K��j��'<�W��z�J���r~��{d�4�w�;SegN��T��S�`/T%#����,eqb��K47��ޭ'�I::��wf�?��[�Xq�x=���rf�⋍�"���9��u�%U\������)2u�:n���\������.��3�&k�A@H^)�8R��lkᵨ�Oѳ�a�<�`ګ#�hi&7;Qԝ2t�{n�f�ҋf��98���`�'�+���A;�9�W�N4��V� ��n���/$-�Y+Ao�Z�;1L��q� 9��*��;������#K#��jx�~�Gdc��������)_^��"�zQ�Nܴ�Zv,:9[��+����2(~� ����������\�G'i�����r�9|���7���~^�	s6b�IjR?lV+����Ъ �F��u�~OH��q�
�,����N�7G�a����Nin1?MԷ��^�W�U�S�^Ϟi_�Y	}��6^����`�TS�ȁ8�B�eVV��x��#q���l�JV&{�D#�=P��o�0�#S�\���|�O��%�q��o"�e?�_��2���ʠȶn���l��J�i�yc���},�1�E�1ߺZ-�fIr��z�ţ!���w8'�k@�җ�k !�S�����Nel�5^4�������+���|�Ոe˕��'�wSz)}_obٷ��\����N3o�2��u�����h]&�;� �M�&]�k�?N����;�����}ZY~U-�R����1ڳ�I[i��㪼m�^����6Z+T��{�ϼʹw�L��4,�2-]��=H�!��ZX ��Kl�s����e�a�M4g�ԐW�S��o�LB�u��9�Y�����Ӭ�Oиm�gؾ�bHCb�T��0~�?s��n���.�U��ZE8)�#P�S-f���[YaJ�j��Q'��LC90^xA�l\���&�0���j���E�]�<�^��$�yM�3��~3�c@*.Ŋ�����E�C�N��ǈ+��y�$H�(�B6������I��bL1Y�Ö�-C��k*�}�l�~/��f]�[�b����5r��!# ,�PZ����ͨV�Jؘ�6�l�Rl~32�)\cۉ�Ч������wCK�a<c BnxPq���7����Ԓ��K�ݟ���t$t���i ��D ��ah���G�vM0���"�L���Z񪄀b|�1V{7�N�O�lcO���g��,c�{�hθlr��}�_��h��w=R�K����!Lkm��*��w^���Ԉ����dE�В֜M���;Xe�IJb�:� 97�ZAuZ�P�e�,���JZd��^d�T �B�=�1؇�9C n�9�ϭ'��,(A��ҽ��������B���HO�]I@Rڢ��u?Ç���5���
4��2�
t�o�.���n1"tE�<�p���ᄀç�0h�Z�7��.<�8T.��b�l0�ڠ���Qҍ:E	mex ��~v��m�>� 2��(O�C��[��g%� |sJ	�N�? X ����-�G|�nٛ��y��S0��Sއ�B�"xv�Q�P�X3��:5J��caԮ�>{��H!�C��8�wPe��I1溠�h<��R%�e $�!�i<4ܭ�S�Kn���tb"�$̻��l��������
` /����ř����q^A@�t�\���?z��o9�=���[���Tyfl����וQ��4�۝9�\8��mj"u�!4�gw֍��L�Ԉ�K.���.�(("�M��P=:E������ ��=Pky���Xz,�a��Ws�r+u�-�S��E�S��l�]�?S"��+%��������j���,�kCt�Ɠwz+������_l}�Ff�=�4B�����~.��h�2��L��֦o^��I6�Q)�A��Y��*�c�,I�N���!HI���~߁dZ��xH�Xd3�oc������/�0ʶ�E/����JG�6x�&�W�ivo�L����O��i���ͼ�><����(̌RD�q)-8��Ns�b�1]��^��%�x��f�;������P ����Y��/�e��+�k~�l��A��[�v��H/[d4-�"��r4�_�d���P���S]��I��*:Ӹ��}�+�MwB߻aH���u�*������__�w?>����>�l��=�"��p����*{�5zL��H%HN��6ذ"4���q�V��Sv�:����+�F��_j ��w��r��1KK�
�����V�=��id����^^��s��� (���W~�u�mL9�m�\K���T�r��3;`I
�$�Ț���%7F)mG4 �G�H�۴���^ĕ��B���]��S�r��ha�<s�βiB��rB���K!�Vkz��k�\�:���	(��]$|�����j��'HS�4��9y٪�T��q`�Yg����z��"������ct��׶�+�:8xN��q�̛p-�m�-A"a5�ɸe­�%䏧���2ܟ �(��v���QU1=�;#ɩP�قBjǔܒ����,AL�9��N�}k���i��.r�&�t�ǯ�B��,�]���w�7�� @>��dY�*K�!�~��`�x�኱6>ְN �'s�ӈC�s���Z75;aH�i*��]��<�0�t^�sr����ڀ�r;��+db�0s s\6�Yв�(f��/�3�8/��!���\���v��c���tG��(`56�bx,�
����N�*���4u=I���Wv^����cP��Z��s��
��^����Ti- rj��dr�)x�d 1�A�f���Z����p�#�'��d�æa�Vc2.+�3��������M0$~��$�x�O��~��C��dJM�B��c�(�k��"�u���P����j*���t��s���p�^#�:�5j{F�9]ɠ��LF�9�X�2NO-����ſ^�ϮWA㿃��޸��sb�D��C��h}� ��T�ٺzx�jA~�5|�mL`�9s����J'M�Զ9CD�cRT>�07M����ain�Bd�K��v�u<�mY/�
�ņ��1����~���]A�|�2[.~]w�ݹ�>9�
Z}���h��0i��,��i�iHGTL"]�iZ`'J�*�\݌-�&�?�7N�C~���^��O���BJN^����P��wnKM<ߌ.1�9�{C�|�<z�*��2�D�Tg��>�����V���=N��L�~��Wμ���Ca]m���v�t'NfNj����p�)�������U��I��9,����0�v�,G�UWB�"9�����A�/���R�śE�^�8i5�����#��3�ni����;*�~�)��	���*l�����S�F�X_�a�H�{����#�a|y�z��ܣ�)���1���O��&^�l�ɘ0��yK��iD���0ԝ��>����s��4����I�>�6"m(!62� @EBE����xbu��2�c����^i�{:�T%\� �馸ya���Ro\��i�����û@t�̋{��r�S�\����h��X����笸�Zm5��N霟�#{�q������C\���3Vk�!e|����6V�X����]} ����	��?��%Wg�K�߼�wp9��M8�{��Sn]a��f��p�0u;h�ۍ��C���l�`�Qi\s�\��"�$��4������3ӟGӜ���B�=V6��/L"��Ě�ww��L�r�j*��R�8����Hlnq�+N/����t2�&��$�����B1siV���#�
A����c1��Ytl����ެ��,+����T���w���o��c�Ʊ�X�;� ��`T�4��5wU���Ҽ� ٞ-;�{�	�N:m�Q".��>&���Y�~��B����!j>�O
/��/uP4}7�Q�����)��;�׸ �����n�h�\/)��y4�!�&KW�7މ�_3��|:��9�ڻ��e�1 �ڴ�q��G0�W����������j��k�m&������*>U��;���*(ZmL������<�jT_����(��ՁȽ�`�6�B��&¤`pa.'��e7���K�2�ɖ ��G����:^�ʀ9��X5Ā�Y�Z-��qJ\<�/"�l���D5�>�r�:�p�oZ*h�&��PK���
2lw��aR@����e�и���?�x��}	�'�q�D��^M,(<�J퍭��	7%��v�e�[ww���5��O�.w���MDC
�F%��]���zaX�=}H�Ti���̲�&��l�%́i;�����E�e���p*�v߅UU�r�붴=�vQ�����0�6�Y����"6�qe+�(����fZ���M����W�fB�\mԠ���#ĕ���D�Y	(����;����˴�_�c����]i�s�=�7���o'UO-/Ŏt�\¶3�ř�t��┷epo������j<5�=���<��J�<\���W���H�����e�!>�l�?���Bԍ5�����@0��^�o~�Dlf$�u����q�a��� �V8y0��G\��^a�V���K���-�=ݔgp�s������+`�Շ�cBC�z"$�*{��v��Bz�G�J)r�+��B;�`{�L#25Ru`�b���0�҄�?r������A���<�W"�l���`KZ��Ll�ƴ�U@'H`��6�+k��5�7�,�oL�@�?�>84�n�"��Xچ/������;Ks�|%�H�CеMm;?z�pl�~��1��%�8ۥ�u�Ǿle��?�qճ4�;�A*��2a���$��{U䊺��Zڸn�kIiӘ0�c;��|?�q�v����@~3oñC)ec��H}1��el����һ���0-�����E��l=)�:�u�ڧ�$�+Ǖ����<zjv ��������4d�R�.'�a˪�S|}K�Zgt6�bu�:���0S�H����r���kZK^w4���!���ɓ̴�%��Z�>\��X�3�v��S?�R��L��7��v��V�^��־y���9zI~&)��K�Ŷ
�@�FT,�(��G�C�s�h��5(�!�pJ�rV/��A�}����p��ߕ�&I&Id�L�q�u��oD�u&u�����/7��]l�$ɑ�ډ����� �<S��aUEN�Ӳ�%�E��r��P2�7�1/t�Z^BR�``x���,�"
����up�"�i�G�g������o� ���vf��4(��xs��i��f��U��T<�2��s�B�Bk�*�����Ei�؅�|�Α�2M����5#y�Z���A�a�R�����K��+mM�ͫ�v�k�B7^	�H|���.S/�aϷJ�X�=��^[�V�0i<q�xu���vw5H���������@T�a��u(:���c���o��I�wCOk��&�T����RJ�5��d?�}�~t7Wͱ��s�-�%�
&���9���1��νj�P$`!3���wZNA���A��?O��E�!q�i�Y}=y~�$/��י�#����o��!$�m�cGc�/��i� 4J��O�h�-��=<_�t�['�z ��{V��T,86 Įj��c��Q>釢��� KO��H�a4.M���$$�E�a�5�j�����&�h8����� ��0c�t��Un䫍>��0@/������󘁁e������([��I��Sw��񉙐���������l��H�څq��=jF�T���d�ch�D��4�ܾd�b����p���
�x�hc���|�����D �%mR	H�K	�\2.��?��G �?8�z����ZVEq가J�M7�_��M�������U>�rہ$��qI�b=��E��`��$�Ag���h;NYo�ڈ�|��$�K}n3H3���b������3H�c	nTQ�~����P�T�=���n���!�rx%�y�'�˓��������K9��U��������������qR-�)�Ϛ[��}a'��%��h8���͚�,�wө�gQ��N�&�@�*Y�K*���q���RUu�D����K�@Gh���y/�MA�:9׏��!O��W�(�.�S�ߊ%E�;�(ҵ�(À��:a"ռ��{�s$��׀�n�-�� ?��_6e��k(���Wa�c�p4<��%0&��$��7��V�&� ��{m�'a�1�⢩Mvf�=����H�`���*��ps��-`fB,ON��Q`��߽.�Y��B�v�R�<S
�Z��N�]K�ad�!"^A��E��^����edۚ�A�U.�(�u$���t�8.��C�ݒt��'|�����)��@TA'���w�Ӎ�4j���͵�s�Ν�ô{*��u]d�4�;�[	���	N�(wN�I�\ߑr��N����q����(��XR"���M;�
�wޛi_-"�{y�%�|އ�����n�2#h}�V�z8V�+��ŵb�N��&<c0�_���J�('��Ԡ��bDEQ�?�+F"������$6�'�S��NɹG<u]l��s// [I��2���4�o��_��_��g6<Y���7"!芦%:����A"�t]!a�/`� �B��$�d�2���X�s�����%���m1#�)��yH*���k���\�w����
X`m���}��l.��0��%���?��4�^����r�N�3π��r�+@fNyU[B����S��K9�e��HT��Y�5����_ማ9c�]�v�0\Wil�uf٪�A.�}(�)��(��W��-,�_+l�?�BS���s�� f ɟ=�sz1A�z݌��\�.8`	���߷����{����?����ۆ��w����Ѐ�_����L����8/kt�|� ���i�Ȓ�#6�6��@v��$���]�Q�}e6i��|T��uR<�)J��4�jC�ݛ2z�l(�Ս3�8���."���]��rI]���+�Q��J�(u"օݹ�U�� ������h�����*,��/T��x[�B�������Ի`f[��X�SID��ߩ>�?A�w�B�P��K�Ԛ��?l^s��i�¡dw�9)M��u?�@�
r�r0�YR~|��i%�ŅFV0�=^�ج�+�}��O�� *\���*����$x�voؖ7�
�E5�9l� C�@C�F�t�}�������]Lc5@�z�
�ヱ��	f!Hʦ}s�n2=�$���ѧB��;����z*���_W�ɵ;>Q�6>Y�h\3LM��״&*#��-%0H����vz�_�۱���7��%�}���	y<�M[D����E$Q��i����tJ����$"�OfC�1��KHZD�oxE��,x�s�Xy��P��lл��|)��$xWO�puqh�J��4�����J���S�7_��T�]��8���VS�3���Y=a�\����(FY��)�+?����5��������J���.�73~X��j*�Rk��͆�"<�`G�4���y�|{,�Ȝ�(�O���,Ԑ�\g����i��8X� 'Q+�`Pc#\��Qֵ�s��01�u�)�_�_r{�֐���� ��[����R~9�x������|� �r2�1Wѳŋ������ɧ��kȡ�q��C��3iL�rW�],G��2�`z��豂V<5/�&�WA��XVsCB��vb��V���;�Ck������8��+b<��(c�Έ��iɻ�2˪�yI�QXN;>��60�,�Ah"��{s���EZ�j�d`8�r�c�,Y8>d��8�U�д6�X`���0�3֔P�S��]��L^5�?4��<�6��ʾAրz�w+��툾�R��r�Zs73���m�Q�52E����������D���Ccaw���T����|�"�Z6K�.>ÃLO�R�9������f�*;8Y)���8���+�tLػ*m�_L�̅�,�G��9�7(������xpP�En^f�~�81��rs�{Aɏ�3֝}L�yG�-B"�QfP^�G�ȃ�G|��t�V��	������2oc��lj��[��+�a��섙WaP�H�\.��d�#`~�%��{����ܻ�0bz��,�j�eu��C��E_�#g�J�`�����ò���D��$/�����V `dƎ�﹂�B�ٌ�1����Y^t��2�-�Q�Y�� [&5���?ƭ��	��-�д�z���8ƶ%i`����y<��Őa��$*��l`����(kY6U��Q�a�*ܖ;�J٤��'��0�X?F9�����n�z$s Y�f}2�h�A�!\߹?����V��Q�	w�͊&;4��L4��\�	���=�⭾斄41-!�e݁.
?��|��U�k�
��:K���fh��ـ��0�m�!vWw�l�84����l�Fcq���n��hǡ_qL�fd`!k�#�
�UڍXY�jڞX��� |&Fz�+�O큏d�����Ta�aH����|U����Pj�M��U��ZA�.�7N�A-�=^�{���7�oA�.��"r�@"}�'2Q!�;�.!��,�2*�:R�9�ܣ5������+�k���8R1��5�qQ�;�3�/��1��ph�Q(�����6�nKH�%{ӕO��IݹK�ߨ�&��,G�69 D+�*$�h����7�v���c1'�z�ʮ�3nK�Fc�1�*�0m�$O�R��#=���D̠ʥ�<Vjn�����_k.�fo�Q1A�	~����:�1�蛅��;+���+��+���Yب�c���jK��oӝ�҆?
t���4=ẝ�)g����H0l�l|�T'ߥU�o�YI����g֩,�Ѱ�8�S+C������v,s��/��L�d�x/�u(h�ȳ�c��.׉��AZ����"��z6�!�-���`�
�T�IQ�Ŭ���w'��
v�|xT��
�ٚc�A3��cz����Lҫ��d��g|v���7{(��ʉ������4�S�]� ]��y6Ϝ5�)V�0���	 �]��-�uW��~��I=+V�peU�=V�w�ƒ����	�f6pTNV�O�� �k�q�EoG�}�m��<O��qv>�N�j02� ���R�\�.nmT�ޖD'���Q�M|�*T�q���
�*��s�[:	'��tm@S�p$p-��{��?V�#��PD����l��輒N��D�=�h�n��׈�6��lFfX3��TD��H/,����d�O���0���tЉс�ɵ���ȉPp�vI�l��X�b��=O0��-N*�����]�ö�T�<��P�l�(���ݲ�6{;��s�ۦ1Q����U/����7�^n��=�"��^-:�A�MK�.A�o���?�e���D&6�{x�R��] ���fP	|�"��#���<q��2\�f����10���������S�
W�`�7|֓��i��v��򫷈���z�n�Z)�4ؠVV�zE��+-�%�ϛ���J��d$�/��t�MA���A���:�7�����[�QV�`����1{��P�a�<֋k�ev%8�|�ʔ���?E+l���&/D"m���\?P�f>�C� �n�5�g��p���c��mq���ks.X*^���6n�"g�~3q�hGkC���`�2�$<�]
ߥ��$�̨}#�EK�j��&�[f!WS���^���R-�f2	�Xe����>o���]M�{bo��S�UvWlNZ5<H�qc�S��ׁL6$p�U���i!:Z��L���#2��#���:'��n�J�q�/5�ے�<i��s�v]�JvGbq!�g��}.�2!�`�+-��%V���>�L�L~/�<��S�aB_
������:%V���lϨpr�\�-�(�gs�����ǵA\XD���m�/Cd�_v0c}Cq�[���� ��r�л�����dAFi������(_to9B�o/���)�46zVE���,|���y��d�և?��'Iͻ'�C��H]��
��6��"Y_�hI���u�+;�ˢ&��� ��+a"�3�꿻{�cf�	��A��Z�r�bd6H6�_-y�ǔ�#�y׹���-� �ƕ~�+�)��B�8��`�bɉ�R.��'B��!Eh����r�v����u7琚f1�<�V�Ye\��a7&�T�_ٻK���K_��y��mb�!M^>$[M�c�Mg|x�/K<�迳�7U��ޕ�M}�7���6���[�Yl�6|��2��Z~���ɾ�|nܓ�l|��@��Y$��1��(�K��>�a��E�7�����\ �m�
�)�P�T�%��Q?�T7��D�zh���d��8\u�=��4�k7���Q̥w�}�����;�t�c2P��%1S�{�D?3Z}���'�1�D�q7�g���b�%����-G]��$�<^�9�[6i~D}��/ל�V��y��&�� �Z�G.��#��J�e1!z@~D*��hi����1����86�F(rk�����#[�ˬ�/.����s#�'�Oo]]��Y��+�J-;R��2���~�Rk��o���5-A� ����6ĭ�4�֚�S��25���C�| �h��@�rv�v���\���F�|c������j�~��I�"uW�X�*Ί�/������y�O�a	\ڐ�Zp<�Ot�JC�ؽH�����ܠ-���0��l�_WR�Z!<�J���H�C˥��]��Y�s� ��p���'��n]�e��}9%6�B��O���'A�����Y�W��d"T�����HC[7��F��g�{,�w�KVO���ҫ�u�T�'!�?&���y!
|�d&;����QK�%�5��ʹ;��8b�Q?q��b�����<��B�*O�&���V�=4���z@���4�8�?T���sț��a�G�d[ �7�O����x6�p�	rl�3ր�gq#��v��\���X�Eɘ�$�i���
�Î97Z�YyΉ�7����� �lO�2�Z���_��䬭琵ώ��:��X1�!�@���^������pi��#�SD�54_p��/��q���s�E��8'�8~�`�4a�3q2͇S�/g�l����`�i|8j�t���B�����qh�B��r��~�خ�����̤Qa�����Aˋ��E��,x�v�:�j��y�S�߂Ն����au���8iFЀ���Y���CP�-�ɥQd���]����'<��(L+�̕�i��f������Q_yTa��Ř��h��c
,��<ߊjL��/��woOΠ܈Q���� �������o�2U����N2�"ݴ8pI
�̩#��k��<L0=�c�z�TH8'5�������h�N��0� ���KTշOw/����eL0`�4 ���C�P���ē+��ά� qw�w�Ԍ���>��2&):�F�h
��Zc���r	�eT+��E�+#8�rg���|-O���H�����~]!�SB��׶�$������+Op$����\oEAn�4j�O0�$,H��7�(���[b�Lg���w�KoO�MQ��H1�~m�e�b!E�T�~�&,~ �u�!y7DJ�XW륌X�=Ja$���Bjphr���0PO�F����v��n�F\_ݴv|j�w6^��x�k�e	��s:;��}C�����n�<�3����b|�k% �t�t�f�l|�dU���{IY�6��iVK2��f]���Fc�b��x�®)���[[,�e8� �����y���'ܴ2u6,��߬Cߐ�J�:6p�܉�dT<�pPJ ������n֠����sO�!�vn��Y���G5��@y��*��̥��������^�˘=vߴ�'�����0Vd��'�x�v�U,���,�vJG�tէ8%_����A�飚��Hr���߈s�n6�n����iUr��S�淠M��Q��Ze��q�"����)����J�r�?���S$U�_��`::�[@a�9߁h�⮯q��z�c�L͝[�nif�g�� �=�Q���X`�]��&G�*��`0虻�e�o��<���pZep�gN���EjZ=]<v���.Y���:�f��AeSd���`��e.9�����WL� �˹M�ph�Ѥ���a���@�ۻ�'ط� �G��9 m����(�7�l�M�hs��R�s��b�d�D��Q�ss���x[�3a�:G��_jlk���J�_\�~<����0��1}�Jn>F�Em�+l��>7�h��|�$@�T�K���qf�j�D��=R£��j�b�PV�,h b�[���(�b�(�6F��k�+J��AK��1�B�����o�7����t����T����7i�=��%���ռ�U�ғ�*?��7'�˿j��%�t>ߞ��v: �:�4��G*F�t��>��+�������%B�V��BT-r���5ti;��|A���-%\���˝,���A�.��u&������?2&�#�t��(
pXL�
��P�B�ð�"�x�����3V
��1�lՠ���$!����H{!<�s��I1�Zmj$s!� =�і�����<+0b]4֌��*��:���#��1ɝ�܁?����	�������(�I���[� W'�x��|�j*3�i�\�xq�1���F.B P��|%/2d[`M�����Z ��w��?`�~H��0걺��y�h���ܪ7�]2P�΋��jS�5T^%���egV�����D�4�;�H���.�2�.�@�t&]�Y�_I��d������,}~�ѭ��	A�"5F���7��*M�A�p�ٔ(��5�	ء��+I|�^(��>��{��Z!��Lnو�:w���3�|kc��>-��-��<�z+�=�}���K�n귇��C)���<�1dnL�/�+�,�C�\�V ѽS�+Ѩ<�㢸�G����g/�c�q��e���c��3�ıe���d�ٽ���.�Q�E`�:�9����)T��N�Jգ�nO\�D����t0��~�k��|�\��Gc?�B��ל��'��^;��G)�ϦR	^�N^:�"����9A&�e���<���&�ցV;�V�?�S��G�{)Ϋ�Rm���3�7�~al��A��rH�#�T�O�APŮ�i�Ƀ���r�e�R �y��{�JV@[������.�ii���P�SɦT+��5 _���)m��}W��E��:2�x�,c��v�,=
� ,�Z�4��<R�t��0ݢ-��ɧ��P��@:��t��>> �}�&��Q�Sdŀ��չ��w�,�#&��$�mm!~���ft�Ls����� ��c!�)���2s\:��
����-J��.pz˥K�*!���|�!�ۇ�>8v�m ����qW��(��`�i�ӣǃ�3���P�-�
�W�['�D����D����cR��F�Y����}7t��!���W[o��Q�t��
�$�§Mg4�SYl��G��g<�Q~�a-�'O�k;�U��Wːl��F0�� ,Cp�pn�퓘o�b���i=����F��>�c9B�e��R}�L4�Ii/�&�)M�1H�$D͆�8�wc�����tf�:�Z$4�`mq�A}`�����H��o���Q��`h�B\4�[�F�^�4��[�q`o�����^�Zܔ���E���f�����j8 -��nG^O����m��U�ۆ�^v��!�O�/g�IM���)eh~�6��U�jet�i���#��m~�Z�t/������[���R��W�s�3��'��3���-�tI4'}O���_�é�wT���,".�+M�_��8���}��<>_�z�����Z.��0��B2W��G����".i����QU���Ô��:rhq�� Pm*<G�$0P[iwc*%��DL����Z����hK̢A�'��F3z��LN��\�O��r����m�|u���.*��������������Ƅ����Ƕ�ۏ�}|KǓ2��z���Ϩ�ua*"Ƈ0����j�U*��1ld��k@i��~���~�~��<�b���D�4�)-��/}��D�f	�DH����RA�6I$y�#���a�1�k�I�ig\���̻4X5IOc��bnc������?S�P������ߟ+���|�IaO8�)*����n����R�j�*i�7v���.���ML�F����޷��Y*ؙhG�D\ض�1����/K�K��fq"�@&#���6E��,�V'����_��
��E^�*���SQ��)Yb��<F�0��R���R(�34V߃�W�>#"��&�,P��6u9
\�96$��u-��"A]�'�Z�F�a�XZ��s���Mf��eb5C�����勊M��$���~��y]F�pC`�����\/���f�\Q�����˴��r�cS�F�����\�J8��HȊa\�z�ݱz ؗKߣOН�rN�qC�r�qDo�����q��B�Ȇ2g��}b��ަ"�o���{�A��B?�#l	�������0�u�Xh/��;'�u�?K�1���<�����e����m��B�}��iz�M��B&�:Y�
�xI(Ջ�&A�#� =q�F{]���2GC����N"b�/n�*�͵0�����I��g*��C��
�~r����ޡ��8����>�z1�l,PlG� (:�U%
kY��b�6\��a�bqD
�]�W��� Y^�>�?�%86�I�������I X�n)��+Y����)�Sv�m����Q/��j����W�]�ť/C���U�Ol�����
��K�qf4���ZEX#�p�>��R	ACyF��E��uz�����!�$���)�kA���bQy�1�� �9X��GxK.�:���ٞ��=HE�BY%C���f�b�n�=�v`"#����?>�
=m���{J�����0	b�H#h������*�?THVv�����w��u�Q=��sV4<kk�k����<���J�A��GTb8�������_��,�0J@��k���6�2<!���D�^h��5=�2���fX[b��\M�;��n�����e���e�Q.�zJ��.���V���l�s�1��|>J�i n��v�m^�\����wbuo�[0	�2M��^"5�,���^�РbdA��ts�۵YYi�$6[�>�����_(%J֕6�a�&�*܄�f�?H)��A4m6>%��_v_����k��ͩ�ͼ�Г��E��^��b���f����ɞO~�5o`�K���8A|�@�=�Zl��<e^�)~�_��4��㌬7�(7Re�ҹb*=׺��ww"��sW��MR���f���G�D��(t���(���O��_�Z��Q�h����:Էn��1�]��! r�(N�Ļ��L�n�5��&w�9'����ߩ�1�����#��S���z摧���-'M�٬�̧���ȅ/�G@�Q�"�~;pl"���hG�{Ա_B����ϴ���3i:��ӈ(��J�����`�J�znk�,�JF󌬓���R�*3c"���q�)��U���VOdU�$�,3)Lk��4��g���u���k,���in�݃�}�2֗e�E��.���׹aiLvGV�)�V��r���2;������ǃ�����F�/�9�)���k�&ǒ8�u��β�=��$a��M�ٞ�Pg��@��Fxw']��K��i��6�~�ʼ$��j�>��LEHA�DH2ȧz%�[3�T�j�P�V*<	��ˠL���8r�����<�U�R��HQ!Hq���r��@��|��5�L�"�	E�e:�>��"���+�P��eWػՒ;��`v�^W'�9+^�q�f�hч�g
��j�������I��Q��`E���h@��U^[(�PJ�iC�R�Uk���ѥ�_T�J�D/O�	?���\7�̠h���ܖ
���=1���ɝ�濝�l~�A�2:@��|�La��� <��H{�I��u���K�$�ɶ���=�a_Đ���Ɏm�ts(�lA���
_j�z��u��b���()5ND��^��E����a�5���{f*=`+��-���$a�:�(��P�/��j�p	2vtp��x���zg& �Kqb��v��2R�F�1N<֯zc��;PI�,ˌަ[5{�/n1��C����6��p���L�{^��mސm}x�x�A��f���Z�ˌ�; ���~�%$��1ID2�N���/�h��2��p�y �6�N��&R�*�#���u��JQ���[�|�3��e,���u[�OpT"�g� ��]��$�����H@B���\��%lG��]μ�ȿ�&ZCo2�qs���>����x���J�b�Ҍ�g�S86x4�S�:H�A����j��{��n�Uԛޫ������g��5�.R^`���W/�H{�ȣ�1� �|���xt�e|���ș�
���dg*)�g�-�k��<b�s��~�Z���\��{��rj4�)��'cI;���!B���z���o�oj@��c?�Źǯ�r���.��08Vő��oz�&���j�x�p�+q�,1Er���bX�j������,ƍ��&( ����b�"�u����+1��y��w�+���vj|�������L`�OS����YH����9��z��|�{�(��3������߈W0�����R�������H�S0����vZت��)�/�I��,���l�K3tg�5�G�\'1&�J/�^x�?
}����ҷْFU��J�RZc �7KAp��}M*A�Yq�$[�=.�7��zŲ}�zk��'����3�A!0�փd��"k�K�,C�;V@�z]�hՎ�X^�S�8k�Fa7l�OyĐ���B'�5*��jI����/�h�����!����3+�s0o)8�|:d�(�]%�Gn���~ve�[��?5�Y��[�6R�����ǑtϟO󪠗)y�4�H��d#�JW�,-n���jP�ɘ�"O����Y5��V�����nG�Py�D�����]y�.0��p(��ėÞa�<�ū~EW�l)k�X|�k�W�E(�a�c>�W:a�*���y�݂��~��/� n<��]��[;*W�p.
u ݽXǬ��Xd��Ӿʍ��R�U�
㭟[m��KRx�dZ��+'��x1��C� ����ƙ�Z�ʅئ�=�ۊQ.�	�k墼6g��i���5�~��˖��߆���,V��71=�>�7$�A%��E�`ȃ���*��;���دTA�Q�5���c��/�+B���k��s�����ew5,=��"�KMp����LEʁ&QJ�§�ø���c�-��mfx
��p���tְ;�u��K��e���3T� 
�{
���h�$���	�p�8�I6ﻓ���[��_W�1^\�ė�iG�%d���ƹxpV�vH�$�˯N��#윜���O��e����M����i+]�;:����Ѫ�ӳ�l��u��(�q�z���4�.�~������f!-��{�⍭h�^c�[Ʋ����$01��6gJ�
4������-���.�b0���D�rW��asQ�Ǭ�*?�ԯ�	@R׍a.=�π�f�͸��%KE8^L޵?� [����I_�A�b�|��5�B�i�N���
b��b�5�X]m<��i��ߎ���O���ѝ�ۙ���S��J�ba��G4��"p��K��j��"�jk����e�`
[Zmk9<���	
bF�B����%!�U�@�Y2Q�����g��xx��%�r�^ӻ�2���]B���ɤ�Hf�?����pk�qg=
�a����!1gmI�.�`�:�7o����b�1ē�pq�*t���1Z;[��"��Z^U?:7�N|�+F��!�����*xgݛ�Y��Uɢ69E����D����P���BI~��b�R�c�B�����Ω�'��T�2'k+Ď���Ěl����+*�F�_3�MW(���a�D��DsQƜ�����o8c�7@g�-Hܘ�T�e��j�Ѕt����g՚�Z{�Hk�q�� �2|����Z��n.2�k�@͉1���U�ض�a��+g��,���:!ʽ./���{GIuP��;�|ޣ��;��^d|L���f�P�u�v�ړ�^ݑ�b��>7�j�����vC?��8���6�y�;<����|^�}tz��E�&����w�-�~3�`RtAe�V���zu�[��;�ӿG� rVpk8]C$�f¬*���K�5���!k�!�_��Pp�UKڎg�S+�VPUg~B���z�_�1`V�Ɣx��zE�!m��$��`��4��I��^�	ѻ�t�w��f1��YLp�m��)�k�Hi�]����6��IYZ�����������z�o���ŵn��=�q��z�.�c-8Wd�U�ˡ3w�h�?�������g���]<2�?.�wj\�ǦK3�<�D(�Z�vU#���`������o��`n02�K%ɡd5m�Q��/Y�N�}X��J����2�����rb�Α�p�=j,b��I�H�bt� ��佛?dѮ�=N��b�*<'�_�@��3'�3O��j��@g�� MG��Oh�U7��_�Ũ+.����Q}g�[��S�' �ׂ8π��
W��U,r�(�͝����M�����2k'{/x������֓�!��'���3�Z)�V/QRƯd$�Y�N��v���>��}(B;y��2p�P~�e_��GlTu�(z!ʹe���/��L]Z��=�0�|�7`(��& �}x~�;�ho3�h9"��{J�uZ����J�x�^|��I�F//��z����8�BC	7*�Uk��߀�������eL�{X�"�@[S��R�j�K����J�۪�Ő����|i�;Qy�#2��!��X̡�iF��� q5L~���NL�D�Oߐ�XE��M&���1�h3
��$HvE�,i�"˟��g�j��+��~%�ZXҀ9�P*���鋆��SU�JS@�����������%�-��H����^5��h1�ѽ�['$��\��i������`�ةۧ�Z�Wt<�	�k�s��r��ž��	/������m�r�p���v�8��iU��t�Q���Eʵ6�*L��9�o��v�ր��`1=~���\����m�|�K�SڗT��}�h�(��֫o���Z�i���:�����
T��|6	������d��^�҂R����&�>r!�@ �C�Y�>���i���em� ��V0��~����ZC.V
���<�E�Ϭ"���e�Z�������޵n��8S�c��3խ���u�Dyn��D�&����&��sn[�%6�����6�/��|�n�n踴�W��X((x�����<3X=5Y7^7V��[<����_��G�:��X�����uW�=��g��
�>����0e�#R?v<�0�{Vgf{X��u�����z��$J1ӔH��Q�R��3�#\��R�S߹�Z:��<����84�F!=F\�VM5s���cPg�'�A�k��#��W����UZ��~������%�c�27d����C��0��?7�~���>����B]�B�@ ���<r�]��sI�`�Q�W���^�+�y��90E@��n��]�����Ϫ�i�K`q������ �i)��c
�2=����%��E�j����_� 8�xx>~�}�K�-1�<s��B�^�FAOy�X������rD�� @�u޶��;�|8��Я ڠ}(�����~�Z%׾�Tȫ$՝��Ei t�V�lZMp�Wb k����Bu�)k����y����B��X _c7��-��V�OzfI��~��V-��9�9p�4�{�*���=q�d�������	u������%�]�<Bz�	��9��/��_Ȯ���7��.�ҙ�Z�T~"��Q��)y!����&��d���g^�Β*Q����Kd�%�:5��t@$2a++<U�J5@��m����Wa�v�.���Wfz�Vx����ӥ�O����7��h>��/%���&�qgsJ��{��b�)�=����9�	W��v˴�*��X��9Bd���z�?���Q�����3��vY&�G���[�b��@ۻ���R�._�v��dVV��nKc�
Na@"�:��v���F�_�������t)�ԙ.���L8A�� �uO�P��BٙN��EL�&U���y�z���we�T8Q�������������Ç��r��񯎧�J�Z�bF��|c�P��ǌ\)�X.3{��#U��>���S�A�'�=���$�<t����N�KSj<�?��2)��_�rG:��U�5�šO!&�{T�Y��8ݍ�5Fda}o����WQ�����{/ӧ�0j?-�ޗ+O9�D�CA OD�2҂�'|�Ҭ&�~g^����W���[Q\h��%��Z���>��Im�;��"��t�j};9�;�2
��&L	"!��ٝ�I�'n�@�9t�;̊v����IĴ�&<c�OM�ᱠȜ+�����a�K�2�P���2&]_.M�G�[��bc��H_�lj��X`��/�r�6�l�r"�x�n����}����Kc�t��^���F�0	���[r�Jq�K�Ԗ�W�7�{��^�To��h��E�	Z�R�"��	\�i�s�E�2��=�����������\��&x��(��<{�/H8�m���X�r���̬����(�P��+����&jxίcuI�2H`Zw|EKG����ū�<C�q$�A��J5�.��`�����9.�۶�U�)�~^5ϱ89SV�;YC��9ǯ
�r��}/�Ȯ�l�釛�n3N3w<	K�c�z8e�(S�Lukg/4��ۆ� �\���P�J�*���Z)�Ӡ�+��C����y��d�-T��m��®@�8y����/(�-ܽ�A����8@ �~����h���H���ؖ��Uq�����wQ>�Y��<�xC� �.�ZZ�(��j����  ƙ�[�2xF��Q��z�� &�$��]�iŁ�����5B��w&'�z;�nE��YhF�&��V1�ˢ�g;+	���A���5&G�%'����� l�w'0����B�s�uJo�tX�Y����0���L��Ԋ�Nx��S��a���|�ћ���)�]��!��r�˩�"�~��m2܄��Y�'^q, 8����,3�RU�`ሐ�����YoP�:EL-��h�R�Ϥ�ȇAT{�` �;4[���W"��@B����5���U^��4}>d�H
�+�����TS�JcA`�?�I:�_8�̀��ӤZX�H�Ż'L��M��I���/�(���<����^j��[%nZtKMgsrT�xZz9xA�� �����)iC����i)?��e���f]=*K3¢D'���O�G�sU�c���|�CL�fwU�
�g�C�Yn�n�f+qF�?��;����uI��~��#��g��TJ��P^Х5���qX_.xW��݄M��2�����/��o�x�Z�v���Y���k�!������y"�dhYn�/��u�T>�8�9�Rr޹�1��x��{ $u⌴��.f�V�;��M��}�S��|�:������� �������m�qŘ�Y@�^�{2.� Z��jS*����9��`�<&`R�I\��e� G�1�lx��@r�+f�Q�Cq��Q�37��CU� ���9$4!�ܻ���qTL�w@V\v�O9k*,=s�q�ў�"m5k(�����|V��{��
.k��+��g���%���弳o�I�������Ȓ�o+y��`!�Nx��R�BQ��(�Y��)?a��-�9�s���!�'E�n7������eu�?���[濭5:�/��F:��8�	�hѐ)7����\�fjSk��(�<�ޡW����*1�����~��0��0k��:�O�kmBί�XÃUH7�К�`\>u$�JH��R3uu��"�$�ɎC&`�F��k�ll��C�
U��C���uc$t�X�����]䘾�݆0��mU�G��[��UQ�~Hf�?2��*�`�8��ڀ$����Ʋa�E�up:/�+{�a��
Hy�A��R��3]J��bG=b.�Z�ߍf&�D���TerP ����^kN�
H��Â�ݳ����Lt�X�2:�4�V�e�8��,3�Ǩ��@MEJ��\�T���u�a� Ql7��Qp��Y׋�B8�V�-�M�?n�4(LG��a|�I����6Fu߈���U�����2��n�)���	cV�x`g �)xy�Y���:�ױ�z���X}�*T�NkٞIWq6�V|8�x���xb�n�,g����&��ob��X�=�Nk���|���c��@��ǐ��z���ʗ�h�q���TȻ���ђ���"�|���į��(��m�>;<��&����j�]75 �E%��hY3u�Epw�>1�kD8�m�c�Nv�&�;�|dZ���퓱0X�̵�:���|
���~2���[R����2��2�"�@p�-�����K�v�N����C|����ESy�l4���a��Sn.1�>�CB��ʓp�^R���c�m$�L���Vz��ڷva��}(���d��h��t6Ax��Ub�R�G�` �h�tT���-b��ϐy*�?�.�@<�C�U�Z��c���n:4��탩WTs>��B���΢Rx����Sw)�z���hUa!�'��'H	cx*�*=�y@�/��&���i	ta�G����k�3����5A����Ǖ�2! �o&�S__�A�8l��~�	�`�f$���i݃��E^H���]��}���&�w���L�շN���#L�i3��4���?��P�?��[i��_��Ʀ�^8fBY]M��E[��~P!�,�x�5�Q�|���G���	���R�*^�x����6I�j��~U5 N!S���õTn��H�8���N?mAxO/-S���l��Eg��wd��:���%c��!d2��R��ΞK-����ṋצ�G�${ݷ��9�Aj�lS��6_��u�q|j�N��H�����'~�R*���G��e�O��O�5���V6��ʪ�Ө��ܶ�{<������3Jꩳ�^�6O0�p��9s�'��X�����d�(!�l�N͜i���鐧�D��!"���R&{4Ga�r$��X-]{T��1q��>3��\�Z萖�W��$���N�U��d�Pn����������OVؼ�ZH�m���o�%S(�6�|)�����yd����N9�U��|�$���ѡ���X�}���]�g7i��[%V�,8[����׋����TY�`[|����Na^��|�R3��]��j
�m�Eۭ�i�g�@�\+)��7;�Ni-�����[~�B�$��E��R�G���U�!q��#�嫙;C�Ti�&R��v�Qp��_�!r#���<����-�`���0��ЛK�r͖�NN����剡K/4
��J ���7M��8;����Y��B���#~�-WT�B�S��G-����"	�* :u���e�
��W�$��=s���J��;�u$z���' �蹢Xx�'�ob~�%���j4�àI���eRA6�����L̊�J��~B�B��R���@�	�d�	����B)�W[�|R����n��z |�#��3jȄAk�
MP���������2�"��Y�M��sJFD��AƁE�������cr1W�O�Wߍ2����xh�Ԕ���\n��.0�E��d!N�|k�P�j%ԭ��_36qY�c�LO��S��b����7�j<�}U�7�1��U����c_��_] :A��ˡ�%�qK�?��º3�EP1�wh�������D�V���5POh����6a�U,�;F?����F������DyWc����Ѫ�z��R�����HUI������6������0b��
�#����&�y�mR��p0��e��g���+����/��$�O���Ƅ�/���5���)3)Y9�&�m�k(*_���r@s�P��t>u`]-c�-\��\O�%���,�[�6':�W���P�Uӿ���o5�M ��o��d��]}�C�w,2%�Fe����Q��ky�"GmS�v�*�X:��^8V�Be|���)�P}6������̔����yX�����N�[BVac���wZ-\74�+{뢈c�z�-��;τ=hD��k�J2�(�P�X'Y����g�=�g)��3���1��Д���h�D��.ru����RW�R��D�%hw0uf���/Dٛ��{��l-�M��x�}璍����J�8d5�\����S���� �1����ޠ�դ�ao���TBr�0[O��`"���h���U�(NܓK�������$�����zM�R�:�pR^1�Tǡ�GH��~i������>2�Q��eGC̺��͍g9��}��&��R����HC�0(bA��+5�߆���9h����t�؂�*6���3r"vI�O�Y瞳���)	9i��/�%���ԁϴ-l"��KJE�bPvŠ,�Y��,H�{i�{�;J"�^���9m���Hp�\k����#�v |�v��0���j���Sw2hũ�La��/ �E ��B��}p	��	n�Q��d���c&���Ծ��|�y?3�����#bS�@e��z
{�`K�e�w��<F���e�Pް4aB�ʍ��1�Q�{�KՉ�u$��Ss�㺇U�GV*|p�� �L�:��"�Q�?�8��!D����ʶ��&l��{ �o �Jp��w�rvvcZу�~�ӱ�-`�9�u|�94���[b��<�eg�L-�;�D�"⾠"����X�x�#�����;g3)�{��y	���r��f
e��e� �B������3m�h��Fn8�ؓ�0����̇t�q�n��~�
��84�W�|��j���8-�m�3�~�j�$X�����1tqϳi]?WV����DM*��X��Q���}����7
�t]��^�{s��Y��[]�J��8���E�Q����Tt��H0IL������/�0�su�_��J~В�_}�o�,G�J�]�򆢸��'!/���4�aN'FJ��+�3<��<ϧM~������xPFn0�.�@0W�i�T&������Q�o���o��XB�$H�D�a����8ŕq+j��PC����7l�d�G@�T9p�l�{![$��������7�����(4�����ef��oI2s>�9�uǨ�-6*�\��H����
E,�/�\q���,�Q����
��:8e1�1ߚ�q��~���Av�<�'����T5�p�y'(hP�^������}�z�f�����řx��E3�NI�`����J	��p]:Բ*ه�=�ai�M������?_z�Z�BP�R�z9zo�E��!��%,M���r��A&2�$�2wN���T�J�˷�� �3��N��^�<x�j@�������诨P��b�Mbo
Z�x�[�`��f�B��ބ�G8=�s��?"u��+h�VJΞ��E��d�#��a��ٴo�,�.]�ġ�R�/X�����<�$ֆf�����Z�'���Bu��,� �����1��E/<f�:Nl`Xc���ͳn��C��$�9vnˍ=�	aZw��� ��-�AGu���N6o�*�������p�퉀l��An�����p�<��1�?�R����?��ͬ@Bp��
��N����8m���^Ċ%&D1��%��~��_���>3JѨp8��ŗv��?���,M����ҋ�r��� ����
��7��Bb�Y�h�m�R��c
ϓ��Y�G�R�Gb�,��H���jqw��Z�g﻾��Ez����9n���
N�C�%��IN1.��պ�����`�2�f�������d��#	���=�mcu��-gz����g�ب��9,O���`�}Q�\b��7��jϹGlCc`��;�Z�.��^tfG? <䄃�&n4D�wTН��EàB|�u �҂58W����/;���qs7�Ra�E���ost �1��@��e�NQ�%�H���5����^
/�=��󯍢��B4mE��T��v㚕�v�����"��	��������NER&�T����P��-��O�1�o�׷�G���2����3�\:Ҍ�S�3	����H�T�M%����<]3�b�wf�.�i!��pӑ����H�Ȥ'����+Jo�H��UN	;�d�����&� >S3sb�̃Pw4��O$�(�`o� cW������=c1e�RƎ=���*���h�~m�B�QrQQG���҉���q,�ebܣ1��*�*��~6]��8����s��>�%�m�գ��ۏ��PxR����#�N���f({���ݱ��Vp�(�	jqz�a���@Hns�I�Py����Ab7��߿*`�z���V�IC��[1�ܵg�i��ن��]�_+p�Ȭ��Ս#6=��S�̉�C=+ڢ�2����Â�2�?�JÐTbR�����jW���]�$7��D;�����qε�pM����C�ČR����T�Z(��?ؤC����$�\�3�*�F�y��7��lC?���r%��^ن�o����&�Eo+��[��"�6*1�KG�1�wS$�u�P>y0Ȫ��׾O���Du����Rm����m����ȧqZ�CbL�-�&���U2�V*Xg]~��XRj�K�~�{�}˜�u��[�)�B�"�����vy爒��ςB��4"����0����ObG�uQQ��iԤ�h��V � ����c�zMW'��q YXj�X����"�k�����NT�mpkNK�v cX�WJ��i��T�at�g�"T�A��,Ԡ�"o�N��z�1q-ė��S��$�(��7�ZonI���%{���$FQ��;,8��t1y�F07G��uN�Q�dL���-�Nf���wa�ߙ��M���)J���T��������"Po%E�E���!�bǯ�_8�GП�*Y-cU�a��_��Vdg�䇲�$mVǿ�<�}�dح�3�|�J��*7UE�j%	�V�R���[%��C�(�����ڳTfIgG�4�ɹ�8ʖ�S�Sׄ�in��*����6ɉ�>a]�<�B��� �}L�=�ٚ�J|E�Xx�U�?t�{v��'}�2�� �x}��U�6�az�f=�S���V<�.�h�o�܊+ACg����0#v'�4�娕/�<�J��B�Vp��Y��˭:��?]��#����2V7e%wz��1�"��O�ȼ���U�־مcg]�(j&3�Y1�R����7���I�`T�J�=��&�D<vM"�i��
�|e%b��['��J�wț�q���f��d�8"I�؝�ʕ��� �9�qJ���0�8(�L�t� !�`���X�{���Xc�Uk%�5�_�v�g�օ�ٍ�s1��~�w��GǪ) �O�q���o�!�ϨD��yP�2(�ی^���wW���'�@-��E�6�)���|�y�L^�}�h��e��J�.�DOZS���ɍ�ߥ`0$3�����n$����^�.�]2�4!���yڶ9��V��M2����
�(�����	[��?γܩi�Kĸ���y;���d� �av�}z^P|QT&Q"0�,�S�~=�s��~xH�Qot���U���Q'*�-\s�xoG�;�{��܅$FL���x�]i벴ɕY�~Ƹ�%�m2=~3�%16�Ww�{¸�Ci�w�n�;I놅��=�Ɯ}&�U(���L9�ΆD�fnC�n������ ���`P��Z�6i�=dt�������g�q��Y}����m���6Tk$/ʌ�G��W�-��ㄲ�N���)!���$Њ�
�R��ک�YՑ�؝���H?�������(�DNh�@g�%����ҽ�Qz������@�I�� ��h��ʏ�
�#d7�-/��Y����������9�^:��Kp�U��n�}�|���j'�J�:���x2��(5k���R���O !��#�Aӷ)�H��[f ������R�Y�8��5�IBRKg�Vy>���d֧W�'l��J˛�1��@)���B����,���������	��>�V�t�T��݉pʾ�B�ʛ4���q5���-v�U�c��~w��f/�va-R�:���(��8iM<�o�dt�X���	���mH�\��Y�^��K��rb�x��J��Q>�c�'�`f��
^rn��C	?����p �E�T{` �1�MD-w2�]�y���\Q�$�~Z��zُ6
NX��t����/��~�(6e|'�H���jS!�v8�7�a�B�R�AU����/ٳ ����H�a]&N͞��\sM�#��]e�'�b[��'��`bI�L�>W�	�\���zg:�e�ں�>�#� ��5'�������C�z����{b^oz9r���-zڟ���T*��k�C'����v�ٳ����λ�s?��{�>�܏>��ѿ � �Q�vMA	z�f_���qY�c��./�z=��G��T땔��ى	%�`UA2G���+h��R#��DEC,�{��<�:��=��M�����b�9D�U�`F�O�zc�.�qz�7�7���W�KH�������Μ[w͵�v�v����RB�yG7����,PQw凍�>��Q_���q�q���o}+�����f�A�I/ܝx��_��c�)��v�A�D����_E_u��n�,e��x���~5�G\6�>�j��1���6�-��?��&ѯ'��:���-kZ�r���Γ����2E;�j�0��l�������W�+���F��坼σ��1/�")O�`Io�D��j�fG���<*�f@ePRN�����[
��
+WMU@�;���Y������N�poPM4mV�����|uh(��������~��|?��OV��P�A΁��a3��Rg(>���J ?��H�	�S�8]@���^������5�/Of��k��d��1���-���t��q��3���;*�=�Qa��{�~�>^ ���H�G"p������h� q߳�D߼l�j�`��]f���[��Jtn�v�@��j�c��D�)k`BR<�o�ר�6 ���y��k+e�`o�����v�T*�>'�1R�M)hh�ߓ������4�\BR�m�"?�^fF-,���`r�Q�.&�L����c�K�k[2x-s��	݅�8�7��A3�`���#o�]�xø� )�c��IW_ٹ����}P�Z`	e>I��Se9�y�F�����BsQ���iL�E>8Upz�3�g}p�`�+ʂ]�$GX�d��_բJ��H��G��1ng\���q<��������a6瓩N�2�z\�)3��7����mZX��H���{��u���uE���|k�H?j �3�u<�-OLB梄w?l�dMm�| ے����"s���%���n��3�n��� ��,�##2~�<������\Y�U>�e���X8������tEWוߡ���l�;�mX�t��I��������uv\�����F9������'���;Q7�
ȣ	��J�9�j>�YĎ'z�'�,)�����Cᝆ��s"���U��z����	�?����cH5�EF�a85k ���'�,Y��Ω�&�k������IHͨ�>�E�����$!��K�A�k�=����ű�b8q�l����'��]xk��XD�G�ą��/-���L0��%��_Vt	Tz������<���!���t��Cϡ�yk��������5�����t�乶��q��&^
V�tjU*r�P� U�2R�T¡0�#�[�H���J`�%k���k	����3G�oM����<�*W��W�
}72[8��w������|f��M�`ĴvҘh8�j�x,^}Wӹ�=�ڋ)��[�� v�����8�Z)�x<�.kn�V����=&v��N27�S>4|��>Ώ��Pf�ɽ@ �<����Z@����)���Q����	�@��IUi'�L�g,���xuP˚��� �L�fz�8�؍���Fڑ����,���|r7�p�@�VhƣP���fr8�a`���@������.��߈";�C�(�H��{)f+�q���p�Y4z�@6@�*�)-%1�j�n~
mNy2�t���J��Vl�L�|;V7���;F?����%#ێ�	�'���Zz�@���Yl'�l��V��2����%o����ja��WV�0��V欉R��i��Ð�.>8���H̿LӰXuq;��i�r�E�C�f2�C��ƭ����@�1�?��=Ȓz�������O�J��f�y��e�MB��f?h�Q*m���|�#|q�����0�I�Z�}���C�Ab��@lۭ�r,��0s[U�q`0@J&�Ƅ��ĳ�A�����`�Ѯa0$p�����h�hҙ��]]Up��%-��[C��F�|@��N���*7���N��s�i?�xC.�S�W�dB��էj�b��5�E��Cn;~�U�}�U�M�j�}ɲ�Q�PS%��i:��~C��9
�!�rs���%��y4�Q�ҕ���\�~�BT�ʅ,9�&�f�Aw�41Q�m LǶ �.L��W��@q�P�!em�C>��,��[���ndih2�8�)���;��5�J���s�jE ��H�A�j�T+������6r<k^��u�NFE���H�w��9�>�6�ު�"��鯈WU��8n�����1������aLV1I}%x��%�E�UD&i�*ƥ�쇟6�z�-k�xq%�� ؕ�4�R���\�T�eݺ��!ӱ���bp�� U���GM��P�ߞ���0��);��u����q�6�A�#������1�q��%q@{��� _h��).i}�6��i�Ȑ3!U�� �+3����N����<�Sflc�
Pй��t$�$	�wv�E&1[!6�����U*ozA.�-�0���os̈́�2
��4 �TԷhUHM{�JB�B_���!���p��pkp��hW���k�S�38�9�ЇHg�h��1J��K��\�c�6��%�T�_3�32��q�K��&)�����VM&wB|A��<ee�s�y|��ק��m��NnG&�=��Ցl>Q��,�����(4��_�~©�q��J>�Ą�s��mAM� �m�%86#�Ԡ�kn�����H��G�w
��c4�ETi*?>�ˣ����w�Y�� _/=1L���;-���]�=� �-�b��,!栋��=N�f;��s�2J\�8K��r��@8���<b�����Ϩ��cr�.S�%,��a<�����nz��>�ޑ��L	��3XBp4g�x�_�F]�_A�����*�t�=B�������9
>硶ʢ��S/!���G���� �/�n1^�GN�AnR�M=lS���	�Ȭ�c�(���3��y�'!���~��V0?���Pr����s�&D��x�VKŮ�wW�">��D���D(��1�����"I�p�� r��tA47�H_;� �<�ȫT#3��(�h}��i��D�_�١�ݾ��:O��pY8n�w��(��Mx�pS��ٳG?�;����DU�}�a���w��od)���\����,G�!G�:�����Ds`�}gM�'��V��� ���d_�,V�\��e^�TU�ĩר�߂�Inj����#�B�2�RA����f���eZ��l[1M��.��:F�q�~Z���+��+j1�5��F�F�������6���ԧU�'�*P�>v��~�_�o��)�M�oz9��X4���lzVU���vYU *-)�d=e����/&ިh��sFwO#�]@��aqb����
u+ 99�����~�����~s}a���U��#���f�.��K���HA��(ILdٟ�H4iO{T	�0�M�A�Hz�A}ə8���W�v���n��x��Xp��H�t!.��A>�������x���p!w$5��bS�B�>>@ݕ�����nd�	�M¶�h���t�<v���H��z�R��>�i�mՉ��P��T(0z:��I�gQW�^�$Jh	�.�.a��'�xϒ�tW�f�W�
�%�pPO�y�� �mu:�f6n�mI�D�"�L¿�f�V�{)�;9���K:;�A��v�>���`���5��b=��3�wv��g�H{J�P�ӻ��҇COo\Y۹��o;KB�o
�<��`By6�hm�Dۈ[
ubhu�0��g�Sۤ}@�?���5��ׂ�5���;�)$Pwk�s/Ύ���*� �q7?l�:�p?�ϋɿO�v�ܧ�LO�M=s�����PԓWf��s&�2!�~�:�Ӓ'5.�6�Pgs!��*\5I7��*�j�`�U7�!�|)+»��}i&J�]�	3m��!6�x� 7�iB7��>2��٘�3>���3��E% ;iE�ޤ}�U���DJ:��xt]t��jݘ�B�;�1��U;�WV�-'NSV�Ҭ�e�K���oI[�x���Hl&�P�����4��p@���z���˴y�ڗ4Z�DX�iS��7nxe�MI;��s���Ԙ���f���� �H7�� wt�q4�XP#����- 9�m72��M1�wT(�`��=���)�����p_
8��U�����\ء�׹�$��!���6�؄7y;��Ĭo����ҹ$J�_Se܉��[����id'���5��|���
���W�3Bջ;l5וz��B�
bÖ�e\O#�Q�<:�x�`bZʤ"�Z�^dH�k����s�@{�����5�4��m7��7^P�[�}�����K�'{�K0'{�Q�n�7�����c���������$�B|��"�9��܆�;JV�a���'�~�.L��C}�N����q��>��ko9!X�!:�YX���Q�0���B��5�1�H�7����icl�P��İ8�<u2���di�1g�����;7���T9$�޻c����k�=4������f^* 4ƀB��^�(���F���!�\�2B���2o�P�0L�����A�z�����C�a#t��M��n�+o,�e7�w����(��h�F�w�"1�|h�{ulޜ�w���T�Pm��wO��O���X��ی{;x��wK�5���BWQ�`=��Ey\�2����MR�����F�.EQ3C��]���Qg��=>A�wq��1�$�,t���st� ��^�j��!b��z��]�R2�y@7�!>���q�0�Z�{����Q@f��l18��~6�2�-�����6P���%�9џk�|�%�:�~Q�
S������f0�=�x}�O'��3����F��A��B�~ۯ싘^��]��ib��8�Qk�"z�~H4�˷"��ܙ���0���ZR����>Zj�xFv1�}�����c��s%~����cK�~=&2�0��g��xI6�*4������b����=���XUx!�U�>W\�u3W�cr�D�0ʣA�|�����v���%�����s��-�
S�W(��.At�#�Q��l���(��腛����:����:חx�B���1т	[~d,e[���(��ϊ�?�w}6A��&�ǳ�����\�{;�Lz��ҫ'�Y��d{"�e�r� ��P�f��o�/;-7#����� �B���{�V|�T�v00�w��d.Xxiq@d��:G��DD�r�u9ήn���
����Z%L���D�g32��9�VHQl� �	�aV�5�)���7۰���caz�d�i����5�$g�}P`ÒV$�RXW�e�}��S�~��̾�[��,��_|��F��^Z��TYP��O���x�N���]�����Ͼ.�����Ɛ�_�Pv�=N�m�	)��?�V<4���j�[G�ɻ�R]���G�{��E��)Z�ڈ�J9������7
��[�~f�${?�x_}�GH�>�l�2�gm֌/�laoZ{�}�����Axl��{ä�t��"}��3i���P��س6�E�&�U±�<��[֡ਸ���t�*ͳ	�z5.]���ɲ��� ��NJh�$代����b���I��`[���(�=�'GB��Ef��B�H��_1���͎�"ԏ=O�Z�D��SGߪ��wQb7q����1a`��P��c�\�4il�/�՝D�|c�� %�(����ךS�;�yh/ai�x�ŵIs6��5\a�Sx D�
T�`��ޚ'��gA��/g�U�u��Y�6?فO�ԑ�}
ڮ���o�����Z����2�?m+H��vt��z�+�����E[���~_���6.�P)�|��^�x�F���ю��&�r�V 8;�ؒ�aj�@Aܦ���P�: ���8)��Ě�J}��}Z��!���>cb�qW�썆vlG�ڡ����Y&=�v�I�_��A�ѵ�V
�����h�n%������@�-��WU{��k���0!�f	�.�璅���I�R#�	��#S���kos�7���`�AL�߽�4\�3�Rð]�g�P���GP0)���L[���f�I|�}n[�3�jk8@����YC"MQ��s���d^���o8⾬�N�J���� *0U;�0��� ��j���Ԉ���LԦ���)v��mY�C�`�0�����@��X3g��f<�s���x��G�!ňZo�]���)	>&��@�@0�>�z���d�%R�3�zg�ufr��:S��VBUo])�rC���Q5�X�(P�R���P{��/��z� �0��_RJ�����'�����u*�ת������"ք������ � �YT����)�ݔ�Щ��ݧh��
�X��j�+�P�O�f�S	3���`�o��<�"�\����&]a �aT�`�ֶ`Y��~Ѭ��\ʔD�G��� �W��Y��2�#Y����@(�D/����S�.��~�k=R���#2�$A��e[D��^}m4��ߩ��휲�嘛�[�{A��_�5c.�ֶ�;3��3��w)�Q j�$E��#�jy�5�xj��=��c2b*S���f;nէH�dLU�� H�(	B\�������@D|�k�Y�d����{Aj.��h"B¹�zy�\�vvO���S��q@��aR,O	Cct�D<�0P���S	P�2�q�{�*)<9��D4�c��y���^_=�j�O|�f��9�B�g7	R�7/Q�V�T�eQTWw�7��98y�?k)�z��4je��;>�k��N%�2���3��8�q+��_O�Ce��Z����R���v�y����G�؈�Op!B+��%�춈R!�W����/�e��������m?����_�mq�������ܤ�Hr�!3�_H�����!\����9��Q���P�i����񊋗I�`�P��Z`c�G,o�H�e��6x$�Z�%76r�Az���-{��6�`����D~�DL�7����R�	�q~��e*$�bHR��l�M��,7���1!����WP�?&4�i�>S*ۘR�8���X,�G��Ӧ�8�bl�$�&��H���"��CS^��rAS�����_w�{���̴��i�c�^�٬0V� fUo�k�֎,���5����~}F��q'���YT`����Υ�'�P���Q8*PoQ�ɾ}(H���Ӎ�D6V#�b�ڐw�����
~�����1�ܗ������5�gӔs-�.�O�K��Ӫk��� ��E���M@cٛ{�?7		:�C0a�������Z3��PӴ#	��E\�TE��a�V�[��t"1���!�d�΅��ȸ�Φ]-C�ru�W���a��lG���q&���jM��J-��Ԑ|�8�<
��d�VC�a�M+�����xש��OІ�P��g�c��� f7I��Bv�����c�K����{9��+����4���z\�v~��\N<�+�?2^������Rq�n�~:g�Ue��c�֑�e��m7ģC�9�9x>���Z�k���fYy���a��*4-�4�?��M�)�l"3뫫K����?�A��+E%|�?����է���/as�y������t��)��˹ɉ��'���{X����M_�sI����\�[�OO�:g��������F��%L/�"QZ"�ެ�'�c[��ܔzWu���74��w.����9M���ӱI��hO����y#ie�ݤCM��HT��<[`�*o�޸j6�-y�NL"�Ї���v�*؞X'��Ү9qo�ʛX����u�p�/�}�VS(�9��gn�(D8�����K��.`�f��13���G 
�e�Gv���h�3�r��y8�p�ۿ�o��q��EX*�m�(}>�jC�e������n�O��~z��DH�z�l��оT����-[Pm%�7:9e�3'd��Ԍ��x� ���,ؒ�E��G(�H»p�i�ʍ��u洴6Ol���Ol����|����IN��͟�yMb�B���Ē˩.{�g��M.-��S�� `+t���^U��|��d?�_'[�JT[�R��c�7h��ԩ�w��|�|�!�^6P�@N���ϟ���K�W ���X>�%� '#r����`l$-5�^y4�-�iWSi�"�W����6gkb�bS������]].�e�q�10���Ә��4�4���!��M���
z�
7X8o�x٩�n�й��/m֡9G�ix��,O�Lȼ�;�z��jw�\������I��,+��B���p�v�Zfn�b,�#��e�|B�k�����M��6r��ܟ���NԻa�Q(&�ge�| \Y�u����Zl��2�5�E2I���3���,�W���v��9���#7��)�Bb���Je����o'���|ު���ZBn!�1����7�g���RK�M��a�`�T���V�wM���ηÙ�p�ds����)���Y&a�� %�*�1�����\���_|txlR���J?f	� ��Y:�V>���"%@��E�_�����	F`J.8�DKp���*�!(�"B�K%�h�GJ��DQ9�(�j=n�Թ���6Q,�\� �H�;W#�dt��?XU�8��ȶ���<m�I.'D���{G�꙰|/FEvd ��S#��/�FA�3_����4�oQ�^��VS�>�s.NIq��8Xٍ#Hqg���
��y��r�� �"N��O<b�7�S&C���֕��`��;�xl�#���`�&%(�Ix�7ֹK��þ�P�XLj�vV ]��LJ.�7���9������2�
�\���y�;h��!΄�j�����+"FU�.��f[��`��֫	g(p��o[^w�_�y`�hV!��V4�V��w -9Ѭ�}$�2��z�X��/%������Z[%��k������dq���t�	p �D�3O���Vj�4)���H5/��NV^��F�h�h��o�<wF�aF��|�����J̌NKgaR����Q����o'f+�I�Dda-ۭ�b-��_�}�J�m���,Q�׀kH�Y�Tj,z�K'O6��G�mPs��Qɺ��� �k����M!l� ��u�T���T[D�-�*;_W,��	26�����"]���~��=_R9��1�=�poC�+���rtaj��O�~�g��8B���(>HZ�Q`�l6`�q�wܬjJ���5��y�"�У)f_m�SR��!��;r������;!��"ev25$W�\8�����'u�e�?z�7��!��Y�0W*}6ࣀ���(t�z$LH �,M�2*�֬�ucҸ���4�ba|P<�q�m�-��� �ABE��di�<�:�U�mQSv{�΋�S��(T�������]�%��wV<p/tBqf#>q�>U��w�� a�_%�V!���į<��n�a &�O�^�)�Jm`b���>��� ���;���p�$YZ1��s��r�ᤔy��~ǭ�'����\9��TN[�#{�dc�/��+�v����Z{�2��2���7�i�;�]rJ&���O�L�U�5�C���qv��"��{3�v����k��lv�+]rX�sY�o�;{�A�2\�Vߕ���8e��Kc�+i:��¹<�������{3p�;����B��Ԉ���r�d#QX_�ޥ]�-�X� w5n�%6�a�4
�6�C�6�#ܟ�N�_��J�MR��� �t��k�蛔5w��Qz��?J�j�Bo^cRrR��%i�L�`/E�t����[�닚���
&���*'�Jf}�%
�ec�0�z�r[E؃9�y�z���'萜A�+H[B�g-�x{
ȱ���������{��*MN�6;��H������h��UL��o|u��Ѭ��^�᳴����QՈw5��p�@t�w;Y���=�s����D�S�l�����76�S<�t|��Hmb.8�{9�Ld%��x� �8b	��-4[����!<E����鱮 #f��2P�qX�  rM�P@�|;_@a��C�
���DG;�n
=��6����Џ08����c�NgWΫ��� gI��n���׋�j >�0�e�K���#�w] fJU7�|A�_�K�=/�#�Y9$�����	)�b4n�v�%I1<pKn�-ˡUv`9�+cUAoñA�:'D6@�I���]i��ȷY�!������
��G DR�r�(n�����O�˩��y�,�OZl��}@E�m�78���K�S���-�6�������τ���"SiA꾊?�ӮwA�ZX��K
���b�i�CГ�*Z랰oz���Q/Ż�C�b8I2��s�3���4�I��+�*jԿu�� � W��z%�4nh˔:���"��@1�G����z�`�|Hc/jGQ��^{p��$�{k��}�V��hњ{���a�R"�鈋�;䭍mq��ўR����ي;r��<�Cے|�+}�� �GjC"�mv�_�\ʃ�P@E�m�g���P�<	�~�~�̭`���u;�fSJ0'dM������!���4
��[H��Fu�T˻�_R�TV��#k��2����jp��!��D��� v���0�F&F�'5��64ѳv���z�	��3�gh�o��:V�%q��@�9]ksVe1��
Q��>L��hÒ`$/$��<�����4�S����`����ȩ�A OL���Dmm'G���n�U(�'�����2������8�џ�7'"qܒ����2�L�#��TGv���N/jᛑ��Of+1����G��3(L�zXΈ�C9���{i1˗�H�鍲��`
M�������S�iԑ6(�G�Н[!�q�Wb�Щ�������t
~�A��"����֏�fNA�����H쵹���
��F빑­��OèF)��c��s�M�: �?�/���9��\��6C����>a 
�d~��J�^��a� �Q��]_l�~#�1ɨ~�<�Il� ���aY(�x����lF��{���:�ʐE����4�n'�`��/}��!���z5ą��
e�0�5'�r&J�W����8��;t�E<�mj4��w�s�y�07~bo���:���阺67���w�n���p�������Z�K��� ���>)�vK�V�\���ۄ}�[�b�%�v>�*���8�����|u��)���u�&a���\w@qn0��}���uD��c��CO���2�>�T���E��5zˁ����l�A�|,礘�����-�Dq*ZlI�n3D,!��-C��Ǜ0.���Q�3���H-��
 �X��0b-W��u�9,2��5������ݸUǘ^M.����q�s̬�@��E�?ŌzƠ7��F�1�7yZ9�d#	N�G����'ǝHZ��gUE�i��Z���W'�0Q��s����K�%��|h� ����
�H�-F$Q_ʦ+�<I����;��;�Оha���.F��h2�"*�f���u��s/M�f���=�_�����g�YG�\��Ln�!	�2�����p8�)�BV���M�3,55�8�,� {"Z3(>�����������E�*�->L�Dq������a3�r�O9TI�9�I�k0�����������ǋ̽.�w����o����g�7'�V���;+�͈�.φ������%�M�Y
�>ޙ_�ľ�$�,�88E��~�t<��kfbc��s�X��3x*@a���ՊG�8�,����L�q[{:[�wS9.%vk\�����&�Tz�1J=�/�?]�Τ�5��/JȡA�8 �8��YZb�-��U<���
����y�X�쿹����[H q���"�ļ�n�t��՝��� 1yTwh����~�V�G����y0��v[�� &��[dVsΓ%��p�)��"ɋ=[*�>Sw��vmA��uL�o�,k=�GL��*��@W\M j	T�of=t�xx��AE��DY�u�xu�G�iT�k�t:l~���	�%E`=�X���n�K�vX|Ҍ��Hd��{#�G\)-����\ZF���7Iji�C��W�����4.
�U�i+�J�7>�ߎ*�S�i�:N�=��J� ���;�.����WP�n�=S��0�W}��/g `��W��v%����)^��?�3F�u���?�J(qDi|?Nw(O1�ʋo�j�&@m�u���J������V���{y�<a�=�A��i2:V�7M�މΘ�LQ0���u;?�T�S̘O�%|���԰��U^
�;tb�{W�UY�)��v��J\�r� 047�����/1���rW/�U�Z^���n��u�F����H e�31cYv͊}�.'�����n�+��&�ki5p�l����*�| :��捣��zhObڃ�ʻ���_�};2\x��v�8-�Xh�4JC�i���4j�ײ�q�z�Կc�aj�O�&r|����R�4�b�LN��b��� �)���}��I�b�vJ�� ��x���d�[6�¾JdI=P����q�@���.�#]���|0���F�5a�&�J���;f��Ҕ��f�<#�`��g��n������������E{����e6i�Q۲�%��y�0}�*�Q�H�	QI��8S�23�e/G	����g~�$1��R6.��32�UQ�}���X[��<��"�..�ߓ*8��w�����E��3��l�, {7��S��5{6��l����7���Jn�G!�Xܹ����M��-��=L�]��X>uZ\*��s�}��^B�����]��Ds�r0p��U�5�HP>���@o�t+�pG͜�%�Ij�ZY䤢e'Ї*� �w%9��_�p��;uvx��K�X�"/�Q/�V�-g��3���5���*����ӆ�L���0�A�ᛨ�?B7���S�'�� �\e�m��T\���Z�0R����2D���'G�V��ǂs?�z�l^l``�,iH��hx0:q���{u��̭'eڹ'#���8�瘍Mf�B;aȃc�t�c��~�b��&�]�ܛ-�RG�V��̜@� z�%�oyO�����7`��Y�n�Krˡ����z@�z �[��-E��ûv�j�7�f����;�$����A�2ة�'�la���!�|�-�2�= �y�yp���<V�����^	ny�]6.��U@��,< ���$w)鎕�	N�@�p��/�e�n>�n>_O�=���A�<@�Jg�꾻�t�T�xp���.^{�n�i��*<%��o�q^|աh�7��[|;=?Y�g�uH��I�5}��&{�<��Dn
erjǉv��������J�v��Eǹ��G�D�Cǅ��1���<f��vw���b��I70�z������*���"/�4���0�^���}W���ȩ��`Y�O�=����b!fp)�-zˢ�B_Zm*�W-]7Jw��_��R�ѕWz^72Q
J��~b�p���|SZ�{�!��i�ai� ������Vi�Q�D��duj�ϕ���!��-�ws����.�4OkuϏv:FN~�.���Q\��-�t���$Μ;������������o�)�����:D���s��ZYaM�M⩯ P�,�B���>��AH��,�����!}�e߃�.a��<y�H��*of�~^�}`�"�����_&1^�u��
Cs7�]n��Y�{ѽNOU�1���p�ڦL�|ڧ���q��Y�n�qD7�L*3Q�=7t��^����%�e�>�,<^F�d��,�|���eI��ƽp�/�]���c6h�{-��E9�b�+�[������V�a;� ��X�0��z"�Z=�Te�ˑ�����%�ŕUg+'��,��@#�b��k���ڠa` R;"T�.��Zwkg2X]�<�yޕ�\�k�}�<gq?���$A� b �ݩ��{3n'��"pZ�`,�����JD�U	$� �8����DI��¯�0my��R���|���ȵ�vI:Bv �a�^���Kudo]���E,fQ!f�80�Bm�Y!ǯ/1|��Ȣێ��/|;���cj�B�'U}��n�k�z*W�N����X��`�(#���?Q����c���t�ʢ5��B��fX��-��M��@ln��� n+�`l��2�?t�&4 4�e�{�[�Iɣ�p�R�/�Je�hR�;�r��;	������d:��Z4f�,�p�y��ߢ�u7�7�͂��:�`]~��e���iu�G=���*^�WV�{H�J.��J�>d�%Q����ϯ @([~Z��N��I�G�/��OI�Kj���T.�xm=�;���`����c咊�E�W5!U�16&|�tl���zkWbcmTj>n|���O͸��.P�i�c�ʼV��ˡ�5�:\����|�Ȗ�P�<��=�Y5
�K��i�M5�[�J�A���>^zۘ)�!��(E�rqEO'@5e��;P�P����m	�WX�{B�T$�����O#�Gk:��Vlz=��)��E������a�hq�7p�xi?r�ǷLi�s�n�Tk���l�'�� a��#� �Ԧ*&, ��6����\��i
;V�N�k�6�%\���ٗ86����NBO� �"�k>YS7���arH��ɳ����_��q�x;��˽���蔳���*��'�����(�g��TN(�rYy���Z�,e,YT���cz�����B}F��+�E�9�F�->ev]�gqH(�$`*Sm�� VZ�XOYt�ׇ6�~1d��V^Y����G� �}����������,�s?U䑘f @�J1 �>��ă^ �W �H��Ƥ�3�`
f������"J���D���W0y��-�b`�K	@C�>��C��� ��οL�EN_�)�oj$��I���.�fS���~��[�>��9���lZ\����{� a2+��8DMl�) �������3իr�YU����<2M�<�ݺձ��8�p7�!Y�.�;�Q~'�}�8�oL+�����Rd�6���)*�M��g�5�4��A͍}_��%L����ҧ2�֩���`����}0�����Y��ҩ;	d5�����۫u<?��ԹV��17�
��/��I
��s/��^$ɰ��
�9��j�)������
L.�.�2�8���(a>�H����9D����P-�	��ǲ]��:5�߂vb(Q�S�� t��b�1�p+NtG��B��'#�A����V:�v(���hσ�@D���X��wڋ#=��rr���r㶫����Ǉ+'+� Ώ*�Bfɕ���m�0}����߶�.���-�?q���9T�֝�W�ힴ;2x��&ͩJ�
쏖��gN�vh�d��LI|�C�	>���tB۪2+�y`�t!��_���-��sAFD���ϰ�)FO�h�����7F�1�����L}wbNS���8sǎ%|��Q�և_[�6������9�v�0���9T� �p.��&p`��6�|��Bl2��.�Ɵ�� ��N�(�.��z&�����@�u4ϣ5��N5���>`��j��&PI�B-��nCCӟO�V�;
�I#��
�Į_ie!�wW5�!:����N/6k��X�^)z��恬�6�׷�Z�7@����+���Ųݘ:�������l�Û��@�40�e1� g�����g~�'��p�u����F�Xa��:[��$6!�*h)�y�,�U���Q��e�]��S������%R�*w�Y���iY��ܯ58	%|yIp��n�B���&vC2�kU����jp׻H��q��*&m��3��4E���޼�����vhq�X[�;�T���9�Q���5@�v�q�R�Nݚ��_V�/Ud�����7�i�%!LE��N+��Iz�׋���c��&&�b��b��n�G���8���K̲ y�g��|,ttߓY��l��m�>=�����O
=?���-� /	y�8����/4v~`��_��G�l�s!�O��_	(B�����ߖ��%Ъ�,e���o:��t�X��]�dH�a߸�$��6�q�|��G9R�<��?B�!�b�	=��t���5�Y�-�o�k�M�c3{��˺���4��ah���Kc�0	�FD}�Vv/ ���J_�(`6F'4MJ�`٨y)M"E1���������
i��Sb���Nkr��	���ȱ[� Hcw\\�D��A��ip�\��/:�7��}1�>�ʰ�ly���@����Cp5J�׹�)��U�C��>�Mg�m�����z_���l4S�QU��Y��VU5���(���d��v�4�+̸?��F�+��bM��wMz]�A�:�U̱a���ڤ�W:�4�ŋ�v�Id���m�tq�h1N��dv��9�$LE�#�������m�#�H�Ï��^,;�hj~\�LY�%��c�������:G�����b5��TgX��u��6�Џ</v�Z���\�2�`�$���q5���(M�pĽ	��Pg�H{����4d�R�T��Yr���,�FP�&RPk�:��W��w]�<���;o��`#���P3	9��ܐߤy��;ݣvE}�e���:�	r� ����d�Q�ŷ�Y���tt���m�8���oyڍ�4@7���T�T�)5{f�#��@��y*\Lg�e�Up �j��]6����Z���ڋY?UP��n�[��v������ �]��t�ڂr$�`K������ֆ���^e�@fث����,ٍ���V,�f��E���>����2뭳st�|N�����X��WmV��ls��j����2k��UO\���> �)��:����ЗOVH�OIK���W��x��|Ie��e���ѣ�{tTF�Њ�v��}�mMsP��%��K����W�)� ɿ�p�k�.c6K����2R����
2���ӧ&�1`�X���_���vw[���A|!���YTz�ߩ2�J)����J�����13�"e��V��8�D�Ƀ8�� }P�-��G1�6���S�g���H��Y�jN��2K�$�Q�C'�E>��N@B��w�m���=���D��z�"�Co,9**/�t���8[ǃq���Ua�Ė�'E������XG��]������86�M����7�t�{a�'Y���ƅ�Cy��S}�w$6ax�"c��4�q��t��	��[1!���~�%|>�#���-��bc���H؁�#xߵ��M�G�"��tS���̆]�L;��~1Բ�S�o���@X���/ݟ�s��,I{ �e0�4�l�����n�Q�s�t�W�p�m�	u��n[t��US�* �&��@�@�nW�[��o�~@$�5����}�y&n���i�%��Ў��v9щ� ;nU��Q&`|Ue�r�I�жƭe��VãM��:|�mChudys�{%�9u�S��J�,h��B�;�Z��t����w���27:�8.��M��覾�-�/	�D��f�?����:��KP�A��FAe���7���Ts�
���hw�cB�}}E����#��k��6lb�+�#N�m{�������ѧl�mS�ME�gqr���v?m�
�v���xok� �Ɵ�1Z�SF��K�^ȷX�%#0@W���\߉�k* /��wBm�w�����.*�FM5f�=E^�ǁ\�!�����L
�P��2l�/lY��J4J��t�m�6t*����k�dY�����݃��KO,�+V2�٤_w1��O�x"��ʹN��;���j�K�Ar/k�e�if��b���N��R�$V�u�S�:,Y=�d���m����D��]�Z��+H�������_�"��xA��?��Y���=3���I�|���l�,L�}��6�ƌ�9�4�#��{��0�ԫ/�$:t���N~84�s�D,����|br�8�q����j��I�Ƹk��_0:��Ku"�'B���:%�G�����e����3rF��]Ĕ��?CMܻ�;(���ߌ���f]0��#ȕ�#U����c%��˸�s�0n��o���4=��J7��g!��&�2ٶ�4��,�y&� 8�q)�2Dk�{�]U��f�
w���ϑ\��I�ԼVc ^��8S�o�sf�8���O�t�I|��a�?����Ŏ�뮴
+�	l�`�2&�ԻO�}�89��e�9����Vx�/�{ G�S�[ο�6�R���ʡW�x��fb����&�a,���yD�Q9v��2��ϣ{�秺3hZK. �[���ͳ��qx�)��4u=@��;;\7Q�	�{��Z���'�*�<�!��>�gX�V����V���p��b�!:�3�EdV��T�g%1�`4�@��qe�J%΅�y�]W��Q��$��#f��I�� Uh������"�e��J�,��ܮ��w����� �"`jm�l���⺳��~�F�yRƜ��>8㴪؏ݳ<�d���~zg4b�U:�/9�T��� Z�L�lU2��C.T?����vwߍ����Y�/�ml�����`c��J�A fc�z��L�3W�q�D��B,VK������.ǡ�^�zf��8�@L@�b�8���)8�"Bz4&��0ֽNb�ۈ��������垵���~?�X+2����+�uDo,���$i�7�z?��/��y�FU<2�V�>�hꚭ�*�"Y���r�7���J-beO�}��-*�Z˄+嵠�No��m��/�E�G����<��O������B��7�U:!#5EQ���g�*Ҡ���_)��ݛ)���K�@�Q�����ߴW�����x�$��	Xk"a������ꭱ��=yq��϶�[t�Hl��Pnlý�MؽG�T̠��}d���\��H�<���y�B�9��@�tsr-3��t�t56Gx0�X��$ >B`�����G-劤@rL�ps$sJv�La1�!'�D`~I�uF%[bPݯ��A?Ű�9�A�#����+�(F�m�w�e.�1.Br�.�r
N�d0G�X=+�FB���f+jD>��R �	��DR<�������Z�s�
LZ�X��|u����a����^�NZ��'�ZagdY�Ic���}�{+�5[��DlqH4�f]�Y�a���|јq	���&2������E-i]�A��I��mrj��T��Q�a��ݓE�c!�~�췯/�u����V�[m�"�A+�:1L��}y���pcw��5�F���I���0C��*��A�r�;�M�� �j��4|/��>Z��{�Y�tt��<�Z�a��l����K#������������c�j���>Z�;�x�nqE���	G�iyY��2�IBH�95�%���C��D���-�n+� ��n�_�E�z|�uk���G����k6���m���k��ϡC�@�.���UwKYBZ=ΰ#Nha�S-�����Rɫ����^t��D<C4����יj�B��^�}�	N��W�ѕ'ڢ�v`���6�ſ��8����$L�<���(Eۥ��6��TG*NbN$�'#?>��S��CzK�U���}���Թ|��n�~�4}T��p��n�W�ͳ�CYh�<)�v�u�x����d�v<�V|���k�����̰�j�D�d��}��r����OJ����k��6�+���D�U'��|V"|��ʋ9��Y�rQ��Y��%yr������������82���y|	�g�99읇��n���4�HTU���i��Rt7���v���<$^beZ�/��OB�J�o1�c]z��W�
-�&�c��zO�k!/$���t�Ҁ�ez��s�q�|�t^W��$�ߙ�h��IA`�o�uFf#s��J{.a��z�8��lZ������`j~t��)��F���ȟ�ݳ܄@���lx���M���_������E�1��M擓�V,=�~��μ��?ӱ��vNdB�ڣ2�z@aq:z~ݹ������z5.9�DZ�+r�,����6��7�=V;@6/��6y����A��B��UQ<�T�QxZ/�?��bYE���'K�D/�+���k[�&�9$�	4��q[~W�hk�[���w�@rɃ�r9$�2�j���<�90C�ڥ��~���P�i߂�,)��0��F�6�)KCuU1A�C��;$s}�:j���Ȍ�U���Q�MW z�p���~�
�I�y\�G����Ekm͌�LN�LaF%gG�^�q�ЙJc��}R��#��N��H��o"�߉bW
*0\�|7�Vۼ7O�7ƊŗU�۲�odp�-%J�~>?�N�V�J^��o�R�R�9#Z�V�c=�/�a��hӁ��V�t�As2 �ŧ�֣�mdC���i�2�����+t8~�@g��i���f�ud����	Bq�9N��Rd-5�@(���Y.v��ݷ��3q3����I��ب���j�����k�0k�i����~8L�2_�4��#��+����!ؒ�N���,y^N����8O����xR�h����ax�;��P��_�D�?B���'a~�E��F�sn���j�X���/�Q��e5�u�ѷ�x�}PD�y=���9����2�ڴ#z��.�؉.��������~A頻���`��&p��kH���8�d��ΦoI��hN��1G۱����������$Y��^��ug�"uѯ�8��2�D�/��]��f��:"��YV�=ԩ��g�H�4� �[�=A�f�6U��i ��t���Go�uB�
ĿX���3����2�ld�tb3m����h�J�2
<��ַ��3��H-�c^�I��̋s1�����{�nȂ!��B����N7�y��a�q�+خ~��z�F�n���uZ�I�?!t�w	3l�@~ڳEO��s!B�)�vp��l�8骖O�V���0?6���N�L��,JP̍G!�OQ��뇃z���4-�����r|�������7��6+�u|�e�LY~�+f�ꪲ44"�3�kYj��@eK�tb�����q���Bԟ^���z�ǬZ���7qݽl���n�}���0x�nЉ��fڇA��ӋCV
�rS����>�zPޱ�埓��f�ݰ�ɬ?oPa���L���Q�2�=7���Dz~_�����!Txn��$ �	)������p|=���U�M��O����G��e��F�ik�)�\�7`��i��>�+K@/.�1�8���'�:�/�Z��R�#��	�C�i�ȏa0�G�A��!t��	���=�hk�^��2��c鿻V�Ɯ:d�w��;��]���5lWG��P���F�m�w|z���.���P�ɂ�9@���d��x�8@ |��.�Q�J3ɺ۸,S���R/3.y���y89��1�͂)z��ml� 4>�_�JJ�z���1]��BG�,|�j>�O�Se�!7�gf���79aJ�p��PO%5/d�� W$��G ����,��Pʽ�C������JiE��,2c륍���K���8`'B�Oƺ��� wn�X� ��ٷL��e��_�c����Y�y�pP�4�X�{��mQ�#'=��n�c�Ik�5QTew���$0.[v��KUk�����τ�7M:48���L�\����V���`ME(qkXr�C��n�����	k	���Os�c���O��F���ݞN?�;�;;K�yf>	��l�(���;�+R
������S�ވC��j���{=����-�B��9�jj�����jy�
�����H����V��dtlεD^C톣$�U����H�0�c�FŃW��PS��P�Ӝ+v�
��Z!�M*���d���� ��֣&B=Ew�Jg;��)jC��H�X*��	L8<��0�p���(ҏ����P�H!���ܝ��
"���<*����s>4y8���~$C��'�/�*ې�Ɉ[�6��Y����NY7��bKSq7>������F�����5o ڿ���}d��\�����i�,��w�3�RyVs3��?���	�M�N;��8�O�*��>�53��P��Ȗb�Nr��_���y�7��U��Z�ε� M�a�IGkl�8�D�&���E:���냪��SC":P���B��?�hbe�LT�P�z;���"9�Xd�����O#Х?#�K����[/�Hۉ��o�\�.����&�:����2E|���-�>�&��%�WYac���Ї�
u"&J̭֜�Q��Tl�6�|Pj����G⨫]�Q7���է�A�׸E����X0�Z��f�[��䃳_��G��0�����+��H��ѷa��P���E���N�(JJ���;�ƙȮ3HnT����z�+�tK�����)�p@�<��-��eׇ!��j�b���%oX<�P�+���R< ������˂�Fe��)��,x%��.?�=oс�~v���N69��p�����Wv��)���.J�rp^3p�C����%��ȩ�9OB�5X���H���z|h�<y�D�6�9���#ܣ,���lw�S"��6J3Z3x?�H��7B�~�Y\�ͩe`?'��KhX�F&���DA�V:��අ�  _)$���u�6�s�?�B�r�r�ʓ�f����{֥F�U��cvo&'!r9�b���s����خci�Jcع]�%��Z�8B0�j�΀�(�$y�)�o?u�z���ܘ���/Z���C��Ry�A3O�ў �0o�s*h�r�?JK�u�s}H��%�)ů�B�����Q��|[���@�5����:S:�|7�����F
=u�+u>��X~l?��(��	��&��#X=
�>4#�5�c8A��T��u�A)%Y����Y1�ld��N���c�w���
I�
.֏E��ri�����
o�̡^?;Kד�|�P໻�z���C�,�L&���N�-�ϭ�W�Yr�G��TI�`�R01���6���P!���J�<7@����rԮ�ě_��Ǟу��(�� �!X�бfTO�6��܈�CY�w�k%m�򌔎�\��&%4�}�Q����Rk�1�T��Y}��΃\ѓ���j������q�`gx�t^~������M�¤��F3d1ު��_�ͨ^�Z���s�h�|m����n��2�xRj�#�o��m{�;st�\~Z�oS�Y�u��Uw��q�=��W��G���G:��
�R�f������5�Twl��z�K�@�1a���v��*X7�8�F��g$;�4�����I���q�)N�V�$$ ���+�Jץ� �ρG��jֆFC#SI�7E�^���2�\g��1����]���@c�u�8a�SfU�r����N�$G��L���г#-�xv�k}"Eo��O�D�O������(�[��s��1G4��s��>��0�ݪc?5| :�,�Ӽ����d�W��=��~���đ�>�Y�:,�=u�;#�>�9%�> �U�:�Ps���kqd�r��T�y�U�E���I�Y���Zn:a�9d_�Ex� W�Xv�?ǘ-��mÏ�V`��=U-s�i�i��<L^Nj���w�ήǭ7�$��xQ�2��j�/����
Q�w�%�;�-�M��4�Z��g�Q�=fJ�J)M���+�Z��mYW}�}}�����˕1+�a��V�Ő����\�N���w��N��z�|�x��|��H��}Ĺ���&2�n�±\����p�rϬ�JiMn��?Fx���qg���Dl<<qa/���u����V���^~9��e>�Y���d*�+g>h�6"(�"��q!�^M���e#{D��?2��d�4�ߵ�x'�׸�2���{�{T����;��ܬ�P�J��� ���W'hp	KQcV�̬��E�kI���.��3��&�H,<LςE���3��;�Yb�kF�7�YT��.�;���pd��ڮ��Dw�lSU�la��.��Z�y��]�1�[œ.�$u6��kJe�?dU$\�Wu�[�3�'J!_�,��G�+1s�}?3u�7u�����$R�Sc%�5���Y�`n���^��Q�O���wL��N^܌ce�~�Zi_���<p����~u��~�;�H���ݎ�I�|4eК��"�f'�Ā@�����|-���T:{O����Gh
��틴�T+�Y��g\a�~�Ox���M4�\Y/�K���݃b��]�k��&{�����ಱa�-N�� ��O��n�G�v�F!2]#:PU�C?�o���6��~��5�]�{ІO�zT~�S�K�H�=��uզ[?L#���fb��*�ƙȅ6e-��eS�jh�wOX��v]^ybK��&ƍXJ�\~������<B�%E�V�Y��Z8���/����rj���i�Н�'?�ed<3��Ƕs���Q���m4���-o���饞�q6�����W=��[==tG*���	п�>s��]��z�y���%B^�j�Y�ŭK��9����e$N[�/����V/�ȸz�Ы��EȘJi���~[��������b����mҮ�>�dƋ_�i��*���T��Is�c7�t���-	o_�eW���k3�5W��@�����xV��Nb�{l��s+��1$j�L����3C;X�\m�\���wpq8��+ԛc��C�IP���^�>�w�K{&:���Tz���4U���tk�"�jH#�j)n&��)C�@���O��� ��D�c-�p��vy�b:c媾=Q�=6�`���3P�﫮a��<F~rG��I=<�u'l	A�k�:4h�O���o*^%{����B!�:ճ�~��KO��Nܹ�ڸ�B<¤O$b�Y3��H��_X��9���ńf�� |4+c�Ot�2��r���Y��$X��C�#�-�>'*��RV4N)�8�W�~(�7d���tl�]X�N�y�'�)_Kw��1��?�\3���`REC��e����!�ݫh0q�z�;�S�4ѻ_bVxB���I@��fyN;>)Q{�t2k���),j��^O�N0�0� �����>�u� ����U�/M�O'sI�y�2@>R9Uf���=+˖7�b!���/7��B_E���L#�G�g���-D|�1ؒ>�[vA�I�F��_	�ݢ?"�WmTw��x�"���| �*|�j`U��1�ީT
��O�g7KvuS���|��Cx��2{��h��P��!�R�vV��D�<�Y��������_�X�Q4���k6w�҉ U3A�^<��/=�?TG�W��LWS,D��㨨 ���X�B��s,��~Y�K�p>;�I��&�'N��++M=F!��|��!��9I\h��,�T����ϡ��280�FH�U�N��Nҟ�.�X��L�ȧF�v��=k䌝"Y�w=�^�uH�Ԑ�P[��Z���e4ǎJ����I37�=LD���U��ͰK�������I �z��C	rY��\^�jXO6x�P/�[�#:��#_B�E�x���\i��
Bl�L��� "gDW,C��t��:��W��'�^���ԾV�a��vUj2֣	�fE� kW�@�u䈳�/��L��ݾ���Cz��3I��\�����W�S�;�����p�V![
	�`9�C}�|"p��O�3o{���/	��RwU�\7�n��S]b0���n��:ZjE��ݼy� d٤�Әʺm�Θo )���L'Wti�����5c��_�B:�no_��I�m�b��Q��)ѩ�6��!HvV��>RO|G��\ʒ!���դ������K�B�Г��U��'�JB��w�:	�����W��'ܑ����<�+�}�v!r�J���:(��\��n�/��ۀҖ^�x�l��An�vn�TLh5%��'"��p��|2p\�'��6ga_���´�v@��M��7P��P#��N�2��@15��V5��8�A��<QB0��KR�-����ĨN,�0�����r�K�@1��R��`�E+bwb慠A4�n"��|�Qm�\�\�A�:�o�{����7�ޯ?��ԓod��֬���;����ţ6���r�[�+�mmIN�M�lLB��\�~�}̦ l���fbL�*p�c���
����������
\e��<(4�7��x�{sRݝ  XX1���G��Eg���X䊿��#Lp��g���D+��;1��/ҥ���ԗ��߀�? c�����f��{�����&+#g�?������z_�V����w4���J`v�6y��v��%�1��
g6TOY~�<����N��`8�>��������{F�V���F�=�4���S����
�`G	1$����b=௏�a@I�Y={k�����SE��xZDz~���ݒ���˸X���0a)��^�+٣�~��4��x.X�.��$07��ِJ!�E�,�������r�~s�hף�f��x|��!J;�1-�Sk�������1�M��5��/��G�0a}S�Ta865�C�q^�čҺ��������SO�sأ"��kQ�ۺc��}T�'�5���u���+P��{YJ8c$ �H"1	q ��[EBICW{c�����#�:4�*��7#���Ȕ�8+֭��1��y��Z�\�X�n6^d�F���UsR?*�����z-�˚��*�A���W��i��p�S���Ī沬�9�%�����Ȏ}��D�D��.0�Xs�[T�ax��ü}���j���0,���{�BG��#�� ��c�� �>"M�t�i����k���n��KYU��Ԍ_��?��|V_�l܏z_�X���wl��@d��F��\����T^����Ex��+jnK\40M�O���m�/�]�;6U��M1�Ð1���Q�SS3IwJ/8��WX�u���@/�U�ޢ�8<;�q�=/�
>��ް��wnv����D������Q^ѹ�&�r�6���x�a�  o&�"�z	��9�<2q�!݌Sv�(#5B�L�����s�qlݨ	�Y]����Ơu\�-~�g,b�����:e�ٌL<B��fvI��%��2��1rz�jrF�%
��~մ�~�%d�A=nO�t��a�S@yQ�,L�DnvC�7cF�ٯ���o��G��N=����Ȱ�h�W}~"��lC�6V��o�������MI��_o\,�=~��,�	t���sɊ�YM��Cbc�����sK6]zNȕb���#]�v����X����V�"hcj�d@���ɲ��db7Z��*IW���w�M��dD��E���^l��k/�_�P!f:"�!N<W���X����%3U1�Eֶ��!;��&t|��[Y���*�O_������|���Y�y���N�����B����W�ƀ:��NF5Jd\�cX%t�Y�u�!\��h@*ͫ`�m�R,�]S��N5+�j7�����[b�����}P��8.��m�Î$:'Ȧ5ۜ0$&��^�B�	J�v�wQ�ZHN)�g�[��V�M�x��0�BU�n�8W��6̤ ���j	Ϲ}5���Tm��mRe��� !>o11����_Y�
2�	Jk�"6Nb*	FIa�u�~�IE�>E���ҤG���b	�P�����ףم�5p1D��άP���\lS��l��I��aX����(]D,�I�>�S�F���
H' ��(�9{�����z����Ba�cS�-IH�6W���Y�v�-B"	=&����R��Zd0�iwߵe�J��K������֓bK��[1(,���)�G���ea������������o�_O��+�R'��JgɈ{"� f��nHg]��x��U��9t�ѣ�%�'|;��"�|FpAG���dl�������{��F�¢�S�1uEg �H䟩�f���ߣD�}��'�痆�
�����1<PX>�R'[r'/r� �����R�/�&{xm
u�O8�s�X����S�=ە�r.O���No.�,+�WjӿV��-�x�BЅo�
��<YOs�p2z"t����!:<��-���I^r=@Yg/c�aQl�=�!�_�Y����w�ċ�{ߚ�k�l=�bO�gq����G\Gu��<�� nza�/���o�(�Ʌp��p��1�A�`�`�d�@�:�,v4��G���]�.��EY��Q�	��O2�TԴ"�<(\�-s-�X{�D��҂A��	8���"@��y�Z]`4ˠp��9 ���Dp�-���6�6�K��c��*4e�*뉌�=��Ls�W�M%�3�a����:��уV-��A	�6�<� �@�:��5��1¿f�):�Z����i4){~�K����9�����!tAh�-V�66E2���+[�s��{�D���V���J �mVYp����I����ð�{�h3����i4�u�5T݇.�&:�6���1�-^,T 9o=�D:��5���3�ߵIW$�T`��4sp���o�<}�׷*d�׆=HW�bK/�g�]M}���9d�$��e�E���ڄb�n&�Om+'��0K�<��o�(Ʉ�r>��q�e�ҙ�Z�C.*/����(�j�u��i�0��]Q��}�Af-1<�^��&�С@A��
�I�6&�iv���%$�w[ RM._���9�sQd�y�g�	�X@�fC���.�P�#_U���^ F����� ���9�<a8��@�wT�#�U�x&�\o��j���͋g���}0��v�@Kǁ��C=�
;�������S�'
�Bi��� <��P`4���`m�4�S�j�:e<V�Y�?�	����� g����g䯱n7|��]N��wI��� ����)U���d��Sޮ[���dOE'�Bb�fV��g�G��c������k��f���=���HC���ҁ�k�a�w�U���e��cT��1�5�]����fGD/��I�7?��Å��I�r�w��f�ؕ�C��C,B�>�ͫ�'�x�������l��ַ
�q�ɽy�һ:�ť��w5,��rF��K�� ̂(�ls�l7NAP�� ��j��4,2���vj �T�������F�H���t/.~�B?<Ot�%�:ֺ��)�rpK��êj����M� ������	0DU�I�r%��^��å����"J|
X������Ǘ����|6*��y�W�s��-����8����`w�,��?��\�������]�UF�"+s��
n�.+D��7j	A3�	�Nu�I}�CJ�T�D���kro;[)�_�Yl`��7��1��d'�<W�%����ni�����J��..kG�\�|]:�nDЇ�2k��|i����{�%
�lc��)���.{ e���ퟁ����L<�,�u6�����'��;f�#�ULB2B���,:�uWk�X�w�h���DX8�cN��0�h]_��]Yq��E�փK�w�p�����8�d��U9*$���[�k�hӢ��'��¦�����N����"l��`��W?�� ��{��$PCc}PA��HI/���
�ؾ�5
��8�~j�qS�Ve�#�f1������D_�P���^J��'���<:3�y�@^��� ��s����x\9��J�L��c�����$'�(o���Nc�3.�ALQ�������i��>Ζ�������YU��~Č�ɪ��mb���_��7��D�V�C�4��.b�t1�HW,��҆Wqv"L�����Vx���&��	,�iZd������	����7v�iG� �����S�Q\�-�+ɓ)�v�9?�:�B�$Ddg�i,�bS�v����	_1[�'��V��&�
�0�z��k�!�b�՛)�y�'��"�{��sbL�o�7�;���#Ei�&�~��Tb��?\��@�\�<>gɰQ�/�c��b��%�W�v��[4*�u2��[�0�W:��)¡n��@%WQH��8;��+�9�U}@���j�]�;�<U�lQ��D�Hݺ��<�I1�:��aN�y�p���D�|�U�S����J	F��}V<�	qY|��`#��"n�a9}�[I�Aџv�A�{�,��Sѣ-7���x����N'��-�j}�ֵr{�oo.FCH�ӗ���"�O#
7~j��(���DpU�� ��}���^(H	\�"
rќY��c�x�4f��k��"�h���ɼ3�;��lT�MP���f�7�\���9A���\�
7F���s������o1i�4rY6!����횪�ʡ�����He�uf��l�u��j�*b߶,/�w�zKm|����!���M� y"M��O�C�]\�ip g�R����U 1𹺡�I}�c���gK&�@�9Qp�<�auk��6��E� ��[��UU���/����t��g����SFqr�]���N/�M��LK��˜��BCK��M��!�~rq7x��Jg�+B���-��$	/����7�h1��7�&ه*�bH���0g���(���_ֈ�Y��q��*zF��l��,���h�����e=��YϦU&�7�T&=���������R؞ޙIƸKJz���..W�8*���{}��%�\k� ��V�3d�#�l�A����ڢ�
=��ϫ�� �"�wm)��3c��!�q�c��#�zI"���Q^ʱ 	���_�9����Q�񧸅WQ"��E���,�.��� �F������Uш�ZF��-�[M��-����YwZ{�����kJ��aQm|���.F�(ߞ��9�ОIYǍ�5:����ބ`�k��w����o�A���f�n\B�"-�n��	�:��1II[s��`_�G�>4ܴ�k<��_�ԏ��F�R���N�ǎ4�e	�=���L{
�1�V�5ޑdSJ=������C�N>ț�Jl�SY���IY9H}$K�h�@t��Gp�M�S���>����i��-�a�{K�f����z�HRYM��$T��f��>��� }�Ħ�
��S)��ػ��sDi[y� ���ZT��ϓ;�Ɉ�������X�X[gc��	K�ģ8`@�Z���?�.ԧ��	���Y��)S�k�q��g0���1��t�4|؄��ٹ���S�<�#���\Y��s��
:��͚8��]	�U<�?U'�e��ĵ~jzfm;�&��� �Ky4ߵ	z��8�ZU��l�����͙Z���r�X����N�$p6mV���V�?H�.['�n/���E+��W����~lz^��݁�ϝ&(�f��1v�䝝��954��6t�⎾��W碹�OJ��e���0��%����>�T9U��J!#U�^k4�+3!�6�^Q�<���oHb�?�H�h�֭�q�bʦ�h.N������)�F+o�H��'���,��4^o(�B i70�ֳ�۱�^2��t|��c�=z`rZݙ%Γ̆Own�<��(%-�_�z�uR<eՃ&j��Fh��v{wJܾN�:"�{œ�(9��1�?��X���|v�Vua���v�M�
@!���ۑ^E(�R��w��<��m��yv��o Kܓ�^Z�����'f6�R?uW>��BcT"�ɖ![RQ�x��^��UQ}2�%����,�n*�2�c�C�x�3}��`n'�J_Z��ӺL���Z��J��e�;B��"/(`\W�Oj5�ON^�9��pP����@��W�P�n�$
��_:}_FW�����!�v �X��m�����"q�R4(��'��^w�'�0�-��K�!?�L�M���cݥ0euF�u3�!v�V>2$����OeR8t��d`p�
R�x���~qA���=�?6����T�2�\v�����Lj�Hf\�^?��c�uV�}���Ӝ��8I�����@�}��ߗ�"�7/���&E2��mOu��0�Ĳ~�$)���I����]Q�Z� >�p�����vԘ�����>a����R�#ZR�G`��YjIA�ٵ+�N���9���*~g wtt�`jN>�������/�@������y!�kUC}�[(�V� G�W{*�H�9e:GL�nqǕc�����P��e�hG���i=��]��J��ձu�Q��֓�.1��X?�lx`*�rL��������Y�X��uݢ}��qt	�6%�WM� ��WtWV;M�C��z�}���Ֆ�l�Sq��O��b���l�|{ @��G������qb�l��l^�W�/M�&��]`|�,�<��_?�[��VB0��[�����588����C��
wn�6K>�"��z1�;�~c��-y�Z�������a呙X�2J���D	1��r��џ(Nv�f�̖�{5�߉ag�Z��D�8��[��Ԇ����	���,8{%��7�ݶ��|/)�^í%;����ݼ8����f��GuQ��9�'HXD�:�w����z� *�.�<�[��ڣ�Q���Ra*�BIe����&�ܣ��x�, ��^kj�u��k�{_\Ue.�{����:c����������n�F)�6tbZ�w���(^�\uqu9(�9���,rwT��������|Fα�&f˽���:'��5��Ÿ���B��H�V���W�����g��0tVF��B��mojz��5�3�o����-/:�)	�j�T3b̆�e�B ���$�LpoN}���M	�4am�'�x���<�X�W6$@���t5�B��o5ID����|�� @����{����-`�ӵa�XL5�������Y4qÅ�@�[i'*;�0w�cPoZ"t%#��Π8�H�'~�I����:�N��3�b�[7}r���r6Q��)�k˝��?�x<���&�7�<_{��)ۺ;&T���,9?
�hץ��آ"AOk��E
�^�xv�|���3Hlէ&D���Yھ���?/+bIf��S#`���K�|�r�����@'g^��;ה�MA�
h��据��	�J�0L+m�\q�|�0t�.Xcٞ8_NXu	�>j9B����*�ܰ��E�bJr�I�SiP��'�غ9k0:)Z�F��P������ŻU�����:��{�ƣwꋊ`���ve�X��X��i�x����̶�=ķO{l�&��Ҁ7�9�PX����iE���/��1�-�r7�W�[�f}ԁ�����D﫣n[LV�����vl*�J!�].<g�^%��' c�:S�kjD�V�O���y!ǎ��{��#���8��,��/�Nh�׷��t'k����!�n��%�"���1^���S.-�V��G�L�qiYJD�45�:�*	�<U:��3#g�<<��մ�-O���J�Z������5Bjʒƪ���F�E���ɍQOz֤^E\�Mח*���q2e��nwN���;��]�~���~p죊����� h�SRn��pK�b�ȋ�o,}e5��_��2���b�����(1���^�_��hIM'�Pgysվ� W�O$G�[�b\�m��h��z�i�����dpIxo�c��6��������⾩ �"Y�LJD�Ǣ���%��.i%�#�	7#vz�c꼿3,r;uԞ�}��g��pP���Z-O��fť?���m4��m�[��*�1���
+�X�]T���ݫ,���_�.y
 #)_��PK����-Bs�X@r�8b��;��XV��A�0tf8pA����u�wG?��3y�
�TW1�Ŧ�#>Mo�F��G9iBL�}%�*B	����[	�h�ky�Rk�J-�sHJp�*�|�)�
K�KE��U�/�(�7�RS%,��mAj���V�0��A������Ʉ�b!q^��P
7��9����4���*[Re����9)ܢx���@Eeϊ�#��S��mi�f�0� ��e�i��<=�8����Ϳ��?3q#K�e�[�Ʊ�3�e!۔]!N
[��O/1��kb��'��J��c�&w�Mb�5���^�W����ןj�W�' �~@��Y����l�1>G���z�
�3�6��O:\1$L'cI���l�����3�t��pΜ�����9�K͋���B�J*����mEP�!mH��������ک��2y��>�7�T���r7�^��nvMW/xa�Lz��@`���A ���`~�[(+�p~���7��Ҙ�޷잖e�9h��~�P�IDk�f3������<c��y۵"�~�2)��\�B����D��/&Ǻ�S�����e[�ש�O,����4�Ә���z�����H:8t��$\�1�k�eq�w�<@3�"���|Q�E���:����y���= ���4�e"���G��(?�[�y~�ćH3p�O�[�P���FSi��
v�D;��[����j�|%�J���	��ش�3Zߩ�ة�ځar��1�v���3����ya�ķ��eߞT��~X���E�̕�Qf�s۷�w6�b�p¹���ϭ�(����Bѻ,�����j�F�#xt���9�a�z,x�ѯofU�����f�a�2��O�o��
���$�[�$.|�P=D�e�\XH<�a��@+���M8�J��?�j�tK?�r5'm
�v�\��Oķ_��!���{M�Rc-R�p���]^~�>�ٻD�[��$�F�"��w?���4�PxG$g�p8�|���Z���yG�;�y��n��h+,�`��v���dD�~�&�W'�x�B��/�����S�� 3��|f���D_G��1(㓆��[aSoIU؋4P�f�he��f<���8�Mb�'ت�eb���A�����k�Fne�������V��aA���U�~5e�y�i��d��/����R`�R3�Ύ��؝c>��|r�$ě!/K>/f�S�l0c����9z7�9A~D��5|�aHq`�ȟ�^%��*��
W�G�<C���j�-Q�nRg9�:N��!5ZU��;-`fD)ua�;���($M�ޛ����
��ӓ_(�;ˋ�9�
��D�+��~R(h�cM�/�����꼏1=�[��9i�!�������s��+�㇥�yR����I6�˟G�>,T;'֦0�J~����v����]
��:k�4F�7DTT�,s��R�7��Ž�-a�.@P�����T~��"IC�{n�2�����o0����&��$#/uِ"@��I�9 s��� .��?��g��,�V�7kai�Kï�9��u�G-�/̡��k;͒�n��Q�n�y5eE~;	�U��?�v/<��1{�Ɵ%V�k�A��������dV��e�2�j��oN������&��\�5�q����,ҝ��D��g�̴�(w{n~����@����1\^�W�fz�P��0eϳ��V�L{p���RV%x�ܑE+@gz�Wک�T1D�"Io ��?��j�	%�i����Zn�̤Y[&�#��C��������������3!��|��@�4y~���	:�}A�j;`Rk�����{��B[�G)[��*
o�4H�qz"(��SZ�Z]q�7'M#�Zԭ���݇�3����c�)N����z� HDz�Kf^ߧŰI��$Kh����7%��{Rs<K���Yk ɀ��#_���QP�*�/U�i�Cߝ�5+J��ȞO����&R�������N���
���V�P���2Q�$b������C1��~Ks���[Çx��=p��[5vA�Rb0�w.t�7��5}l�C�n]cҊ�Bnb"�a���s�8q��4t�L>���=�l"+���\�`���H�B�=N0��m�Ra�y~���lzr�mV�i$V�@:6'��w����Ϛ�'SlL=N�ƂͲI�@��^�<G%�Y�;�u���T�aߖ���Ǣ�	+�AoF���)\������ �AUs�P<���8O��p����k@�4���
��T7�9�["�#��=@x٤{m��Ҝ,V�5*���U��=��EO�ף�E��?L �OS��a䲄��fH1��A}��١�sZa�y���C;=T�nϯ"i]c>Ni��P?���.M����9e���czA�meF
�'ۗ��k&� -rW��˭�l9����*r�{��cS��w���|U��x�?��"���Xy�2�ع@W��B8L0~�Y�
��F��6��z�HB1$�{7N�m�EǶɄa��h�4�r��r⨖�P�@(2��o��%�^���\ê G�aH�ޫ����@�
�=���2у�dk��ou'�����!�F�ii��lGu-��)lf�>����1�,8pt��g9�}gS&��PONN�E<;���D����en�{H��,���Z�P���;��Ue���vxެ��4=�2��Kl�h���g�m�j��C���\R��p֮�Sd{�����h�L���'��y~~�X-b<�
�"|�VV�!i;3~ԫE&p{��5K�j`Z��/��c̙�\�H��	��r8��g�|)��μ�z��	�=f`�K��uJ�9��{��:���`��ZT���3�J���1����G��<�iF� +�g�`�c`�QۗaD�w�K�@�A���n�}�̍#���yZ�G�/�2G��ԱP���#�-or��0�j������&N\�z�yD��t���v��n�����C����qlO�������f�ԩOp~���;@����0:�v���"f�6,/�!�t����gi��J|����Q�6RKI�͓�q�Uͷ�%��M��� Ìor�~�R~[�E@�D�n#��6���Z~m8e�I�C����X��G�%�p�f��3<��Ύ��S��Y���d˙k��.F�:)q��H������ �f �b���]S�<q�V ��Z蠟�gZ?GkRBr~��W{�R{66.�u��C&���Ԁs�:����~-܇v�e�k�Vپ]�5.(�cy'�G�Y�?��QM��[�Vk抿�-#���u^��m�}�Ԩff>����i�e,�y�Q�\��+�&Wn=�I�䁨�-d�B���j-��$����E�\K�}y0X�;����/z:JJi]D�qI���e.�%bg)�����y�SE d�y�
�1�_����j�3G�f[�tx\F}#�"�1�q_wA���8j�O�Y�d�p�f����8Aۥ��9]g8J~���%�K�S�Qak�&�%�����J�����2�k	�Pn���l��Bk�lJ8�QIy�]����g�7��'ɔ�H�AM4v���	G�P茐����s)6��������+��m���s+�>0�=���?ʑ�0b
JǏ��Hu�ڡ�V��Z�4��;���1��㏑�&����� �9�-���-sR��v�N�g�ԓ�G�?x��a�&[��0��}�������h��]�>���U*�3�,��?�;g� _C�-MW�S�c�i���
>PCX@C�Q6OP�-�����߁v�K;-̃��7?�;NBbh&
�J��ʑ�Tv�x�߯p�?��!o�)ț�y�l69<���1j�r��4U��R9D��eU�@<�a��+{r���tq,Y[�a�
��]x�n�v��t�UՆ4�]{��3�:+�����f0:�ġ9>�s��)cN����ϼ��zE��ĆJ�a��H6��S��&$�Eh��_Ϲ,o�}[�m���Kv�v�|�'Ef�a����JV
.7��_*-�!<��U������E�΀�)X�wP�t���gy��g}�^���5��3�#8l�Z&)�5��}1�2r�
	z�u�m�(�M���5��;^R�+��"8�C6��{9���?�	���� E:(���a�.�[�u�i9_hèul� �C���S�w�o�"*2C?���xK��8��}�nE6ޣ�О:}!yP�����h����ۏ�֜:�4�뿏mC#뿬���b����
5�Q�V	��B�NKO\Y!�$�"��e��of��%�i�N��P'&n��|O�.�2^P���m�Ag�6z_��с��J��ž�s��� ���#Yz�<����ȥ0.Z�+����bSR��fn�#��lF�ǀ;�oqFB�&D3�ftrǱ����r+ �'�3��������ȅMsڎ���E|p�z���lRJ����0�[ͭ�[~w�1\�!�'������2��:?12c!v�lb��c�3�o(�g�gJאO@U��0k����Ʋ��0�D5�	��Z�_.ɡ.�[�\QSc]�%a���-���>ѽ,+<ns+FR㣂���!��#����[��K�»|��>�N��Xf���ۓ���o��(<A��=a��e(�x��磻���8۹D�8ԜF'(���H�W�j���!.
�jlI��HC��v�����[�_���Zh%)ɭԇD.�Q���w����QO=h����`��ʚ� P>+:"�4�� Y4Z.�/��7�,�دU)�������{O�	�N�Ϩ��\�	�flQ�G64�����66���)��qe�������e��M���l�aO�<,J�v��"��\s#�5��O@�"֤�cb�l���oI.j���2���.��Z�B�w�o��,���G��>�*�����qIEg�*�����(�uS���-)�z��hU��;��)�m�Je�|_Y������"��D���c�7�P�:�	�D��/��}%�)��o6����]�
��(L/�z�}~�����}��j(�JXǐV����o��bɊ��y�|^&�&HX��R���L�8Uttm�e��ʔ��xqٮ�;��s&�`&��Ox­[|���"J����d" H!�>�1��tx�f~���-Բɒ�����~�'���f[�Դ�e��7�X��L�*�O���1�O�*�������ĹP���<V�w<����	��F		S���N��4�(��Ȫ�M(�``3�*)vK�lw/w/۶:�3Yr$�.d��hDJSM���m��P4�\p���k�R��BK�պ�N-c���u�"��Q�<��2������v�Q�$ha^u��S�3�mG��$�S?�uSQ�$׀=�c��V��D��P�=xIj��9���gxh���8m��w٬��󂍗w�J��c�|TѴ�{�|X�y~�� .��Dw�AnUe����ߗ>������75�I�����]�����-U�h
'��#Tu��Q�j��$ĥ]�5��Z��ԃ�UW�9v.�>�7�3r��C�,t�X��Y��S��GD�o�9��p�.Ē(���kh��)�ܹ��k��M�P��\^��w� �k�[�>4���z@�X6~7����ٸ�,��1�n7��ߝ(���JL=�$�?韃�'5DN�x�!$����0�R�v�Nv�d~�4@`Л<o`!��_aՈ,�5��8pv��),G��
�I�2�u���Z�g�S�Z�E�){p�Ħ�v�0|�.z=��	B�q���h ��\�����Apβ�R(�Q�&�ȊM񁍹3�]�G'5���fM���RP5j����WN.?�_>p��&�eI���V�������s:��������ds��Ny�j������|�<g������ebLOm-;X)���*S�nM*�y[��]c,�xr룹���}XE���.3�0b��ԏ��"�qYFO1��i����f%�nP	�F)�m��Ջܠ�埼G@X<M/b�h>�
!#Z��e�M����!����oͿ��U��hl����n�7���8F&���p�j��Z�<r�h�< ǌE7�Sr̲|�:Z}�X�J>���v��`����Ji�_9��~�^r�+5�"U�CS��a��\��JД�ĉ�����(�<�>l����(���$
�����;�1��?��.�^�<Z2�qn8|��*������Q���dtկ�j3��d�ht&�W=c�	md������}��V8���()w0�̿\��A�YۮX�ɠ磟���m\K>��#�
`_(����yZ]��>��	������"���� '(�ہ���Ur9�,c��8f����`�$���\ �I+�8�А8б:S:9�7�#V� ��M�����:!h���wh�E��f�>�	��@[�q� �>��*�S�P\�i�|��G�X^)<B�����wZ�\,(lhn��w�d&�m�~7"�q3`�?B��#@;��`tNs�"= �)Bp'�
c��+�T)�2;Z�k��>r+�Tq�!WrU���i�hۭ�� �_mpHaw�	OD��3��K��4u��s��~�XdP�q���g�|�����$=�7�Qy}N��{�|�pM�������7�xC��^�Pz� a�K�"X/�>ϫ��Փ�~3�������}%}˄Yv�j�
�b&*�E��X7K_ZA���5D׫�QںK�G7b[��8����8OHK� R�s+�@�/�����
��޷�i�c4�X-+v3a�"�A���<Oll"�v��v˱0׺9w|?���k`��j�D���>��	����2�&�Rİ`'X��M��[������q��8���캳��\�kY�N>P�[�7��]gm}����1�VY�>`k����ш�0�O1��V��y}���Di�~VQ�ikq�>�������@W[uh���}�yC��zZ�@�z��'؟�S�י�l��;^_�cuUI�*3�[��f�7!���l�UIr/q톈�ڥ� uuS�^5Ե�#���R�CK8:�;_�)�׶H���ia��C}�4UG����F����Z�>���/�GV�i�գ�ǚ�tS ���	�W�o�ɖO�]|D-!6�Ɣ�K���-�b���9��-8�C�1�䷁��޶%��=1��ȟ�KQ�����_�f���M��uo}�w����1ԂB,+�(2�g���L��Ώ����>Y��{�o�
��N�ٞ�2&bʜĦ��j����u3�]�Wr� /�=$n�6��+�`�¿���R�*̌� ��+!fW�|��@'�c ���ټ?}�Ǯ��k�%R\w��\�$8_e�<��7	�3�,�_�-��=
F��C��^�U)v��M�@Ug9n�C�ڃ{���4җ)�ip�IX�}�7
%P�2���C��������v��\�IjCb�&E��2	m���������f�,`[H�4�ӱ���T���mD j��Ը�C^�u�S�] ���V�_M���'�)� K�a��>�t�8e���T��:�(a�� �c��Qе�U])�&f����)y��"NgU#���r;YT����?y������՗�#����Dw�PL Ԥ6Ƶdʵ��*I �r�y��-���Rg�\�P�XF/��/�$�����&xHq���Xu�.�B�����3d3�W��;�o���kJ�=2�|�	���he�3��Y��g�
���8&�ɷ{�Q'�Xr_���0�,��O�M�G��3��;��Q��`Z��ʐ�a*�;����G�*�L�$3�0y��0vE�ȵJ}.�*���堀l�$�k`/V�Kf��"�ف��Q9���Ke���P@$9��L�6L�	���M[jL��~�]������`A��ؑL����ԻT�Nm�?��Cu[�To�[63�,�m󃭍>��]�;��w��I�ms4ա��Ú��lp#��!Hn�_�N/p��ρ�no>�}{ޓT:�I�������Xz4>w�-��qr�}�g�����w��Y���>ɛ=�;-�-�^	#���d�ҹ�e�u��M�T�Ĩ��#IB��*e�M/��������]����@b7�"����+��'ÍΞL��Nؙ���M"�����]1� ��<�\��⬴�{��%�-����̅c@�׫�<�"�\�W/�6�9��p<Jj2]�UU�<a���iE�W�7��`��{Q�������? 9/����	�pǕ�pa)�c�l^�v��j�.��/�
��XS=֗�_q&5�'����&f�p���_��(�<�F�*R��I/���n�����&���f��M�{Z/�S}���A��`�	�=h iI=ٱU��ʠz{�e|�����3)~�U�#۝��#����lP��/]V�WWE��T��Tw-�]�Nx�6Ȼ��0Au�@����S�"�4�S�����\B�u��i�B��:՞�o���ǁ	NDBM�ڑ�?M{e/ʎ�J��� .V�e���`�n����͓����&����8Hk�)���0�@�����&3�?�9
5mA��YJ�'?oGZ��)g-�J�O�^ߍ?��Ƹ�.a͛���k'gt
<{|x\����7N?C� e!l6���bg�+^��(�����LD���uv���1M?��$�To+F��+�7��g.ڳ��{�yG�(2HM������:b1�&���s?�Uȼ �AE���Z����W�G�@$�t���A�ʺ��O�x�)�v�d	IShbi`Ǥ��6�iʭꨀDb��[浍[��w���ސ�Mk�քkHl%����b��� }loqZ��!+�(��¡��p���O3<l�Fn��y�� ��e�ņ����E�8/�%�pD�{��������Y��	�e�x����ןڔ����٩M�ckb���L���<�g���>��U��A'���w�ݳڹX߹�6�V���� �Pap�t(H\������
�uGy����	���Ev�H��[�Hvq� E�g�������K�C@LK�죃�be�m��.�P����o�}���H>�ޗZ#�ܥeů���	
C$%�)�^��
��a`����x�0�5��]�����n8]����%��xJӂ�z��Y����h2������33�y =�!gKA��m7�
��µ����ʎ��)%.v���kx�2c�����O�jV�/�I���\�G��	�kء��G�C��/V"z0���g���-?�I;$~Ѣ��Y�pvDe��?�1�:�����gr��g����fӵ�W* Y^m=�	����8�X��݀��qAA$�>M��$����WMЯ�.���e;2��W��^)Km2
lI�_5C(��mM��A��ܪ!#ĖԂUFJ�l+_�RC��y�I1�k�+x���<��~�D�	��6!��<��T���1_��`W��>|~�K�k���I���9��1-�P'��U{���~6V���o�ঔ\�{�;Z.f�����Hv��y9�M�G�p��J�h��H���Zұo�z?�_��ޠ"��^#�Ͽ
O��_�t�|�:�g�1��Ҍ��و��� O�ɪ�i��ԅ�|u7��e�A�s�އQ��$�E�BQpݞ[�бz"��j��?;Jm�#VA��!���-�!�|fJo�c۴�����4e��>��V����(h�P�r&gx
�0�?�*���4��Aϋ�A����[��#S�9]�V�[]��E���ɹ��@�1�Z�銊r��m��R6TKl�펪�a.�S�m��K���(<z�'�*`W���Wti����nLj*�,p�?�~��C��N��1���"m����Z�n���f��.q�~G3`ݟ<�Z�W�|҅3��~�!��4
�8�����fg���OS�e�O��(���� 1�N���40lM�9~M�zV��A�OB毃S֏uA(�j�V���_]D�@Y�±�g�C��� �P?9,�V�&ʱ (������"��#���g���G��[�P���S��)�1�|N1�n>�����H�
�V"���(`\%TOI2H��sA�g���O7�����\�
Hs	¡��,L%U�B��v�l����"}/��~#��M�oI1n�0B�¸�� '��7o��Z�޽���^�hˑ�o��og�b%����~�`�	��2��C励WՃ�0�Y��K4����Ǔ�Ć�j��t#�"�������*�[���Ǜr^�X��h-)��d�"M���m{�Ck[���f�[ssw����qK���O%�8�΄f�Q�^&��{N�F�x�̗���ں�R��K*h�,B�ltF��s]�M��0y�!ɒ��f�{�N�����Dܜ�:�f>�����?X��)?#�)��*aw���m�F:�|.Z�:	B��r��*}l��YGv
̒�I<J.����w~��JIǠ���(=_���;���8u�m(t�j���5�v�h��Ro�uL�6X�F<��ܧؕ���EMa|�R���3t����0����@v�]�gA�J� ���_V�x�^Qb
��F�O�+`���xH�����d�[d�)	�Ɲ 8���a��g�Ѯ��Q�l�/��8SF	�`O_F�!�~�����	�M��_��9���"I��"4�.�
?�->�px�C�ҘHe҃�����|�c�ށ�+h��;��;ݣ��
�v0�/ʓ-�E�7C'K6�
U@+J2��С���b�>:S����;�ߺr�'������0ol,%эJ�3U�7-`�=����uu5s�L{Lp3��_Ґ�xZdژ�%|O���@��_�8�F7����������S�x��83?i8�~tŝ�"�9��������dri!�e�N��j��*DS&��8�6�����wb9�#(�OcY�!E͆�;iW��RL�t�[���Co��B�V��m�ol�r�
�'*�2���H2�@f���ޝ���*n^P�U�+kh���Cd�/��3�L�m9ׂO?��$W�}��BL\g���`��7��S�D�&�GNJv�Pmi��0�J��O�
�P�<l���T|�d;��u,�����z��e�8����jm����9����ZsK���"�����dȮN��(�����Ζ`�D{���� -B*�mܚ��X����>c>�#z�����yKx��=�k+�՛)��;s��Ed=,5�Ȯ(\�`�Z� ֎��*��
0I ��-tڥ�Y6	P�L�۽T�`bd�V��)������p�*4x$��c�ei�f�ْ;�o����[��&�5#h��Gk�S��R=؟,�8og�ܲB������A#��"��7{*����3,k�&�Hɪ*�l#C�?�y�i�B���<d|�~�]���'|�7ږH���S�6�ۺFB����v2�ص#nt(6���@=t��z�<�"�@����D��i�b�,G,t���ȋ5sc�;�ߔ[jh򾵮�Q�ƈYZ����H%�*vSº)�%�\�����h�d@�M?��L-���#ER�iF���*��D]�K�CJ����&�dA%��k]�j�}���[�l��w�7߭��#�Q�Ջ����,膵�9>����2'<	��$ו{����\7�F_��hQp�����Yh�(�����x>ٝu@\�񆀬�_'$�~��\#p�Z��]� 	҄nݖ]��%y#����	YFX�^p�+$T@c�U�H�>��2Q�#j_e&����}��N�.��=�Jwc|B�$wG�.�(�}^�8`��Q��O>e4^+�S���E�(�+E�X��%P.a�֟�7�ɤ��#�5�E��AX;���������<����5��x��ɛ���+
Xi�@�T�8h����̄P��&��2tg��y.r=Q��_�� �d�ٝ�H�}5��_jHhݬc3,Ńil:+S3��P4���eȜ��▭���W�6=��c7�3͵��$��nX(����!kf�T����[ز�ëW\3�8���āo۫��S��Q���1N�T<{.�u�.$'�ͺU��Ȥ���$>D�5M��bp��or�W���A�+�B�0�g�4�@ABYY�J=�r�7'��Fc�n\�����C��$��x݂�
t=!5�h�c���L�4T�Mt����m��Y���Ѷ��!�(���\��qMp�~fL���Ѡ�g4�M�s0p>�O�S:��l��%�U�T/6���q̈��X�t�E7���;a����T����,_lD��#�N��wZjD�^���L��T&@,�uih�v���x�#���������
�7�r�5E8l>�w���0�,�$��󈉘j]�:M���K�q0��V��s3}#0��9#kؾm,h9�շ�����JcP<�i�'����I�3���n|���.D�� .��K�{Z��1��	�C��i��9=�>��QNQYE!+l���~�E�Wѣ����G��:�eC"�7�?�@�	���v��S����{���Q�/i%:�y7���9P��ńFu#1�
�;CY8���YPyU�'Iz����k���z
0`W�2E���i�{0�(�05�R׆�-檒�9�t�8!�+J)l/L�����Ă�Ĺhp�Y"��aj+ �`�����{��a� �17�K+���Ļd�6�,�d�(TL��-q��p5��7�`���_�}]��ǩ뀣Of 2�~k�R��<�P9y��ё�	A>I�4W+��gy�ݟ�߁ƙ����� J	���yhK�- ��u#K~>�D���R�L��������S��f )�y* ��"����Ui�׾��;��=�ߜq�����ԍ�5� ��A&�� ��+"��`<�0J�'��Q."\��� ���GD��v�{*��Q�=֠Q0J3O�k�8�co��9FS>j���A�[Z�v��� H2�
���g����Q�	�������6�k�"l����WF��8�Z<�Z�y�E�Ւ��ξ<������P��V�@������x|p#?���q��[�yAA�(���A�뚃�J}�-���0��|m�8�@����o�(�iV3������Ւ��$���!$�XvRPV��w�e�GV���$3�����}�m2��K�T����jɴ�@�zƀpin�f!J�ZHjw8��@��0���~;�u�3��ŧ��gd��ٽi%��[-�E�n�{P��[Q���,��m����}��!A3��7p�^����������Կ��S��jק9���7�ͅ�G͟�k��_D���"o �l���7�>E� �7V`�Č�ZY�zj9�'㩶	� �������=���f1����=PvƲA�^�5��@�֫%�����f��"8l��J�s6��a�u7�YMƣ�	A�����r��j�z�Q?2t!�����!�r,q׽��K�h�z�4���7����R�f�Y����b-<�ЧG��@?���FL*����GDRH.�K�!���%�|g7.ѩǲ��.�u���*Ŵ��š*,�S�/�� �Л��]i`~CI�Dݹ��lx��0�4f�s��WX�a���jV�x�����u����rΓߏj���#u�:5*��yϹ�A@ .�h����q ��`|�\�jV���p�Ek��l&a3�2�<��d�T�Q���������ĪZ0�#P��ω�`��r�~�7���@]!ݟ�x�p�q��Jo*��1�ީֳ�CZp���8�{h��bW���pTY�p�Ȕ��48�/��}- }��>?�j埛��n�,w��p;a<�;Ëz���T��vai0�?���j�y�������\ǩӖ��B��*K������:S=s�k���8)&R}�)L�n3A4��M�mY��OCK��mt h��d��׫*Kh���0�K�u���i�?�Ax��gZ/;FE%�4u�ae|���_1�"%�oU5�t[A��'��d��茏j��vTynfA�����)�? ���ߍ�a�3��;��	�:Cŉ���??`�ܾ�i�L2osأ�e�2ą���R���n�G���\{oy@�`�N�JS�z���|o�����á0��B�;\����W�T��ϱ�����EF_�����e�u�����T=����Z����99�2n"�gd>>/�9C�2W���ތ/��}o�X��jvR*�9�����#��� &�����A����u�?�������S0�®-Ɇ��T���V��H���_F#���e(�׊�vB�
��,��X~��hsnQ��=j�"%�
	!����ǐ=��|�Jz��8��3H�qd��Ä<v��H(�N��^���Tѳob�S�gS�-��.ݰ93�b?���l�dS���bб�񌔕]�kC�,��Sn)N�^]�������&>Ѣ���n��4��F��=a�K0�"�DL��\'B�.�^mS{�����ZsOM���wlk���C�a�
��Ł�bE�g����iB�x�2����9�w��,�>׵"�2q@�~-��{	�|�1c���>�����S�~����a5K�О����l�*K:\4��s	CҷN��he��pv��.F rNbx�& �L�S��BŤ46��[o[�� �-3ft� ���	�Fh�o*�g�u�{�s�:&/#�M�m����S����U�S���X�^e{��(L|��
���د����j��i���)�:����L�K�X��:����;J�L���4��]�<[�u�qe���Xk�ͨvz�d��gT�k%x��o��=3n�UC%�{�	���H��m�[��WM#KGF
)99Su��O�z�3�QZj�R-/.;v[Ҵa�6��o�e����F���6z=�k�F=C�6�7d�_r��!�fYQ�4�Liﲿ�<`!Zw]����@t�[�T���D}���QV�1w�s)G��T0A^��c��?t�v	$��x[��ƨ]7�b�ɖ�}&����(T�|���2(��	�CC�/�B�������y�����_�^�5�d�����2HB2k�9�ܶ*=T��؂L|Q/tV����H�9�b��-\�8����|-�'������}D��3�x�j�����8y��q���)3��y�C�	╢*�b�^���%��*9Nu�w���>�ԉ��a,�X�}c�o��IE���i�������-����'<b�Ԕg�6=ĵY�e����@��@���'h�ew��x+{�q-h:�LSK����q�	�:�!{���@篍����� ��;f9I�<���}PMR�p� P�	u)螔Jú� ��Gʧ��䘼���|����eu}��T%8�γ��0W�����t�Wh6�h:O���^�M!1�?���{�������Y�+Ѕ������au:�/%&B�ҬWMg�	��=�q5ٓm�i�Я����dRo�������^ �V��|�݄�#�;�`eoy9�+C*H�k���<(3*'<7�1k_��i�*f�EEP2Z����r�F-t����j�+A�ٰ �������w�BaŶIW���6���.b��`�Ď�i�E�,Yg�D$g�@�!%��ϥ�����GK�c)��G�)�+l��#�^R|��O���X]�C����z�8��6�A������F���n�bӇ�"k[=�*�s��2`ԒG��ba-u��t1��^�_M��P�\��s�t�t�ʐ+��Q�RoQ���eA�觐�R9���W0�f��W��!)����QI�]�$��7��+�Zn��F �Dr0v��y���DzL�tS��nۼ��L�����z���/�fL���zi����֏%&F�at��ఫ�N1��2�0�>+q3�0��X�q�&�1�:$��N��ט@����F�#ߠ�Y]۝0a���d���m�Q�ifD2�I� ,ԀW��9/*J��Ƀt�+Ev���D�)����6_�wv�m���=��C�j�I�!��B�
��ӎ>�s�֑�~k�Qʙ���-3Ȳ�aTg��@v͐�����D���S>N�/�����}������:�w��\L����[��ז�sZA�&l�K4�r�N]	c��dVZ����V2I�v����
�#D\��c(Q%��B�4.|����U�'�X����H_�W?��O��m߄4�w<eA�^�K�icȺtp��]���U�u�e��l�*v���)��[E�����H=�,�Z����K�\���C�vK�r�ݜ%��-�F|5`�ݬ!.�P?��:��E�����\���۴�}ȧ������?Dl��b� �%�u��F�t�g�P����3�7�Rt��.�e����K�V�e��@���ó*�m�Hkm������ܱE�����c��c��r|��F{!s�֙��i���qQWp�pk������]�Wd���Cj� "?���I�8/x����V���o�
�[ �au[��5}$�ʰ�E��i�����EM�B��dS�VE֒@��M��4�$��aX�_�v}#�2H|=�
Z't�ܜ�V?+!E'r<4����ll=s�짲"����53�������0��Ü��,u�=¡�̠����	^|�`d��Á�`K�������Al6TA�25��	�jm����A}h��_�g��.M���m���jfh3�v��v�� #���9l*�v��V��_��J�N�� �u��\�i�������kV�t9�"[f�x!%)=���L��0`��[Q����n�5��wޣv�Y��WySi������Ap�����D�%ë��p��Ϧ�!@����Ys�v(S�6���q4��������6a0_���$+���V[�./(�Y]�
�� �.�uhls�@kS'�)�(]�|���V�c�����������؋�(w�Lo�;��̇���r{c�&-j+������k�����E,P�lcgv��k{���r�&X@�Q��T%�#4+������uݸ�*�#c�x��1B5?���i���|�
����yɠjɍ�;g��i���NU�����Q��;Ӻ 4�C�r��n%I���B9�ƚ'�$���-�1g
g�
*A>fl�}�d���r��A`b�]��'�2z��M�塍��
�|X�u��`1 ���=���H"@lXw�Fp���wD�)��2���Ρ���/��E21�l��"?�Y�8�⃅SN8T����	����v���]�\H"�D����"3�v} ����*���o�u�괓[� 	�����_�2B�C<]!j�1_�)�8��|,��T�#��t�f�Z���c�5c�f�'���[�Zp7��$��W^kt��I:KZ�f�o<=)+��$��I��A(_oԠm!�Q�H�a�\�Ԏ����5PJ������2�j�^u�Ks<�j����4�<@0$P���ōhц�Z1W�RBS��S����b��+�(o;z��+��tQ��h=��[e�;��\|�g8+f���ǶP�<���*nhZas���'CG�o����˴�24U�i��{7��-9�E��p�b��H��^H��Ђ�ϻH�xN���NJ9R�%�=УT�jy'�kqQK�(�*i�$��%��XE_>�_a���c�
������Pbu���DR�<�N����οeׄ= ��i?����e�mҸ4	$^��|E���E��1>�X`�2:��h���n��,�*���������sLӷў��nÂ��e!�	���Hv8���/�&���qxFm5��e��Z��3GP�ϸ�~�)����ax"��{��-�r�^����+q����%�$M��xm��i�W�%=v ����Ps姒���?є�R��f�G2b���p�@V��(n"���z�%��w�G�%R�3 ?��8�p�l)<(P�c�j�0�VP0�@��0�u��ҷ���˿��p�(j/|�A}�Xh��P>s� �z�;8�[�5�U�u�]��r��T��ɶT[����غÆ���*�)@D3wB������̧ 8֜��l\�ש�n8{q��.2�
a�S�mU4�Eµ[��g�wg.��q�l���D�dA�lAOm}+�4�1zD�U��靪�/�w*���!�V�Q��!�I�*�����ñ����A�ʕ����:���e��y�_Y�f/y�U��BM�����5bu[c���=�y��}Z���N��U�G���V�nuw<S��=�Z}��� b���1�'umy��9��m@H�����j���9�c�{Xޟ������k���͏�M�JnYf�0��v���r%(?��J��� 7�r+���H��6~���=�t�W�&�2��ȟZ��P���v�B�\!$�w�!�J������	����Smgt&q0&�<y��7/���s�S��2��(�_;Jx8�W��!�c}�J"ZE]�t2��X��f�p	�p��S�����`N�̀�Z�OJl��ҵ��QF��>�y��+�\8x�F���P���c��I�KaZ8���M7��7��u�Q������B.���R+�y-縰�#$���&�I��A5��;Tw�#�Sy����o��Q� �[�{)�(���_O�܌�?<W��v��
����"2�X��-[��Ɛ�L�����d��ׄ�� ��D�U0���?�W0�`X�k�/-���Z�$�V�ρ�܀	�hB*�']raj(*5����?Btr�T��0e>ᗑ�*��)�2��P��)�K�M4�I���I��H��U��;��)��i	16��)�<T�ś�f�V2@�@��5 @�s��s�������H�y�� a?��eXj�9�,�g���!#�>��\^���,�|o�]���5��Z��ߊ�����4c6��N3@B��i�����}B�R��O6^ߚ_Y�����J/�0����"Ć3��J�z���_@��U�Es�x�zl�@�R�4뎃Y+���QL�7i
_�,�C�@����c�����.6�oC�&lS�lm#�K�w�3�9��(�η��3��fWI$��
��G�p���f�fj��W�k�jA`Q���)�4G���˯�ި���?,��/���+�a���u�U*=���?l��~Ȑ��y>?wB��c@xH��m��H6�G��>�o�`����	5�rG:� bu�0�3G+�wx����V�����|������@�Yd!d	�.3��=lg4�<�pxw�MQˈ9����w�x�W�>���Rqp����h����5�{~��"5e��i�&#�3�߿&�����J��~y��[mMw�QrQD��cz\~ژ��^���z�P�!�D
Ta�mf�+v��)�5�� �<|G�l�1����k0�G(;�*@\� ���K���'QQ��yf���"��k��#0�\R\�Nn��?�X�`��
P�m�'����:b�ߣGY�c �r0����ZR����S���-{��ԩ�W��{dc�	w�l�.W;iܰu���(1�R����Þ���c�;6K5���q�����h<�oO7�����XЀH�޽
�l�����T�Lk>� �[�cHS���+�٧�P}=�����4��x���:x�c��B�f1�A^��ݖ�7�YSt������l1����P���|r	�2�+9��sό���Q�Ǉ��m���P~���>��ȼ_�qqf��~_&�Q�K��C3���n���v�(����_�zWoVa��!��/�����gN�V���.j��qUi�v��1��瑵�>`m��9PaS
g���±'̴��F}MCo�����sG'd<�_<������5�va(<�A�'a�~�U�q�ڔ�zxL=��/�|�K���a}���.ʟ;qu?����b�7��;jr�fd���:@�v�	Уt�l���y s�b�$|��^,�.��Z�u'���RX��q��M�)���%K��.9�6�^ f�̜d�j 콄Vz��@XƏ�W�R�Ç/��:��S�6�6��}mZ�_٬���������󛝈��,9*�R�K%;���׸���W��>� ME8�ν�)?�q|%���Y�b�e��[�Z7��'�t5�tG�%w*���T��4��[�fߟ�O���LV0�A��<xq|#ŴW0넸�}����6 ]̛����-ʱ�v��V��'_�Ac�K=�h��
X���-���K�)�x������#�s	y.��@FV����P���Hߦ���oTF�.�E��E����&$=��q���[F��^/�z�a��}���TA[�x��t"4ϣ�Dc�j��@�}��E/]c��#E��rG5���E��×���&P��Is,��V�}y=P���D���M�I�`�Q6�$�; p'�Z\�1)�I��>5]�t�9��%y�*أ�n��~�h�����Ic����P�^�����̍eL�ƱL	(�\�β�@Ķ`T��WKo#|Җ�o�ǎ,G�����_��׸��0)������88�� A�/�tï{Y\S�,}-������i��]#�+1����>����*��eN��rO�q8d�����x�j�s�ʥ�M�R�8�A��=2���a`���*�i'Ë(�W�(`�����R9/U7� @_Cw��.F�Ȱ������I'���Z)�e\��!l����5�* NK�x��L�#��ݑ!�!��K���//�0����jY���`(�!��I��j�����[U���H
�L_���
&��v���j�,���K��Z�}(��g�$�V�����c>�r:6<�Ɂ{�3;s �e�O��a�|�q|+Y�F�Vp����+��`�P/��Ә+���m���ó�[�0|��%�Q���88�A�%t^!s~��ĈH��Q��{,#[� �6�ab���R������ԟ��4I��P�H�pn��E��rk+��IY?|O�&F������?�T��}x6П�~�n�b"v��^pV4�y��ׄ���+�'��'ezf�!��z��)�Ŧ2��9����ϏVˍ�2������b���[D@8%"_�,;�8�����gF�E��b IGa��4�����_��CmX#e��ހ8{M���υ�s	Vpk�Hd3�oT�|_����������&��=�G��L#oA���m�CU�")t=9��df� &�>D&��^���]�
�^����83 ,k�L�s���?u:3S�-����(�ߑa�n8�4�\-�^ο9�y
* ܕ�@�}�C��o*�Xp{\>��Ϻ��#�6��L���p߂Ig���9&e���~`���N�Ռns4�X�)�����VJ��3%��#<�V���T����~۝�#�F_� 2CUN�f�e"~����F�+u"mD��Me�Ѕ����k5��b��=����fQ��7&�gVИކ��e�-��}k�@{���pd�N��\�#��p{-��T����R��(��=�mn��kӸ�ty��3�D�/�*6/�z�P�\�'$ߦ���OGT8�c��Hr��Eo�A��E�^blX�C2)������
�A��O�~�Ч������L@F ���gFu3���H�X�-T�ц۪B^>�2��A��1[����+X9���2��-��F�Q ���@UF+˿�IK��'3Ew,4�U:�#|�C�����2��C�_¬'������qf:L��].>R\2���;p��%���mT�ѥ���I���X������.xȏ@@���OT�����-���e{"P�sX���O�"���D��z�3�+v�<j��}��v]��>UN�EdHq������Ҧ������ǥgN�3v�S;&n�":�����Ȋ�G�+�Z.�k.j5��}����.۽Y�pO�*Z�@���+�N_؊�.�����9PZ�"�)@�3�pAV�ѯ߸��s�|�CD���.k��CE����91�:�p[���@;_.ʻ�|�:q����C�<�O#Zʣ�g��!�:ٝq�6�F0�}r�gny��ݞ>Q�Ǡ���/3_���(9�,���y��^̍I�0k�U��7F�O��!ǖ_(9��	�r�IU��-H��ڈ��	����SО1h��4��J%**1����B��cȡ����-&���;����< ����p���������|(����l֕¬�GZ8�v��+��}��ԖK��P�4w�&��kݓ��ǆI����t��*[.��\p	���W�k����8U<������f��5�=�!�fȤ��bE~i�>����ؘiD]pBL��R���D#�������`��4�U�K5��-Iķ��O?���f�+�����k��&�e!��;he�(ٙ���P3%�7ǲ'_���8�w�i�%w"�v+C�*=&�k�N-yjz/��`�jHɳ��M�0/ �%��R�(���A�����:�|D~2ö��Gz���yT� ����/�9;6.F"��+k���1��v4��
�k�^��
�X���$��U�����&�mgӹF�����3gs�+<)�,��EN_�V�ɷ8%k{:q8��;��8�6��=/�$wV�՝�hC�;����TD�Pzrۋ��l��!h�މ��k§�;����,�1�6��?��Ó�I̚��-{��������/sa��/:Qg����s�������BA�q@���Mg��/�� *[�F��MP9���Ѩ��"@�#r'����,y�H����<ꘆ�l�ՙNz����v�e{L?�ɢ��<Q[��!_��b2Nc���a/ �Y��ti���NZ�Psv���|����5��}����סp��#�R�Je�pn��M0pPi�DH��
� �QzN���>������a]����Х�p��C&,c),�9-ƛ�R����r�a�z�AA�ӡ�����ӫr���8[��0(`d��7��q`n-�l��eC�Q_��������s��.W�3�2�ڷ�%��'>| �;��Wf���;��C �/�.��Av׫���=(I�rk�%��7�H��� �(���'[[�]{�}�>7�evd:�&!�2<�ۖ��~��*��|WR	o���d�h?M���W
�Y��;� �8�,���^#�~��<?�@�Y���$���(�"8grwE��d	�p��D�1�D!�w�El ���VQ���I=52��X�����:Lj�Y*�5;�M�ܧ��o*���=T?�K���Ո�.�ܘs��kt����t$� �P�]
�"W�����t�Ψ4= �1b=�}�.0U"*w�5��-�GB����`�	|񅸔��P�B�(vX:M�� @�-�˱�\!w���N��R��.g��(�-%�)4�0�����B���@����"&U7�b%@������O#R/=����`����r�VK�o��W4�)>h�J0jI[VG~��JuR�p��=���I���E[n��&�B�u=(E�&V"��H�6�4��~����{�V0c��G�l�6��j� �ИC�7e~�ȏg8K��+�|n؃���m�4Gs�����q�>���2�����m�8 E���_j꼾��*�g����d�d��7���/�L�B�[B	*���E���.ͨ� #���pA>p!7�\�}�Co�ԯ��n��,��+�R
&�֖,K����;�ɼ2u�1��J���;��C��BZ�^�L�ҸR�P�W�@�[|�Ys�=�����3�.�ⵜaR�����CGѧn3�ˮhE<D���QZ}^���j�Œ^���~�v"PKԳ݊v��\t8���)�xǙ�θmؗ�"d�g�u�Ҵ���# ����Ԁ��Eo�\���K�boq��,'̥�Ld����p�x�:B9�&��}��22�x t F�KD�`�$.�^��<WӇ����t��  z|���z���tr��[F�i�'���:X�:�X�[�^��	V��+/F�8QPZ����\�j��O�o�o����#��(
>+4�,\˥���&l�׉2�$5�oi�h˺�@�_yhayR�
҂�
�x���Z���f�F�QHT_l�#��POY{�4��ms<Y�&�H�R5�^&�A�Ѕt�%����P��a�X����J:�L�[�>G]�[�W4�ND�=�oʋ������)�ͻV;��O���@likIb3����y�O�B��1��fpw$5�=�s�;N��4��B��1�.�M(+�y�R;
�6�F'*VA �l"B���1xF�z�O��>b��6�3M����#�,zĳ_�d>Df�ۅ!N�Y�kO��Qj΀A��^)W{���H�ǝȸA���@����������(I;��(S]�Y�U��S����i5^Jwf".��΋���O��*Ȋ��������p#ދ�h��~��^�F����]��5�����"/>���6� B/���B�Y}�&�ϗG�M���+Qp@�d$�v81\��ϳ��V��?NW?���X4��7E����K �m��=��w^��L��|�m^�d�_�M�uJ ���
ps�0G�RK��<����=?�I��rB�Khҡ"���<�]��N�9�������cU�Wx%�=��6^�'.���:��wZ�,�/��4��2I���M�#�L�)�[Ok����D� ��&W�7�Y�+d�仙U��m�hVu�f(>��|�J���x\�lJM>�c�=p������Y,�ϋZl�o��ػG��� ����BA<}��!!W�8���V����ĪM�ۣ7e�vn�UAE1�gxt��j�Lp�X43<�O�d����京v���D�H���˘��b5�Lj��b�73;�3u!���t��5q� ��p�"KWw[�FEx�V?�� ��ʬ@��wY�R6�6���n������ҩ��=�f�-���J�����TlP/L\��S���å����JڂE�;�n�-�/�
��x,�37_r���7)y����p\�d�Ԯ>�њ�f)`�0�����7>��M`�گ��rz$�������Tw�d�¬�p�����Y['+��+5��:�s�P�~ā�a���hI8� ��(a�ۡ�*��
��|\���>���L�'U��ӈ�v�@��E���E�����Qp�v�[-��t}4QN6v1\�Xw��	�ez%�?��)��"�Q�����t	u�%��w���۰6�J8Ox�-.��w��9�{Z#x��BMH\�I�Z�}�e7ߥT�ؒk��k~�
ĸJ�Q�(�X&<-��!��O擗 ����}���(.��=�+7�?@ QP����zLzr4טy4�����㯀�;0i�!4 8�j�VѾ�N���D��c���]��GJ�SI��s7�i,���TQd�*f���[��¦�rÿ�x	�1�i�_c�F*r��it�D��c��p���պ�:�HW��-��V�)��ѿg���:mJЭr�F��X9���8���68�n��C����K��*2�B_��l��ޥ��~������hO�w�p���ƌ7j��N�N�m����m��ڕ���4��7�^�j�.U���n��1�]f �]U�g;����h^�s��F\�ՠPZ�3<���.�<� �6��aF������^��׎�e���6B��6~3X�`}&�̍����C���]""���>�U�>�4�����󡖲���p�����r��p��?�9Kn�����FXcI���h�>]������n����a$���Y"`G��?�`�˳�g��Ǣ�/�]Q�AӊC�����s?�P��޹���V�k˯a��&K�c���sRc��W�������N�l�s�9H8�F͵'��e�-^���#��*NQ6
|z��Sy9�|,��t���(�AkT���,�hVRm�?�mzP7����;A|�`��QJWU�*oR�_I�2QD8���z������9JK?h?���E:+�i%9$�?gy	�a)�騯�v����>Zz�A�\_�h��	�mŪNoG�O�0��h�O��qr�?�J�k�Jm�Y��kܗ�Ȑ�i��LV�6_�95�t��R����<��?�D|��g�sQ�f����vʩ5�d����**r)p���D(��Y������~�桵I���L���ԦY�������%s�Ym#@Q�`م ��Y�C=YNk�&S!�#	�
^�Aw�|� ���x��]�=�8��9��{��k����d�$ڳ�R����ْj����!\�3���<��l//�e
�}{�&�zܲ9(�7Tb�� 9	� 5kQ��Gz�f��<�4j���(���m��&�s�م�N��&��מ�(�\}z���< t�3�W4qvT$U���C|�d�� "����&��@q&�Nw���.I��Y�$�p�~�L����ы'N�1�8�>�p9�,?�ȶ-V)X�c�����;��UZ�;�
������>���V.��1Ǥ�
��R�9ߥ�F���&k}YA�&Ңa���#w?Bf~8��P��y�(��Ի[�ݜ�k �&q\~�"���Y`5s}��p�u?���$M��gT4�K	��';��*�!C�����K\b
��'�"��"{ܨ���PRذ�x��������_&n����g��X�M�:(�z�0 P� u%��(��C|�܀�$��+�# C]p�����Kr�ņ�� ����
�OY�@���9����w��<i�p�}3�_�3׆Ok��=�*1����(���}3�j�)G� <r9�e
�A��ҭn
��h�!K�� 3l%/7�2,��f�T�󦷭'(�֟ �~ү5L�\��d���@1������v�p2�Ǧ-�=�;^%�JUD" ��?�n☇3K�)��ՂڥF���&�=���et9ۏ�R}�%�k�R��=���_�a��K��b_%�:ۙ�Ah���#���^��.*��@*wA�8ƌ��1�TA+=������!IG�!�x�E3�tc��2�w"�j��t����hv ��M��.�x�������۪�c��K[b��ޙA��+���v]�j�P�F���[
�������-�8H����ׇG�U�y"��E��ĹM5������b6m�|z��P���P�� �)��?BI��>���Q���b�uOtlc��N���=�������5w���P�qM|.̉��=����l���ʶ�Ӓ��{z��5�3{��_����>:�=T��������3G)�m�'4�RΫ��Za������n�sT���H��KCU�qĈ�1r=eLsw>Uȫmȓ�Y����X���s�c�Z�p���`����')��^�&ɞ5���夒4C'�ݶiQFpfi���&2�G �P��4�^�ݚ	)T�C��̗���Z�ze��i�F#k��d��t�&!{,����;��@�L��PS��`���hM2v%,�o�y�BNRn>~8�=�u�4��%if�}(��1��Q´ޙ�.�(�չ9���w���E>ߌ=��#a��%����r�����Vv��T��5~L�-BTҴ��w�6rq�鳊X���"��뙨<ie�;iO܊�2�[�-ro����:b�ץP�h�z��-��L����׊�~!�J[r@D+E��IB���U�\WI���s��ɼ�Q�g_����:Fj�W�fF�C��7r����}!.�G��`\�x��>K�la��M�����B���U �/L�	���\)I��`)mb���Stu�inH��ݶ�B&����?e[�Z��z@�8*�j V4�F�q����i��-����TocE�
�N�`kH����J�U�vxt6l�p��n��W�)bM�]�FU�v�>mr8h�֠E�SCFkI�k��A�<\�o��L�&nR:]�f$�{��$��B"�l���u'g����[�(U�{�-̞};@B%������͵�k=?���W����E����P�z5lR��U�߄�y=Ѣ��	��>~���)\��_0�bB�r�ż��tW��A�˓�jz��V7࿸_M>�,�9����PӇ�SV~+5���6�׵r�OՑUv�&(���>�n�]�� /y|5��<�kz���w��ۜ?HJ��Qg)ס��|+��+*��m�O�8(���~��k���4��=l�^�������3 ���.�`�d}黖~d�a���Ѯ?�ۥ�L�� ct�O��=�ޡ�3�v�+���"'��J��	��Bj�� $�6�U�bw(�<���܄��X�G��7�c��{�)��XjHP�zՎ��U�qo��8���C��Zf����NӸ��#"�wІ�5��)!�S�r�ȧ~J��BPW�H%�.�^�#J��e�N`a�yA�9��PoR�?�F#r�B��8�M��~��/��|�O/OO#_0I�����{�8hHma�#b��kOH)�����&q�S��N���/}������m!�����]�4���7�hN;�G~����?~(�l�6��|�W�z�Uj�����Uo�<�t	|{�	:O��9҉&��Qs�����.�u���}돠+_�В��ֹ�k�}��{Ӟ�A�>߁�C�DH�2ֽ�IV,���V�D����+OZ|V�<���xV/�Hu��Y�{i{0Ww��b$��%z65�yV��
����kz���6���հl���1��6R;�Ƌ���Կ��;}^��"="��_XD-?Ǩ0�ڃ_.5%&�>r��B�iQh^1:��4���̘�#U�$e��%!�Ič���)��M�eX�(�#6�.�D�@+�I��l�?����Y�utc��v��\����*�SZ(��lYH: �A�m9`�Y�϶�ڴ�6���r`l*	 �f:ʢz��:2���{d�G�tC>u2g�9��15ᚾp�R?{�t�)
�5�m����l���_l5RV�i�4��H����į���vI4�?���-G���dz����2æa�N��\є�n�C "3��#BsMh��J+�m���:d�c�+T��Ȑ�Jv�����L�|��͡�) �m?�����sS��ז�j�1���Q�(b:P��4~�
^�
�/YƸڻ��@ᦎ�KHH֡�^���;˝��QN�mԤ3�*
A�0a�Ap�D��r슓�tHl�5�rY��r���aq���#$���T���=����������K��&q,WۗQ�X���<�<N%�ϔ5�����v}������F=@L���h����ΐP5��	��e�H1�aJ�ߵ�}N>dbSֵ�]�a�UP��"6��V�=���X���O*h�E�W�:P�əs�h=4�����(C�� l�����ƫ����>�e~�'��#���Ε��E琙�89����x8~-D,��.7U"q��o'V�� ��a��'�W��;�%�8����H���|���`��������̢G�w?Ϧt��x]� r���2\o�.�G����j�b�2��N��_�����ޓ�aH�b�P7� ������>
fz iۃb!������ �ѪS�h��c�ԮԜ+<�,�C9�,�4~��(���F?�&?�!�K��:(s���Y������ fdw ��N	��k0xQ�֘�'��ϋ��asl"�w�LқƺI�M��G�2
븆����2���(�h�ז�R0�%��Ӧ���4=�ށ�T,�2Ώ�	�P���Q�A�N>�y}�k��辵8�����߉4����S��
������xCʬ�4|�6�0t�c�n�����ݜ`�A��m	�1#J�S'hӱ���ʻH�Pt��4�CT���^U���`��R�C�uc�V�?7W:����A!�j�n�O�
n"D/ ڬ��s��;�� ,UEyB��?��{^s$mH�i�dg$������������-��է�:-�&���_ƪ�\k�:,�z���7E��st��[��T�U�ͮ�p}�yB%8;����r";Y�@�-��A�|�B.�H�����i{���H�B;�@�M�vK��xf��X�����pe �}��3!ߕ����yT�������q1�>�e��L`'Ǻ����z;��ځ-�b��¯�3j|���dk��6|1���At�B�{���E}Kc�'6�ϦO����֗_9gO��	w��M�t���jG*9,���gO��+M5�>��S# ?Wh~��[� ���J�<1ÆjW���K���J��/�1���jTO�Ud�-]36�ł{�k���k	� �M�(���L�����������ʏ�s��o fD�h�o�!�ɿp����=�=o`�<;8��@X��"cH,]z\��Pr�.=XPS���7�	��TDMTҁ��HP�h
����"�*�[;��|���$��.�PC
P�����X)���B�e4¹��!��|�V�g%���馟D��mV*р��{|�&�S�v=d����Sǜ�RF$y:���bd��O%'�� ����a���*�u�����������]؞PDy3�Qvm�d�(�W��&O�_={��,�#��覬=�͈�¶+)d^��Bn�e(��c��H��x�AƏ�=���EE���ƨ�!s�����b�A������;9��B�e����,��4�Il�T�*5�ao���H��� �`�HzT8��q$�t])�mf�o.�s�,�����!���B�2 ���qVnϡ���%��?6���u���ZI�{��|S�-T@@�)���%���c���s�ؕ�H�Ă�-P�T�x�	�}�Q�
|�p�#�*�L�`����/�A���H�}GL&ՂK+�+���S�b���)�r�o٥���+Yk��Yc}� �C�*(B��f�h6^%A.����}s��)�/��,�CMU��I�-C�E�UzdN�;���%|�AT��|a��	��­�I��C�tb��|j��T%�FZ6��$��4�����B_�-���p[��ߍ��$&�/�� a7�76���2>���O�X+�VKl����Vk���(&LN�Et�����7�E�'����ψK1���bHj�A�L�}��<�F_���b*���!}@������Ӽ=G��1�
[3Z�O\x�C串�^c�C�A���w`8+�]�iUgN�6�9�#����vDr�߃��+Y~�@2�ڍ�T�
�;\_�[ �FB�i�1aS=�9��a�"NTj�X����+�D:��xܽZ-Q �)���~�]�C�ܝo��[��\�6�4��Cl̃����Ud�8���_������5>jաU�zQO=����"_��7p��������Ŏ��=�x��|>�6������!�����i����I����k������7��5���ä�J���U}D�;@-|i��E_�1X�H�Q����$!"��d�$��0$�����%�JL���t�p�O������)�o>v��o�D%����(C��O4��A�m #��
�������CX<�h���c&�!l?DI���!t��=���g��u�jY��_U���xV��>��b�@�>�
f�������X<;2��K�RDu�<y�������Q�{?{ѓ�d��R�KGwE��g����7���#r^_�ǵU!��i���f2Ύڿ�ע��uq�k]���9��_�y2�v����t=�E.�ޅ�_�	Æ�hq��%�%�%pW�Ru؇j����=;�1�o�o�p�Eҩo�����/��PO���(��5`�be�	u��@(��-�+���GJ˱����l�JuY�e�����F���lᆿ"��]|1�t��uB��ל^Ϟ�b��`��bwCs�!��K��O2��u{$� �E���pR�U��0)x�b��'|m�RU}�̩�ڥ�][���d��:'�a�+���������]���B�
��o��r�@˖�SİMNf�$�y�u<(�%gq.�*c�bڦ�g?3xs
�wum���g!#�`������-�o2t�������!�4`I��ʘ����䗀ډ{��%ͺ�E���c�Z����r��_fA##K}:rl��Мo��e�Z�d�b4��!� ZO���F�S�ygH��-gi�݆�[���$���Vc�MLu����)y�����%�e�z���aN�St(~F��7�nG�S�����Z�������Ƨ�H���p]�Նh��}����R@,o��G�	���{``R���̯��I�3��@A���3c�e�@&�*�g{Y��G��N�5���v(HTzxZb8��<I��댩c�_yJR385Q�]���tn,�L�B����'���\�!6f����FH<+���qW�3>�eÝ�s4�ޡ���tiP�g��QRG���YA����q�h6�
�N*���-+@H�����qZm0?����������W�[_2Ǉ��,��.��s�1�0r��Faiw�����q��I�� uɞf6 ip<^@Z�FS��"��V���{5/�22��/�-x ���!Xw�������b�.2�L�Q�d����''c�|x�Uj�c��hy7F���kt<��-���	�j\�٤��X�g��l�n���_��z̽��c�.��k������V�I���j���+z,:��,�JD�k���-�l>!:���Y�dĺ�a �^���	�� Ց�������"�����%�ꖕ�?8|~s���fJqG�_�h��w4�1��?C�w���W����F��,��*���� y�6�}�n��쾪�m@�0C1WIH.0���=Ś�*2[��ʨ�"^�͝��l���Ce����-�A�l˳SA;�{(�=5��_��O퐘���P\`�q�����A��ϲI$�Gue�ɥ6�@�'�97u+6BI2�4���_�eY6^ ���ЧBw6}���] ��B�h��'
0d�". G<�&	ױ�SF�n���
�
����k���zc�t-c��K�W�h0�Ł1���RY��QM�x�2̕��}Av"HN����i���@A�_Y��q�e�?Uj��,�W���*^�@�53�ԑ&a6��1�j:Hx�����L�
z-�! �r���c儼\����2 A�Nf���N���cj6O>���J~N9G+���;��Nښ�T�|�'��)�Aq� t�� �����h��%�êE�d�o�7ޕ�N��V��"9���������WXDk}9�"AWC`jx��`S�cՃ��VWpd��xvR�ّ��
b��C߂��J�]��g�jL��`/�,¥��A!�_�r\����LL5����M�0Y5v;�@f��ˍ���o'`n�ċ�"��l��FD>����yg���&[��"��s�!�Ԇo�?���5��7�Y���~�Zu"X���r-m�r&8<�S�҅�iq�Aj��9�3�� ��d&�O61�K_��8�@2:��=�����+7["nU�~t�A�6�9Nn�l]uR�z��AU&S_+����.$'�����n~�;Ȩ%Jg���X���|+(����F�XE���oz�Ƙ�;o�a�
x�ŉ�Z
�K�m��ჿ��a>p�'�]�GhU�H����1Z�^����0��KkI�m�S(o����� v��A�����a$��J��i͗�>�.W�5~Qs� ��&}')�Օ�1K4����*�ŀ�\�Az�p��}�����G�K�_��Dv9r"Q�#?!Kc�p3�w��R�a�[��!$V�KA٪���;�B����T:�����Vw��YjX]g}�àa�D^(WcI��mɤ.�S~��� �+}(YE�3[f��,�d��^l��FE�0 ��5U�'i2W��P�:�_Ӛ�eP��cAlD@�U�;\�G��?�fU�j]��2�ߺǋ�����O��{���vs�1��*�q0Y'ՓY�]�� i��,Hin���x':uL-!{��N���tSl`�u�ջ�����W��\j@vn��0��J�̫]�ɐ����o/�0&PM�]U�#d�I�;W��t4�������ڎ238��PQ�Q姎����o�����{o�3&X�{�}^����zDh-�S�����X�:Mz�؀	.k�IT"�0�Ư�r0�]��lڪv!\Y�l�z���|W�������$�a�=A�'�&�P�&����9*�0,���G��Gz\��.��n �Q�t��(�<R�����w�� #p�D�i�8^+�N�#�į��+��a������(�*G��ty�u�!�0�l�R[�#����mz�~��X����촇�Lol�7��}�� �A���5���	N^S^ʇ�u�J!��jg ۋ��қ�B��6�c��R(w��T*S����^�N���Q�����D.����ga�F��a���x(�A�O��(\1\Bp"�cE��<;G�B��i!m�BX3����vixk��ҟR�H.�j$��_�����<���H[��P�/�w�Oi&$#Ah'���pY������,��IR�N�e�v���f@��6M�����K���,��T��mR!��-�5��Bv�4�``ϛq�Cb��A�F¯[Z�;�[�!ZD9N�-�k:�D	)���/�V��N��ꍞ�4�(���˭�L�!��E��Å���11!=���V�X�n�:�4þ$��8ޣ�̳����ͼ���W�R���a�gf�aI�z��{M#�\�_��>%�Nߒ5ʛ�;ـ��לgt0vl�(b�EY�D�jܽ��qY�*ָO�p��%!��[�3�@�n��"ց�Sg��ծ�Z��m��������4$G��1��m}CzI��8{5Щ��'��	�t���?sBЋ��b=�u8<�A!�B���"��j�+�<��Jo��NYgI�֋N߫����hQ��.�rF�N`p���p��W3w�ǸzC�U C�6��8?��6Ү�������^o���Ɛ����[����T+�i���:��ڄ���� �%�j��j�雖�U�ܣ?90��|H�������h��o����+TX	?^N R����o\j��mV�o��cǽ:a�0ut�A���������8��J�횏9��J���GQT,
Өo�a�&��+��nU���:�R]P�~��6���oM�s������'vqʙ�P�s����^��bz��Wu�(�����S�OD�� (��y��~�ng��w>��M��6��EI��S"fs%�(ҏ�o]�=�=�����y�����Ⳓ�c<S��-��³6v�*%U��]��-��_�:�G�����7���#���@Ψ�%��
����������٣�E�R�#cA�4�*H�E����X���_9^��/����N�it]��N+Av���Z	1��6�Q=���	�]P�Р^Nm2�]1
��^��x�:��!]�C�_c98���,4�/g�5�GA���E��N� ��F��S�2+NP����}=�@���܅�>����{�����������{�p#n����i+����΅�X)2hX/}��0��"dӄ/�&��k!��锟`�m0�}��y("C�c[�y��w��R���ߎP�a�Q֫���ݚ�wFHϑV��K�>���T�-�R�Ȍ�q'	I#��D�e�lw�)]��`�����T�pm�B��#XZ�E���P"j�vR�u��i��ߗ�ݫL�ѻ�����3�0��`�F(��r_6�&SL�>TWNF�#y�%�S�����jZ�Is��eͤ& c�Ū0և��0c;e���Rku�`�x�����G�M ��K��#��V���2�N�f61�ӊ@��ۢzO�/[�/�3ck�?|�v��aJq���tkYRyp��!�֪�!���/�CER�5!�����6[�N p�Pi���'[Q
�Eu�YAL'}�5Ͻ�¿��ܧ޼_�ҟ}7��cȽC��k��@�A���?&��󈗼��&����7݇�;���h˪n�K��X�0����h�b�|�p��C��02���tq��0H��K����l.�8�s�YQy�V9�Ny�'V��^���آ��z3�P�
��U&�-�4�6��2�"u`�MHD�)�.�aޫ��Ͼ멵�f��Wh�dR��A���r8��p1Rז|��J(M?C �(2��;��C%U�/Ku����&}�}�E��82rx��C�C 291�`��ҁ��n��-֥&V|��׋�һi	�4k��y�HA��~d��]~�%�f �A�}μzS~E�2,ɡ�Yuʯ�qL>U�����G�)9x������]�U�!eu34�HJ�ۨ����LW|�/�]�4�Ļ&bH��!R�a����`ϖɒ�Jթ�{Ke��x7_�~l�f��"C9c�}ӎ�1�k�����Jhw-(�� �%y ����s��0�mɼ�lm]j;�):�鄶<�=���MyK7�"��1;�K�Cn�4Nx=�c���&��Vp��usʯ'Lݗ�X��A���`i��?��f�S�K�����?F2�@���؟�o/�����EIo�[� �P�m����\S��CX���b�1�}���X+�4��yg5dȌ�&d�G�X��ՠc�ݙ��ĝ���јHvgo/s!�IagI��bĦ�L���I}�a�9^����ד��!᷵���]�E�+����s�q%\%��?x(׺���Jq�u�د��a�,�F*����3�ӷ��|Bò�նRc�ΖSbN�z.w�h�U<2��Bt󓇖{Bِ�'��!?p˕+S�Ԙ�Li���AD�������4�EI��.@��D��轼!��K�QV���}�*]�DM��3e	KO���w=,�N��B,"�J!�hu&�e���RIM�B~�=b�X�7zjP�(j����Z�X����x'����PÁ��}'(<"����+���z���=!�sr��,K�Ѳr�L�j]-/N�6&����Oԫ���'W�k���˩W8
*b�Y��K4%6��	��1�����em�
��b���x�Գ��Z�}*�m\��m4��׌���kAnN�x��8���?��	T�q�~��|(ę|�pw NH ��6}9<������J�2U�q���ru������~
�楄y�|��k��C�4]D���mL���FK�0�N^�VV��]�v)xk% ��D�jlg���(�PNY	#X��+��I��CHҒ����y4YH�QYgj ��t�<�蔸�$ܒ��`�/ ELxl���@��\">��Q'�g�]�2]��L'�B�z�P�����%��7o����Ch|����Zy��cDM��}�JlO�^}��@����/�K�Cn�۞j��$ tD�".����4���J-Y��(?�0�+a��A��aM5��cP@�<)ѫ&*.[���v���h�[�b����0��9����x�fcA�q6-�j���k� \�"�3Ƭ2���|��w�t�Y��+�����Y�$����&��	$O���y�p<Lq�N(��K���ػL�
6���*�Xl.!\#a��� ���o{�W�hF�Fg��L2?���P�n�,r|?+o�ϻ�Z>����u��ݱ��*��=n]��ôl��'���:�E�!*0�=�U��M��`��%�h�����|�@>��D�jᚴp���S�l.�Ƨ*��ec�|5y���Le]����&L��$�'��U&�O|
8�!�"���QZ7=^ӕr���CѿJę�l�2龿���m��V�A��5�;J�z`�͛"W�%�=�ϭL�fO��=�W���$Z$�h��S�~��|�	d�%�Q�+(��U���3,�_����`+S<�u�O��s�!2ӓ�����$��0�c_��[��/׫�;�/>��kd@��S��Q�@`L
�o��U-N]2m�xr&#�~D��p��1c7�05I)ݦn�X2�HҀQ~,A�_����L��Xَ;�B�d�RI����xI��I�:�k�
7vs�k�����}y���X/i�������s���"�&9���� �aE�R|Qyd���V���	X�S��U�F��F�����4�5��C_t��3#�v6����a�K_S�W�Ăk��~�"�$< Z��m)�K����t�����==N�ŕv
�N�LI,m��`���u8�1��hGڐL���m�5q����QIv[l�irϛ�;d�T�����;��T�4�4�9
Q���X\x!�qO���l��%i�d�_-��>S�3�@��~~O�Q|�|�v*~k~4W�� |���a������0�1vl�U�@j{��e�8S��H�v|㳜t9�e0V��!�j��f��B6��=��(:!�!����8�W�v���&H��vZ�kh`+m�򼌪y|�y����1�� 9�#C��$���x�ݭ��H&��L~*t;s5���B�3�F/����K�6+7��g��.��VjV>��pEEōM����;���jI#X�`{�_#�C2�3$[���#���4���g��`�y��E�����[��w��W``a%\��L�1H�\>GB���Y i�'�5���P�x�R��� \р8-<�4�
��ZFF����B,�[�}��wo�䜟����x!����&l���v��P�+~�k^mc��V>ݲp�ZQ��}�:���A��R<<7^�Ga9� 8���4��^7���n�1���S����%E�q]�(ez���8-�����{�x�Y"�U����)]��B�D�������4��@�'�X,(N�����:�,�Z��Kel$]&ޡ��6`Ѡw{�#�^��^D[]�ͼKɀ����Ë��8��x�j����<��i�)��lK�z��
���.��*P#X�m����B庵����{���}5�Hu�)�=�3|�	a�
�/dD��D{�)^
��<�L
Ӗ��]�p���`�LC)	Z�)��R�C��6�w�.�ύG�hE(W��/	�X44rr��U_SK�J�ޗQ���LIqQ�M�ܬ������?�	�
PI�b�<�E^Jd�E��ȿ����ѬmD��G��բ*��1#/KZ�g[��ԢJ}ՔE=M�[~A����K`�WE�֎3�PC����s�(��j
���Q�	񻬾�	��'RQ�T�7�a�fp�@�,��S��ϙk�Be�h���[��m���5
n��*�2{�%vǊE����,n��E��/7�?���r���{B�Q���|�?u�xXO�����g�EIWG��7�R�<��k�§a��A�����Y�߹6po+�Yw)����t��h��*0�]h�5Fc�+�����Ӱd)[׍X��l�5	�&�c���5�=q!mg�싊�yd�F�������3�'�CxiM�j�g2(��MN�G��l|�W[z��U�oiK���y�EN�lV�����-XL,�fV*���l���O~<:�e��>��y̥ߨ����=X8HL0�	��蠴����	�x�W趭g]�;{�iJ9&.��j��Hk�C�n1�ta:�>��iё�B{�� ŏ]L����fb�L�6�М�1^��o�f��~�H8J6<V1�Q'g��]0�{�=���-Z
����.��l�	'��o5�W�������%G9�������J03�!�j0����Nu�/Q�T�6@��������?�Q�Z+�@�:���$�C�d>NJ�f�T�ڢtnf,j΁8�<�m\Nx¬ ~����!`�,
g���"s�'�z����y�	"��«�V����R�1$B�h�T�<���u�����~D�0�"�F��;z)�tծxLlQ*��ѣ�L9+��|G���T��������-�l�������f�W�6��9&�m�{Y�<�?{q��)�kM���*��3�1��3��;��Q:oP�4QC���?�~cN�ͺ� wh�G3p��D_���
�0	UK���m��:^�� 8"��HT ��)sz�M:��|C��T����&�E�
��A�U1C�I�����z����\ %��T�����,+�X�L�a�{̙�e��9۫5߾��}V���e�7dr̐f�4��}W�WX�O��$�R�mYra�/���:X�;�ЌoB-t��L����P@��� q�+�r{y���Jxp5(�L��'�&�yL�g���ѥq��ѯ��Z���`�\��.��?]�F[�W�*2*=�ء��K~�20tW��}��	��<��2��N���>�s)��*����f�/L���ɨ�ZN8Y{q��2��B|��X*�0�W���A�4z�,�F�F��Dw;��40���nV]U�F��d�;?�6<A;̄k8y��s����*+B5�'�Ţ9�T��)�pB�����"X%sN펋��ӱ�����ܑ!��1�{/�]?��Q�e���N������Ӝ�
�<!�@��-�8	��|��]G�i�я���r�h�􉁚v�e/��ɻ�n$��M�Wt��s�^>X�[��c�4�qU6V�}N)�2]�!3{f�Kk6���]���f���E\���nW�'�L���n`1R1	Y�a���|	���"�@(�?�<�V�J2(���-��g����k��f���e���{Qe�V鰞܏�
ʘ\��%���2���B(���^@+6�Tc��PC�ٷA	�4���M��g$�����t'����h�PN��_�j��R)�B�m�Ր�F��T�-�+C�%�\���;��a�����dE��̪������w��KP+��|*���I}���g9ޔ��'T��fV����oɶ�d��m����ʚ�#l�V��+����F�I8�#��čZ0:��*��Lk4���4�J�����gM5	�e�_m��*�o�Ӭk8��f�� �ݔX�U�!�Qf��\�q�Z�29�6n��R�J�!�oe�����G�k�Ct<�;�3X����ïx���'+�)b�+�����_�Hm�5F��e�5�Y�p0$ng���-O̺GRIO��P8�z��V�y�<n^ b�R�H�2���|��
7^�Q*�%�6�Ly�*
9t �>�cf�T����a�o'�`�{�po'HSԹU�KXm1Ue4Årđ��=R���}�ѧ!3�_�S����Zb��d��Fy��YRxW[��
������k7g�2�� �%3��&r4re�f�����a9^"�t;����'߻�p
dy�9�b�s4˂P[)ULQ-e-_��>�+_��bH"�Ȓ+�ߜ�ښPěvʽ-X�L��5���݄&���K
ӊt�8J��eT�}J��Gu+�̄3_Gڼ�t��R�%~�7��g!�)[����F(6��k_�'?K��,�y/?v-R�q��T�'$EuJ��p�����Б!<RzIId�
���E�9��H���O�df��K�G���9/Zɻ��`2֛UP��?e���-c��=r�R2>�G�y���w���YI�l�HX��:o�Dy�5��k�OsT�"�E>��0zg��@r.5�w�]�uܞ�ŏP}��6�����נ�>�]?,���=�N�jp����0y`�%�Jݨ��ԧ�gRZ�z\��B�n�<������v��rK2�-:$G&{r���x���^��+�,�vXl�I�,J�z-�l�=uyލ�1�������9�(m���+e��\U�Q"��Mf��SC���hE��-�W-��H��)�;��V��j7�=��3n�t����~n��;�Jd7 �5g��'�۴3��ѕ@�K��/W��op@�
�)ŅI̬v0q
sNof����D	�������.d�ks(�!G���-�A	9G����H>�V�gB$���H7l���A�%u3)�L����1�����3�וy�|�F��I��_��D۷$�� Y����E'N�A�'�$�|�䫿"��(wNO���j@6��������.�^�S��cZ�oY����U�(ߨ�6@3ܿ%�xW��YC�y'
!�X�.`���Q�3�CĲ���Bg�e�����c�:� �$�}{�/t����&ؕ�H=orH��ZEr�������#�-���YR������H��v?�5�>�"pә,v��\7��k+�-��1�3���BI���}���e��/�����5��%�՘*�I��̩9^�?�ݶ2��j�NU��]��R?���}5\k���OƦ���I��%���ZH{�7,��TvZF�K�
�،�� �2}��u]5ۆk��RP�\ޖ�,�lPX`���P�	!C����*��܌V�e@���+=R�C�h���~b�ْ���s:@��Y�Xa��U��>�� C��O���s"}X�?�s',��#ع�rDd��C�l0�<:�'�zv��]m6��j�t.a�r��a�6�%�:7c�{}n_��2����FV��ܑ�&�a�(�|Î�����\1R�O�q�a������2�bb_��R~%�$�س �5�D�p���:���u5I�M�H�����@��i�/1��/M�����!�b�x��v2�g�(��	�};��Bl�m�4K.cZ*�NBɯ�=X�Q_�� 	N��ȆpL���V49��!hz�`|��nw�����>d���A�����)��E5^�^RB5�������h
��:�%0����k'�Ш|�#�P:�(h�E����k��P�H�n7��d�$#�{�,sv ��KT��������!n���	��s����C��)�����B��ȗ>�Wo2x����n7c`�d�7o �Aԏ��ڰY��v	�y!VkT�O��%���v?Ը��Xi_�U��rC��앁�#ӿ>�D��M��e(l��6r�+q;_��G��N+��1h�Vr��Ĭ~"����P�0H<�CA���x�����6c86�e/o�^M�.�0p7hpH󻟯�%$U.�
$�����ۚ�����)�XZ}�zA�T�����^B^S�3�--�8Ѵ�s�\F��C����7�/�?,و-2Q�,J^���'e#���F��E%V�6J�m�d':.mV����Iɳ����՗bNF�1��/��}���ĶUD��v0~%S��+�����8ȌĊ�m��w�� ��֕�Gm/sp�E�]d���<����u�PN����o�#H����]j��{lq��)D].��
<쿝�د6<�Ѽ�γ���_,��4?W蝜m�	;e��
�ݨ_�! Y8�ioW�P�q����F ��!ҩ�D��8=
��`�e�ͤ��}F/h`��F�O�l����K�:�挎$��c7�8�8ulY�b��dgp�D%e~3�(���0uu��݂�/�=R��->�)��Q4�j��W=N�f����%9,�- ����P��r/�ᨰ���<Ɩ����=�D"�6W���J��e�53�N�C�E6�~�Eb��G��I�T^xֺ+�M�fZ!�v��z5?���}�o�vP��^�N���FU��3�6<�sy�AY9��;ܴ�7�I�y˞cg��gk�5�*T;��Ly�� -_��z��5�Y>�0~8�6�����2@N�q����=�oZ=n�4G6i�uv7�Y=k7�v�T���)��$`qQ
{�O��&󓗁-Akᨈ¹;��Wr�Q�$0����_>J��>�TG��z*bLL�>�5Z7%��B�HO-Y����arB$��H�I��+�_Ν����Tq�����ȩ?��jQ ��e�����)�.�C��{l�7��!(��{ޅ���S4�Խ�_�l°�j3�j5�Fo����@���՛�@�ء�I�e��]UPǙ�-,�E���ݳH�n�-��!!��q�uG:�N����~֛�w�v7a�B��=ޅ���EY�96	�Ƈ�{!5қ�@@D�:��m�g���B�0�v4�)������ ���x��7��&x}�� �uMؓ�����*}lw2C��NN�!��b�ƀ\��� �>�B�j�U�θX�+A��z�T��q�_M3oU�����Wr�5U+!�'�����&��j�ͷLkG3�fR��"X���VI�I�@����$)d =f���zQ�����4��k�./��E��J<L#����w��ށ�O�D�|���V���B�4�	ˌ��Ȍ&���T�ޖ�;>k��N�{DR���q`I���Y�}����>+���%?o~3���"x0bk�W�D*��8��7��`��l�I�w����|�1x�Son�������6D�4�G���A!�`������ N�kķ��Y�?�2���CXKW��x7Bp�L��+0��ͥY	����e����&���,�\=s�r�iO� d���d�|�R]_v}UH���%�l�X@���<D葚[���z"�C��s��)Cs�t�.'U*m}T��d��s]\.�r�a ���v
�t�7�$kh)���8�t=��9r��p�Cr�k��K1�_C][���Wi�N%'��L2`Π��V�Jq6�o�](�5��մM���vI���7J1dݮ4M@�QYe��0�LƔ�#��#yV@��3;/�׺QAS�������w�Đ��Ƥ&DZ��*��8�����cp\ߦQ�I2�d϶v�x�^X�'|�Z���.�e�G���\)�au�|+�i��X�[��튤杉�ޥ�hv�Йsbu5��|P\�v�����хui&�_"Z)��T`w������GO��z�S�s1�*P�;!#��9`nY���8�L�3�a�v��������X)����p���>!��T��U�;�Ⱦ��-.l��zJ�zA�Ʋ�^��C`Ä��'��0���?,q�7��zA�s�9ss��`X,P���Z��� �-oRޯ��}D�|�2~֘��W9	/��&��dT*�����C\�'�x�p�.�RЀ[i����M�L��憪S�iw��;�ǔ�G����g�W�I��B���2p$�B&$��&������0�*L�',{�
Z�ƚ"T�	@J.�7m&2��GJ^�`;����_�^iR����!@®ې��$<����r������Kϓ�|��s����&y ~���id���Ah��Q����
��vR����M�$f�n.Sp�^G#`Yr9��!�*�o��	Y��>�A��S"(����%���)�g�C��q�],��1���ܓ�FY%o�x�`\�[5�@񂤜��Q��Y�&Q� Ɏw�<�[&�{�������vy�G��뒷�(G��6�	AjR�x֕��l�0B�L�z�e��d�fQ���o�,��ɹϞh�7�l�7����8zp�+x;+�-ǚ�`�d�Yzo�:��?�ƀ��?s~��N�Y�O��g���I����q�Jʧ�!BM���	��1��iQ3�@X�35�]�Š�y��w%�'u��h��}絜_$V���Q�[]"^�f�G�q�wq~.qT��?a��3 CC��A0�s�_.�ket�z*�]ew6(��m�mŘ���`��P�NJ1R�֡��-��g�����Ż �W;�v"F�q�|
Xioaykծ���[��(��8������|���Ϗ��g7��S��M"��a��уߤ�yW���Q�~��j3?������
ivb��sV��)��J�ؚ��"Q� <[����XT�̙�u���VC����CEފ��h��׊����d$~9+V5��XWQ��T�0�#�P��K��;�.^|�eg�H>D����?���м(�^����9`[tt��&Ċ`���ӝ��F3�g�1U9b�|��ӌż]b�����?儮k���a	���������}���y�� �L��b;Y�Ă�v��D{<�)���&Ae.�y8�ǔn$�K&U��o�\�AL%��Bf~�[����a3&P��Wd���<�~lr���}�/�k�N�(\d_S.'MnN�}���쎺��B�m�L�׬��U4 F;���氹�%#���!���
�+|��q�3*�e�g�����6XQ�r���^_��o��Ai��xU!�&Z_��F���?�؊���^�yhTR�cK��<F��O��	�W�ǃ��� �Ɩn��OfH��_��a����L�[�fkJ���\�+4�Mq�Ӆ�c��+`7�/5�Gdj�K����b����sj�)Ҩ_J�1,]��}��/.̓K�G�:ԣ�9n'-u:e�������#�Bu��7��[GFƛ�
#Nh��!�X{�gy��r�.�%���<toɥ�4t�])��v��}(�y(���=�z��W@ϯ��pQ�����]��u������(Y��Չgj�V$J���@��č14,8����Ew��ò�.D�u��Ä��3�[>��7���U쭊N(��V�b�5Q��/�;�T��fh�	�<�o�/
=>_�(���E!���IoL)�I|��M�5@����Tꔿ�E~*���� ��$3���M�-M�����7����	8_;�����C:��3�7�"ݲL�O7K,�ܲ�k`�_��U��t���Yݖ�5"����\=�cRv(O����Uyv�� �u���`�����Bu�Y�}A#
r�줄��\�7�D�\�"nF�J��'!�w%�Rj3��u��� ��-]�Z��%�D�}�{.o�b:��9N�hI�,(�,xՑw�~G����]bQ��xͻ����]��Cе�>�G_�	b�֗�l�B�.��x��/�ߐ�Gx"Ź���`�!h�����+T��������p0(.�}ǔ6fƒ���HdI'����� ��6N��� �R��G��w� gT ��H��|���A����<�Nd�ų�:Z�[��k�|�-��@;&-��7�����nh�����HG*wT�J�������M�$�.�h�Gb	�D�9#�A��Sv�	��(��BM��u��w`�28�X�<5�����L��+���: Cadq��l�!��"�L)E)�|��˜N:�Qz[N� $A�@i��b��9Jg�Yz1�#��b�g%X������4V�Q$�+����d(`i�I��Io憩�E^�f�P�	o�@,������7Ԩ�L���̊��8�G�WU�-s7�\�1+'h������ �|)�"����;Ũ��b%R�l	Y��f�t0�������)H��"BM��XeM�b��-�!��4����S���s��{y�k�����%����M0��H
Qq�n��J�ZZER���1<�:���o�S�e�(O��Xʇ�ߠ�P�Y�i1ӛ�imH! ��u�\��ݕ���}D̲��a��W(��h�����k��'[��Z[�2N�b��͎_r�Ʀ�V;�i�:Z�F`��	d��`@���ߌaJcL0y����ɠ�䈤U��4X�c����5��lm�4�]�~8�5�#�+�X���/����ku��ߵ>˄���1X�",�Zhn|��?�QM�}; hW笟|��:�ӼޔKcU���qPc�j��}�w8���D�GA)��5_9Nv����_:*�Λ�O��/%��D��'��7-�����QF�W��wF�.T��\~1�� \k�u������Mp� .)����,��Ʃ�'9$����-�bU�����[s�8���y�&���/�u��m�׵q#����G)�E��܀d�m*' � K�%�^;�ՋBhl�&�	��]p��صk�X��hQ��Bw�P팟������2[75�/h�S���w�s���`�6V�5��=�7��G�*����g��0��%�����h����8&�!'Bӧ_�`W�!��:M_	�M�ʜ�1���q��N��P(�϶��r�_� Z�0�p?-�P�숪���I��%Y�uAs��R-=�}�1'Ң�?�����^vu�0y1鄧faBR�7e�(���r_m��B�a�F�_��h1t!�$��3Ȁ�[@�������8�nO/4*�?.�P!TtCWyԸ��^��"Sm��X�f-C�)����X��+��e�.�D�K�=K���Z��s  ɥ�k���f�+i��X#[�4Z�w�$mz������)�c��ΡC���Z��As^�f�����S���7�C4��ŵI�FT�� 4H�TB+��?�����ClAًZ+�KY�yL/�%���ײC��>����q�Bn��K-�F&��*�����D�^�,N+U�,C���ڣ�#�#u��p�����l��j�`;�I5xи)X�G���N�-�t&��Ub�"sYK`%V�Z�=!����{X|%{�ʻ
po'�6��-9b��S�f
�`��؟���䄲�'�&-�����,Ģ�+����X?��ۚ�*���0�%?��i��?�,u���� ��O��
&NC��0�TȌ!��܆"+��I[i�\PLա�>Obtf�����`?�u�DhF�wu�C�����<���WF���qj���lR�����هf�F�"g��8PAw����,,a��Td澐@iAMլw�W�z�@��S�<�uiVϪ
��f9%T�̽�r�h)�y�z�[9,��yM	Nj^>�u��8Y,m�1tV�{�'h�`�kٍ��l4-T�
Z�G;E�T���ᆸt�wA��9i拼��qD�>���x�,3�h	H�"�Nm�������2�|"s�����9�Z{�}t��y��Q��V�8������=u��ݍ�d� ���ڢ��C(蜷=J�N�n�O����3��tmǉ6�9����`�Rk�0fY�.C�ͥ}�̬�d�=���9��1��M��CeM�/�-����V�R��<do��E�w���S�m���G.�Wc�oGˑq�����x��*|���ų�B��X2�fO����2K�%
�=����G����<�+ܗ}\u�V�����+�����s��#��˱n��o�Շ4�/��1N�%��V��\��MA[_����[lr���+fŜ�u��bN	�c�p�1�
���K�YVûx�)��.Ub;۠�֪�'�����&��]A���߼���"��d��SY�����C�x�g!�SS"�tXŰ��D�U]��o���ˑҬp��a$�#/-�};{��Ĵ
h:��1�5{���Iz�#�̏3h�#4�
������Ms[�)ղm=�>���x���#�EX�v3	�S �[Y�(i��1;*eH����w �U��m`�u���i��(]���ѓ���,E��t/:)����k��ó/Sw����f� [ Im,��1�}��_� %�_"��}OSsv��?�D͢��&��v }$�\�[lk0�'o��5���˞�g���1�6z�oTY�3[n�N���&Hf������F������&^���xG�01��X��X ��/�2���r���0����,���<��� �����'�����y��T!%ow����Կk�͈��?3�LO�0����%�ILڅ�&4"�,��~=�����Yvy
�
�%�/���=��si�pj��b�|���W+o{y*G�,��������a�������$�����5�T�5����3�[��Z�^�ַ�Z���0|-�3WwY�nh'M|�|��.��n�hB5����'
�Q[��].&:螺	�*��ʂ�ҥ�d�{1^������{ր�{h6��d�0kO@r6#�F�k����U����f�F��^��?��'��0_ L�x��c�ی!�I�_<f��[�C���!��Ǖ�����$68ƈ 9K�����f�?��9�o:����.LF�4)��l��s�Ɯ��"�{+Λ�p��� �`�~%���8,��G��Wx���r���{w~�1gr'|�^�l/(9ѣ�-}��r�']�������}���L .F����.��N��m�埯u�f�s�����E����/��)�Р�9�&������c�S�W{6]2������cAЫEa/�PߕP���Mމ��Mp��zlt�gP7������P����]F詩?�7�]Y����Q�dL�1?�%�@�Wt�<HĠ>4a�\��o'/�n�Sǧ�y�I��BQ��r��א1M?����y�RenԄI���9H��I����|q�|�	�?���<B�p=�)���h��VQ�^o�B����@�m�7�w[���x�[�a�.e������U��҃���4�w��z|�m�R�VM�XI����u_����x����`�+�Z-��y�IU|*8��/�/Y�!�F��h�TM;R�%ٞi���<��h�xA^�p�J��Ӗ�c��oN���G
�Eo! �BR?�P&��}�O,!�u`X�MSV]��(�?�ເɸ
ޱ)~�F{Ժ%׉$� ��1$�+�(��X��������Ę�o m6����G L����0:QTl�R�&�s��Z-��2g�R�y���,��{1Y)��'L���u�7�[�/�P����3g\�$?�	l���A���J�hm,�L���])W$�\�bx��e�g�/
Jn{+}��U8ƺK��ɵN�O�HPW�7�b�#K�N��K3o�)���7��m�2��ļ'�!����(&���v'oH,Q�DW��ƅIv��76��
cX�A�JpoՐ�t����W/G�g��E�e���GcQ����J�|�D6���_8�FFg����F�J��J�L��E{۾l���{���k�� �����*��e$vg��:�u������5��'0Ԓ�66C�"l��R�玅ȶ]�]��7�,3���=��Ci�:���-GqI��}��U�K����5ܡ�Z����'�U"n{����*�@�@S�	�lx:��9�m�Xo�:3�ث�if̿���K���<���{?I�O�m��]��<Ó���]�b}��(6���9�����u'{D�OyA4b96����{�Fn]G[]%;�n�Ҵ)Ա���eN���5x4��l��/|*�,"ȬcK���_e$l�s�}E_Қ#:Ԛ��jnt�T��U-����@B���/���c �(��@�u8�u|6"#�e*�J�C���ۚ�q �W��t��R�?������$g,)8!�l_���(P[���Ŧ,�k�ʓD�2~#4R�4���Z]�j������]"YĮ.�uh�x<C��!�LkCiMf-�"xU^*�_�a�_�2O����m����� ��mG\��Wqk��制B��ʌ8�G���7\��k� E�%DP������6j[&D�7��5l���F�P�K�&��-%�Q���M��D4������%��S��M���1�������՜��T=���M�����銐ٜHM���EK��c=�(I�q"�P��5�r��������,qM`_͸z�2i���0��w�K�X!�W�<vt^1z+۽[5U=���2�y���3��CN[�a^m���01�&�`�;܂��GνX�ܿͮOJ��*{������'�=��tz��Za�ӄ��*�\��z�<�t�:��d��F��u�غ*�!�muϽH#��O}d	qmu�:�i�QϘk)h�]Z�c���@:&}z��0\C�ui�ᮬ���l�v�Fy��ͨ�=g�1�MtSKT,��LiA���|�4�u�[��@�i�@�0�����)4 ��5���~��]�	JɨE���غ+E���|N�2Y��2�_ *����N�֔B�_�vª�|&�;�GOŤ��6�a�����v����م����a.��~�L�g5y��f�p�Q_<m�[��D�~
�g5���]h�z��o�ӎ(�"?�Q�<���FV!�,O:��ފ"v��1i-mLZ�QO����޻eiQ�('���Uހ��}toX�؅--h���t�2&Oѣ �'���f���n�*r�b\%(N�����%Ă� 4�ҷ2R��t���R��&��39`�u1I�<a�Zo���U���Ӆ%�$�9ZQ2���x��$r�otR���^߫����o#�? ��!�@|����y�K���������xu�N�{���B��ᓪ3�[d��ܺ����� ��?�AH��8}9Fθ]OPk'�=T3<��JRaLia�`]�zm[�D�룙
�u?c⵴S��"�Cb�x�c��z+�����WkVg��Ah]��>������� �	=�N���YD�˚TGÎ�yP�F�+ς�&���G����K<���a�i���ړG��ԈL��h ��%��z�)CMx��8��T�����99ϒ|��फ़�;r1�E�o
�ƾ�`>~~*q�7_�i:K9�K��	���R[6u�oLx�]P)���#�ܶ+����P��r�!���-9F���h�Z��ӡ�]@���h�VM>�C}��M\2Ѥh䁉,�����=j���z}(�,g�����1/��zpV����F��.�I"/���O�>�RO̤�Q�y>��p&���?�R�B+
έ~�m�Ҵd����\���J��P2	�ב�}��T£���H����P�Agq��c��l"�q�*�8� b�P�Mo����?�4��IK��V�v�c�+�Y��m���QǛ%z8�CH�&{s��_�_D@{��A��^�q�K���]��bm�+�:
p�85^�\��^��X�U�4�:r�o栩ok6����F�1ò�n>�"k;�hT��J�w�>������O<�9�#��(8/+���H��<����E�9��]JJ|����p���	�IDQ(���&�s��ؽe��V֏J�n��!V.��/�qP�B@�2@���GOP�L25�[ֻ��AVȂ����b���V+j@��<�h�'����3����6�M�d焂�'�юg�L[~b1��G�Q����X��[L��v��I��0���af:+��+G_(NXM_����=w�Y�8�)j��c�_���+�յ¾��'\-8_V�-2���>��)j�Q*(S�H�Tܒ�,�S?����kZ�}�5�'n��ywk��jj�_����� �������_	'���(
(�:�Ú{��`�ZDН	�+�Jy�%\(=����Z�9�6u6>���[��БT�����g��C�=�8�;u�L�z@�_O��,c,�(��ӾÃ��S�g�:x�>*踋
;-#g@1���Q��`�C
�33CP#�b�XK��1��� ��Q�-���<("�����������UI@L_���&\�ieCV����:]��d<^�A.�mZ�u?�1L���%�LJ�Yd��&L����� �G�|���{?e��������شUb	�H�t��2F���;e�>�B��k��Z���:���!���&�WH���Y>`͎d[��Z�6�HD��JR���X�YV�#�0����&��[l�b�[�C��3�7�B��/��٦�i6�4�;����] �|#�׀4ӫ^�TS(7��&����IQԨ2�{K�M�-��Bl�/Puu�Fog��޴�ßK	�J-ݹ_�)��"����\(���hS�X��b�ec���3�����Š�G��v#gwz���wT��SV����l+;�r�g��>W�_7�կ1�����C��x,Q�'i�s|ϋ	�F�<��x��kg�yr�C�L,���ߌ�e�}g:�rV8R!.Y�����qʕ�k��Z$j��<������3#Â���&�f���
����gs{e�	�ʐ���H�慴�+�����?�Z^���K!��{���%�����Ù_�I2�p�q��c�e
@[��W/S0��)�<��J�n�C�C��/��z�85����)o��� ���?e����fKH�4.��h��)�^�����+�4&�Y�Qs�.k���	��3dK�x��Kt1.�4B�pM���\��k??nDJG��4ZA�?�K��Tm�'��:{��#�^�p?2**�X���y�yki���d�%��V�G�I9��k`ކ� #���/��K�I��+�tn�Ⱆ�=p����NOiW��]Z
b�bH�b͌5(0��P,Z�k��R~=x~q�C�J��t:0P'��VqS����c�{���R)��Nш�*"�I�,t�4�;wߕ������1�N) 2�S�(�'��WE�p�*Vc�5=�$�S�B}ʀ�hb��u�� 	�-�'B��W�� :�q��]�,�Kg
���.�;�^s�]����	_V�u<�5!�9�Z��~e�۬<uu�*�!�i�F����� _,���<�3�ý���{��*m|?]2��# �(i���o�y5z�@q�(���o[į	vR�F��;�u���y��t`V��n�_a�ү'{�d&SFW�'�q>Y��y��09&'�<X%dI.�:z��9V��Pa누u�`���%�(^��5 jރ�+��M��o ]$����������Z��A�SM5�����ӟ����('f���qMC�"�$�=q�S�A�[Q�=��Q�Ԁr#�Hr`C��+XF��b1��c�1eE>����ם�YY��KtDX�Nbvl9}�t��Ф����Wͫ����a^���M�9+����(��9�ZG&����M͍Y��'�z�5���E��`�?��C�|Bd���W���Ϊ��Y��T����o�^��ʙ�i��l�hg�7,�����W���������4 �m�Wg/BΠ�*�:!
���dɣ _��S<���v7~���2�!�i.7\�qtB��FH1��q;m���$��������x��}_���U�\˷ �����;�Yse,�6,�{�k�L�co?�:)/��r��D|�	<wx�B"��X�e���C�/O�p�5HFܸ�]9ơj�Q3+�,b��� �Z��L�d�h���)�H�6��'�#��(�ї��$�B�an7ѣ�*���3�x&�A���Zu#�{���=%lx��;���
�0]�XQ-, ��_Ԅ�=Ah�3Dl��c�_���A&4��Kh&,��zey��1��%�%Ԓ���z%�?�L1�Li��
�|cx���C��>�$�P��?o�# �V����$"Q����q�w�&�ع��L3�1�D v�@�l��|U~���dÆf�ýgP�1�	2߿e ��f�R'��YE6
���[)����]����Ԑ?���NN-}CV�%��'�B��7����sN|$ �E�˳zƸga�N�=IB12��Cߺ\�h�88kҐ\ƥ #�>�jF�y&U�ޟwI&F���W{�̯�#��ۦ-}����cD�P����):[ͬ�w��:�8�Q�s���v;8CR�#����l�~sےŽ��C���.��ďGP�:屴�+ۅ���X�A���c�� 
?�(��ɲ�,P��J�`eK�t��iT����Ӥ�f�}���8~P�:E�iT
K�Q4�5b�/H�A�v[��������3���{8��W<�E��`/׺�Q�3�p��� �1�P2�B�z/���u�S�C��L3�y��o���,MDYaV����o��8�u�>��!��^�R�y���)t)�NM�ɣ��uu✻d���J^	n��f]�]�.K�"�s��A�����;ݰ��rr�Ӵ�_���K^+��M�&4gN���No����� �����z�,�y|�����x�`���J��8A���ṴP��2l��9��3�6�N�F�>�h��f������ϯ6iU}B��.����*��POb1�4w㷒�I�z��.��}`��%�#P|��V栎��&3e�tO�jh�/|qZŧ�7�`�33s�5ʟ=m�Y��Tp�ST���?T�V��~� @2DתE��#���h`��Y���M�/��	+��{�0�`�_yP��>� �X���O�ua$a�Q_��G ,��E�#�� 3%xt!�r ��l� q�I�dWN|!!��S�]�sJZz}J�a�"���Ս�p����oA��Q2+�G4��ü��TP
��Qɤ�� �TW�6~��lj����V��a���f&&Q���v�-�4�G$��o���|	vF�N�m�<F*T�yh�Y�0��fN_ v�6X��?{�k�C���Z�
�'���x��<�Tk�g�	S�i"2��,5`��f&�O��zj���y�u�6������U�:��-qҾ=���������]�Ê�Gg02u3T�KF���\�ȼ��U�<(�"˻�ƞ�@����[�2xv�hG����P��t��W/�<�����g`����
��4�Z��������������;܅* ��/�~1�+FaC��3+���/`ΰ� P�r4 �M����)�j���D���Ҧ�]����C��L���n[�<"���J=�ؘ9{\W] B��*76�]��\���]���
���}�Tݩ��
s��飏廔`o2RXG	�M~'�G������U�J�@ɨ�kf`�B� �1�y:"��}�(�[}�D�tZuT~�/ʺA�z���{.�R�V#��AVy�l�"�S�6����@�CE����a.Ȑj��ʵ{.�N��}Ah�~߻wV�8�%�֦�^8PX�1��H�#M"l��N��_ϱ"p��s�C�U�2I�E�1;���}�R<:������.Y����ۖ�`�d���8LyG)�J��bLob�K*�`:�c��C+s�d����Փ��H��>�'e4.��\1��$W�s� tp�DP×�T���<� -=^�):�T�0�Oo�N�뜈�V���@�~�\t:iV�a9�Qb
��c��
v�������wf1�t��E��^~�/�j
�[�:˒�+�uvc��Q�k�j��B:L!�,F�6��*.n.�c?>-�����'��ӄkX�����a�!�1\[-�O��M+�������&�X_h�Je��i�l�f�Ʃa�� 搵I�[��N)^d�'�\�kVD���!Ҁ�I)n[��1:0�ew� ���qb��{��i����bo�PC���X���K9�"LT�����#HefP�fjt��x=U�����哹ّyVk0��vT)Q���B�yN�5h��R[HF��ͨk.iH�6�]07����׹���{4U�o��O�[y��E ���I3�1��A�������ž�#$Dm\��-��_�`pk ���-Ϩ��?w���C��2G�!u���${&v'z����1�5��M�a4r��F�Ʃ`���e9&�P.~]�iuX��,��G'I~��m�Q�@��"���KJہH=�u����)��6���'�o�1w(���x�ᶖpgm��#�H0�����Y���g�(
w:�;�k�^ �@�ZC��xΛ�\ʠ ��/c���.^GO�Q�5����q���$l1��|���L>b���
t�n�2e?e�hC"aVf]Cp�Y���,]6��7;M"�ݯ�(ׁ̽�s3,c�� ��m]V��\�l�2�;�L��æ�
��%HsF� 4=fl��ԇ�\�Yp>�	bx��0��r��~���5��]Vz�R�H.q�=QL�s��#;G���Qf*�Xn��S`��X���?�{�{�� ��\9 9gTؓ���_c��Gh_�М �yp�zu�Vnh���^	r�����R&����	�ر\nEUC�nd5�n��]��'ɽk[�)j��78�UE��P������Bw��c		����o\y�E�T����⠚��&]������"�:U��~;Ɂ((�F�٣ˌ����h��!������q�ꋆ����B�:��%�Tŭ�Z@ :�l �5�`03��3|-x �_@q���_��Z폋\b�{Ҙ���a+�-P��8���]fP�V'�>��(]��[�8����;�'I@��
v�(��,��1+�{ # �=d�ev�tyg����Ľ�¾.����	x��FRS�9-�7��;��d��}�MĚ*��6D�T_���R�']�������n2`|#�̑(��o�� nA�tS;o,��V��EoK�Y�h�$t�M�>ӯ~�(��3'����M��E�C��^�����<��@t,ȱ+����3X0��x��&k˻7�`��wL�,�y,H���,vyMDs��x������.����j1+��/L�cg��-Ӝ
I�9��WI3z�&q�����1�V�P�G)?g�!�%>B�F���n��D��ȍ*����6�����0�aT� ��_㱸�(j�1�ؘ��R�"�$�HI���k�ck����X�uvU|�h���3�����}�b�
�&ɪ?�!��Bb��>�~��͢J�3To��~�m�C	9:��v-��i��B8��а.�rw%M{w��F�H)Q�M�g�rA�G�ݣ'�#�(��I�O��Ⱥ�0x.���
�Р�U�
�����F��U|ח}�L{�ɽ)��lem3�ѩ��u6KJA/	߅��:���G'kk_�)�J��Y�(O\J�G4���`X,�ꍚx�ߙ���/�}P��
��^镘d&�f&���-V����hO����x�$�;�t)�8��)�"�0��¹b!����nh@MJ`D�=Q5~Ѥ�^?�&�伧1��&�� 	��ٮ?.�+��6��Wp��A�{@o��?3������z����r]������E��xf���wg�H�慧�� ��q՛r�A�AIG!��+؛��b�3��Ty��2&�������k^A]������F�;�ݸ��})��"��P�N*~۲����}*��>N�}�4^)o�ow'v�ڍ~uJ�2@�yx��~�Ϡ��Jx��ƅ�(�ŊS��R]c��_&�l�Gh^r�G�0G����d��th<��se��rJ��h�վՐ�7`���THt�!���t�����{�еoֱ���b���uH�6�/����8�	,���!�lO����d�����̑�P��C��{��M[�g�C@�`���\�/'z ��P�o��F����$�uGOl���sB�h�'R��9ۅ4�j ~J<�~�2b��.9�*��!��I��J������^�J�x�|	"���j#�}��@�ئ�Oj�.�H*�����.,��;��4��z�y(?\J75�r{4�c��QO�w��B� ^�����q<ĩ��X�R��
k�a�A�^�;1j��E�ʛY1V���,a����ܑ�Y�F�EZ���`4(e_�z�s����Uq�U#�ս=T'v���j`�� �t�,�")-�"�3h4�6�&;�E>-���S�F+ �"dI���� )!��MR�I����+�/ZFi��7�{Wћ�N-�y���t�����D-E�n���z}`��f֭����&�b�k��	�;�r��!�huU�JTF%��ݹ��l�|��/|��T�qV��Y��2ؾ��#�h ��,��\��ݦ�ó�&�t�g�f�4AT����s��V��d����"Qu��߂���I��26%�ԻoR��A�	�*�05!,���ߟ����C|�m�����,*\����c�m�H݃���.7V����/�j����^��j�l>���ֈ@��d�OhC��e��c�t�: _����.aY6�n�\���v�M`8��+𡋭���n�91��'���6�6���f�q]e�ZW�h����/��y�$_B����e�ށ�ohߘ�T�2�H�{�j���e-,���l��n�Z�֑�'��Mu�u�Y�� V`w�rRm����Ipշ���D�dvL.�]13����S�����o�q����f��FI}$j�
���>,�w�����[��k�/�N��US����Sw+��L�a	ҏ�aJ:�n�����ݧ����:�=���I�!�չ�<�4p�}/���\�� �;�Fﶵ����ܬW�gTZ`�*�\/-Y�XnQ<j$�{��!9���55��W�#yVVu�3������x�Mme{�<���>_�d���ʾ2M?��7�?^!�F�O	PO��r�A��� #?�ិ�[�$�'�z
���Se�s*W�p9��+r�:ǣ��̷h��-+{�|L�-H�v�ˣ�La�Qěs������I<��a��ʜ�����s�C�rI�VPGo����xq�F͸=Wg�bA�<xEP�P��ف�	�Ĉ/�5౥�j��O+�6�L��@�ܖ|���i��'�Pϫk������S����.�P'����m;ᜒ��Xq���j�̫ځ��4s�,Q�O4�����-�I%�1c�3%kU�&z���%�aП����K��6];=��Խ^&�U�zy�H%Y3GoV�![Y` �x���v^lQO�_�����51�FF�pK�U-o��cߜͺs,!���^6��
q�ƞ��
{��ё󠻧���`�M�}ξ�OK��8	��	��X��{Hąs�-��K���m,x�ݓ����+s�DZ�U.U�X�/�m��g$��a�O�O����/PX�Oۀ�m
mԥ%� _Ɋ���Z�W�%��d6��Ox��C��6�K[,1d�W:p4'��z���u����2clnE����g���	=�Q�&$��E��bk�D{��;���})�u����xQL�}��n��1��O�y	V���/��s��_y�U����Fa#�D��l��IGV4\ԑU%N�W0��Ή4��l&�� �&")6�	��5�;]�q��YN��H�O��\����_W]�6�Г�Iҵ͏§	���0��M�aq�n���l�U���S���G��D�7��g$k�
ߘ�54�x����X�1Svt<���
�I/�o�Z�!(��db�����������S�-��R�L�E�:a������:?�2镕�)56f@�C��^�+���3�QK�|��E��y<e�4�1�?Dc\2�R�L���+���5�o��bM���|���7#��$硻GŴx� ���a��'q^~NX�[l��ͭ�f�SVz>��Z.��E�G˒���l��A��~@�[�#����)�s�ܐ���gv��`�S��4:B��ףw�W��DC��t�/�Q�8f�)����J�ph�E+�}��C5R�t�5�TZ�J,h�"g��*Ўz�u�履�ɰ9|ǀ��I�i�j����1�(�WC�l]�����*�Q��T.^���+�*At>H��챁�E����Y3�.�eX=eq!̳:�y笲|AX�]��S�B�vQ_#��$�݈a!(�
z�4D����� �4׵K�Z슈3T9ڴu��S�.��b�S�Q�s����_C��%�`���#���;��B@�'IiY����)F�2H�H|X�f6�q�_�=:�KV\�I�? E�)����b�#�4��_TOh����8Q����H���o��i��O�����k�91��I70�dG��1R:Wz�-\U!�W.�c�qJl�(�?�0�>�&�f�4-=S�nN�D�t▗��|n-� �d���iE��6�lDx����B�v�`,��{,����;�Q �D��О�U�v9�b3}A��I)d܃�ǎR��E!���� #��!�ʰb�!���v��D�����r�X-��{o�gjJ��װx����DD���(/8|��:E�)�g���4�i ���M5��9HQ�����҃�j�7�7&!��?��6�e��W:�}"P�`۱Ɍ�����k��z�Oӝ�{���4�"s�⎷&��F��t� ;wۙ��1J�G����PB����`px
�E�C�K[��a���N� � M��c���?_j/��Se�y��>#<�2#;�iӰJ�tm&p�y��fc�8�ؔʟ-���+��}[�3bL�*:M���:o3�U�|e�D�����,�N_^��l�NMO]��~u|�Zd�]'�A��W6������=T6����67q��V�j��D2���k!�6OƘ�m��^@,�K�l/6X��P�����͐E��?��nEj�xX@7A���_ [��N�����%|�1:��3�g������	�\p��ݑ�$#^5]:�/���^W��ٖp�'B&�i�k�U%d�͑�%ל)�Z�gx�ZeE�6��Y�(e�<,C^�O��1N�c���n'z���H�Qj߀��Nq[ܮ�]�hb9�b-|])|�΍B���JI���j��wS����A;�wms-DH�`/�����,����h��/���#���'jJ���8ƍŵ�&ݣg��@��?��k&����W��P;EXo3Ȧz� 1r������M�/�em)k1��1ʪ��S��by����`��K\��g�>�7G�.�F0&.k���F�om�.�Ě��͠�Q����n�=���	��(��⸞~K�>���qfG��3��2�j��4�u;�P�P^�?nI<ő�VPj���b��r�����^q���I����yŦu�(`R��x�a\�C�q���W]�ߤ��Uh���<ݴ$H�ӥ !_#��$s�8���P�~�sU �i�bI��+��k�/�oe�^���G#sy,�:�yҰx�C7IKhb�1��J�F0��O�z�,�{H|�zS���k��p�b�?&�4�`��U`�V*\����L����u��3�7�b��Ol�u2r�4��s��J����{`��*G��6�e��2z��CO^����.���ԑ�]?�������eOh��E���U�R�n�����V����)�B��Ն��Z���C!0/\R��4P�i8�R����h�-w���=o�)�;y�yj�<Y;���>���YKI��s?����̵�Xǀ<�V\����FJ���|���9h�_�\3g�ǳ�&��7��E��r���󩬀_�{�>Z��&8�m>��2B���U�rY��Y풱�I�	=��F�n���a�O-W���(���[w�2�l��9�䬑�͕J��	�tZ����������f9�p��U�u�2��Nl����sdk���gKP�M5
ՠ�����T^��{��\x� �ùf�0G��2�z�UJe�d�q�>���_2-�aT;8᣾Q��p�x7n�Ԉ�W�գ�Q�+Gk%X��Y�8�Y��g`Jz���t��z���Z����>ݯ���I�jCJl���[��N��'5�k�k��㍢�J
�i��i��FP֖�!2ݱ�"C�]qg_29h��;��9|O|��&b�X��Aq�`�3��֍.�;����H7z��;N%*���Յ+��'���>�&��Ry�EqTN�ݫzIc]�bX������8�ҞL,-B�Nǋly�.����C���u��$��W쭗�l,Y
PT+�>����6,�����C���ư������_��o�������� ��则��bw��@�%��E�O�閃4�_`�g�'�Z���#�&̾������?p9���Zf����u�.������'*��84���n��wY"3٧���|E��F�Pj�'�'����qB�pH�{;s��W�\S��!
��ǡ��1������q�ϋ�^N���V`�3� �%�ٿ�@m(��9���x�?�#ڛ$��W!�vA��l&�=�߹��O��8�kG�UB�K�gZL���ÑTm��I��$�_���&F����L���s�TA��C/�����������HQ@�ǈ@>�˙
K��l�L�aP�Is�r��ÿ;����M�\�ɶ\C�.�_��8����&N��i�P�ymklvQ�$vG�� �]3�B�(�BB;�M�Z�������������!�XK�ޜ��N[҉t��#��<��m�����`)�$OsS;��H�Ьx�:�`V�@��pْS�P:�o2�)���~6�5��?���\_1�*\P��8��ئ�d�������(�G��1�Y�LG �x�IbS}�;��������d��{c�DXkn�'��e�y~�.���7�B�j��T@j�[W�z��,焰��{�MV��ˣg��/������/-��ug>^�*��5�l�)/;��*�DG�Y�:g�G5%�.�����8왘�A�/8���ul�p����Oq����3��$̘Ԯ���y����3���/n��r�3��WO�w�W�r�(h8W�Rܺ��,Y~�Q�J�C���I�-"�b}���n(e�l���,_x�{�>m1��[>ԿxߢWy���ރ@��J�.�x�N$��)��{���c���q>p��w?�oQb/8�|�d��(~X�@�CI`R��զ	��g�	��Cp�t�������QpK��$J	����w��2�2��7��0����<`�RT��{�<�g��%ʏ4� ��6
���U�a�/�!'�51G�β^��.����!ML�H�xI�%�%R̅�b4D=J�U-W`�ɞ]py4 ڸ���T���u�u-3��	D"�0�����i�h�P~d�;<�`�����Y���4��H�_)��l�B�S�o|��"-��Mi�v��?��@�Γ�Y���W�r+�QRӐ����p�@)@�mv�)`�g�fOW!"	�0���9]�%i��d^�S�KR�UFg��#v/s��wQ=��/��9	Û��U�Jr�a�T2����$�.=��uΞ�'�	�0��v����B3C�K���ʗב�7c�����G�ӌA0�ʬ�n����a/s,�Q��d"�x ��9�e��� �v��g$]1h���K��>��:;�*JKC5���"g�ࠖ7DD@�:�k7Q�~�AE���&�vD�aƵx:�nUi�H�fR�2�S�NC81{	g~\�]�_,�7^��*s0㫪W��?�`s+1�22`FH7�����(�c�����O�e��t�Ӵ��<��fy������ wW;f��#�F���8���0R�1W�l�wD�^!,u������ͩ*�8a��k�����4��(h�ɗKQl��+�FwOZtl8�e�kث��;��Eͻ��!�eI.�p˽.�٭��� ��$u��xG�B 3�H��k�E�G� �(��v[����	�W��:8��]{��� ���x	�>�D�5�U(�&��sc�O�Il׈np��i8"ǆЫZ(�1��ȵHw�͏��)b�gg�&�W��5��U��'6��5nw0Ϛ_��2k5���,s���a֬��y�|0C�Ar���I��(�CF��t���>������3DWR�?�v���� �f[Zq�+�͡�����uj�dPs��y���\���v%Ƕ>��~�	V�o�m��d*^7�W���4g�qz`���?Rk���X���%W�s8�$���x�A�����՜9O�x�į�j�;�h�"3P��ݕw�n[�l��3EE���u���w֬��.Ҡ�D���A@�8�u��Է�k���������zI$����&��W���&$#3�Є������=�PW��T�Q����Tr�o��<^�*�T}g��}!aO�PN�St���g�v�k��f��RF�$Z?����i��Ζ���{����G�?G�i��D�X�a��fp��Rț�I�.�S�Lŋ�TޔN:�������f��)�����'�E���'m�K�ճ�>R��8�n�Vy�Ց~�X@�_�͌�Y��'�N�:�&W'u3:��Za�%Z��N�)��W�*����	j]|b��w�9a-TT��-;W�l�t��p�2Q.7��G�����IT?�g�y<������2�u���������*T��*�^ �<�>�֮���x)"d~�]��22�G3&j��G�U�_D�`�=�4��A+�M=n�
Q-�NG�ʘ^>VsW��E��|�}R��9����*"�/}*�������n$u��f�7�Ö?���824��<vs�:I3�m�-�
SL��$� ��������Q�Hu.:�:�����5nf��+20�xa�|X	r�a�X:�l�����|�U(9���h�\�`Ƴ?�Yv���D9s[#�v@��O�v��Әb�0�臎P��a�	OF��l�a��z�*�n����iB<�Mu�cz�i�<��n��ϯ�;Gq�E�x�u�zn�I;�Lg���#��;U��=f9��uqQ%j|W���G��5�%R�L�濺yY�U8<�˄3GI?]'![n)N%�5[�(�f��MG��k��5Az9'�QQd���<��ʦѮ�>�$xR���$���"��3E��܄;��_���$9�˃M%~�U�}��|%���������P̙�}ĘW�=В�u�	���3up�o�́���J)G�o�Ò�q�_��Y��΂��nv�G{���j�%�\Gm�ԨCW�&�U�6}�,��L����>3J��|8B6s#�ʠkX�K�.]uO�f�ù��]T��)�����	����N�B1/��O�X�˃�*��"�n�w���%�rЯ�����%'������i�����V-������*�.�����6cѴ�if�/?��W���6��z~�&���������[V��Uɿ���+�^�Qrd��~"��������L�M@��~$ l�2��	�v�aw/�LRr2��	<0ւV#T�7�7�}rJ��Ӽ�;`aO�٣(�ᛳG9��>ӭ=��C��R���m��P�t�/�]w��1���-�y�L٘ �������и/#�ӂ���݃CI���":�k�z��Vԇ�쒚A�0���Eg�����[�����Y�������{��
Ӆ(��E����!��h���'vdZ�k�X�������XfV?5�b���ƚ늉2��x��}�ϛ����{i�i	˦k���jt�<Yi���>Z�Ȫu�x#����^�-\S����	H��LW}�nö�ϡ����w���PzQ�VN����^Jh<&e4��w���Yڕ�iP�����ܜ5�f>����A��cB_ךm�ŋv�Ɉd1�ni)v�*]�7^G�R�T��t�9���:�LlI�=�uW^.?@R�^m��y�:E7�o�<"�к�p�un'd`e�R�f�צ���<MU���9g��!4�H�m�ԁ`��υC��y�*�v�_Cer;��|�Q(#�U5!~�xɘ�B��+V|\�@z�������y�'l8�u�%h�W�/Bi�m_�+z�@ ��)؛=dЍ]�S2*�*yU��R��~:J����,��+],!�&E&,t:ė�&gDw\�V0�r�?$�G�q��T�������zz���LCm�=�W0�T���"�NZ�g��%��U�ɤ&���0q�S���!���}��_-��'"Q����9B-��O):ay����@Q���C�ۏ��J�0�Z�������db'Q��������B��<�ύ�
U�6	�ɜ�Is�70������&8vu:5���xtJ9�u��s�'��&5s�:M��I�\�Ll�E�j� dP�GOV���O^?	�[���6D�]mEz���T#h,�\�߀�x���9��@H�cX�r��J�@]�TJ�#�<���E��EQ$��k�#�.JU��x�e�[e%��uN !#���4�2� �ɉ
X&�h❈�i��=�{��׍�!!·6\Z1�%�2ܽ��#Rv��+�B��Q���L�{	Kl�)}Ë�.=�»N�oTe>Eq[Z{V^�]��/�b�p�2o�Gr��SY&-X٣@�ѣ���:�0Dk�C�n.�������b)yi�f�5N�ӆܜ4y���Gkz����)��;��uE�u��y.y�+_�_���# à�Bn�r:u���F��e�Ĭ
�$ ���F>�����/�yzC&�˝1�|-/a�c�B}�㘲 `�9�\��� ���]Z2Z�XȂm9��Sz�����I���Q�u����7��qY����q�VD8~>��3#>�N+�)���� 9��&`�%�Ԗ������p�:M>�4,��O(��c�#o�3��$�ix��&o;�+l�Z��^�A�ք�i҈�����ƹ�zZ:�f�����$��GO�����M	�.�3�@�=���ӣ��"1�V8̕5ӑ�P�E��Cr��3:t��d�1��t�]1��T��٤�5t"ޯ6���$#� ��7Ef4]m��b#�Rd�oQP���B��0�h�Q�$�'읩s]^ԟ��y�����W7��)��ђ{Y)o�-D�	`��|��:!K��M4�k�������^����b�]�~��	[�<���h�U���!����h���4b{3BAR<b�(���_�Q�i�zAx� �tNFA��d&��TK\�#deXnj3?����*U��m����Q͍�D�3��C��R9鐓�u��m(��<7>�;?�Yc����`j �)���������3ǽm��A@~IRM.g]��>����w�1L�4�]�,�ߔ����s���_�G's\@��Ǩ"U����?]"t7�7��p��JW��C��_��tm�Z���	}���pPk:��I�V.�'ſ����	L�-�S$ ,���5C�\���,�� ���,��J4�z��"�>bqi���Z��Z�v~�	�D*r����*�D�̚$�s*��$U�d�4�oo�eUJ3�ۡ�"LCQZ��c{EZ�h蠘	,K���=B�}��N�.����|4
�}��+ l��OSN�Lۮ~�X�׶��\'�8]o�t���7R����*��9�:���WI!���R��;C����O�84���W���1b�W�(�|{�>j]��P#v���e�
{�{�	�����'�SuG��H7��N�/тr��m���C��羦T!�my��qd(k-h�O*cw
H��|�e�����Q��x�!�)�{��Y	�}%�dVr�Y�n��clO�g I{>�ɢ��0<�͂����WZn)3q=l%-$%=�r������r����wk��P����aݚ	�(X�zם�	c6a��7���2�����E?D�+��Ou�i��r����N���%�,t�ޖ����7D�BQ梍(�Zb�#�8��G����-c_޼�*��L��<��b���@j}�����ۆ�,�!WI��"���5������7�#�2�G�@"H�<�|�CX�h@�zun��.-�����FH�U!�u�'c�/mu��$�
	�1C�}�P&�:1j���	�[�B����$ݥ9w\�Hp���c�����dȧk�9M�:]��4 �P;
���pU��f�糠KI*�^h~���k�]����<"[�g!�+E�������X�|`G%�4����RN<�n��י�E9\o,s)����{��#D�r�A4�� XG�����?�=L6���eX��C�I%�#De9�Ul��C�6��������g,���P�x��.H�N�fiGP/�����q<=2��ŷ9���
�)9s������{G��G�'�Ƭz�^���Y�Ǔ��X�
���8��oa�M�J<�n��@?��}V<�aB�G��/�?�ul�r�D��zx#��G%�?��tYO�Bxm)��Ĵ��ϻbc�Q�^���g:.P�	����"�������΄@����1��HR8��z���m�����l�.�C� @�I����J�*�W���Q>�$�!Q��Our������*�V/ ē�@.������ǧ%��Q��5|��?Tw,�V��q`ժ wa�e.k��￥��@q�]��^5>AG�X�'8mC��_]��B5%Xf��J�G_����>GP��ֻ2�ucfd��펔��̃�'�hb�����^rQ�w�7� �"ϒ�N����ɉ���`����1��o���
ǒ	i�����-��)�B����h؆�2R�;e��?+]�"�G�S.t�J��έ*�!���t�7͐�'!6�-��N���*�@�5�C���V�'�S�����eސ���l�ri��n���g�O�џ�v�����������M��;H�B��b�n6��S!����'�<���LC �P�".��S(	�0~�:	��D2[k���[�?B_K,�����<���E}�w�vm���_��ɸTX��Z�ԝ��Vٱ=}J�|ћ�m��h���h����� �6F ����]bx��=9�O�Y��`{҇Ǡ�pW�)���B��2F�L�����'Ռb<������v��d0���N�u���v��$K���&v�x�Hi_�AŰ�x`;�)�=���(a��;��ŋ���j�p��+��m��t %�{�'WW���ᖂ}E`)k̉��`���CbR���{���ޱ��pM��Q�Sn	S,��PM���O��(0��f@�?f|��~�
pT�����%����:�m}�P^�ߡ|��%�^�r�l����g��>��b���6E�:or���% BIޢ������5UKւ;����<�Ѯ����SN�]�؅���FMxx�´}L��Ș�i�����I�g��69�fHײ�r��a�V�3�Iٹc�Kv��)��9��`�J����XKv�>Q�S��1U�7��U/+L�DRr���QS��Pp@�ᜄ�:�u[�g�� �� ����<Ȇ�Ƿ1�����AG�5JT��xne�Y���F����	����f|3�縓���JxVX�, �)����Vv�.sů������y;��;��M�h�I� �}f[���"+�H5��ܦ����7$NQMxf��^��tjr:+�?�*lހ�����)F���o����@����u9_��1�R[�$���f���:o��M�9��Pӗ�yeu8�GΣ@?|YM����P�����(OUr�ն�0���O���fI݇�k���{�4�C����������6HɎ ����h+��+AE��(�(S�3jۊ��}�K���ߦwWؒ-C�d��Θ�z�RD�m���Gי��n�T֜\0P~hY�c"�S������d̾���բ�r�	����4��_a������A�?("���TOHO��S�! l��̨n^�20��	NU�;P<��s�>A:\����C?�O.#��Vv`6�b$��m�b˰��4��8P����ou	]��M��fy����}�H��+a����1��'���R��%n��2���k����3Wm��e�K�5h�6G��n]3�����lҶi�+<6��ݭ��T�3�<K�u�ӌ���I?�V�q'B;[��b��g�]���D�P��`�At̸U}�S?4-/;:��I�%�#m�M���+%�Z���± 0�J�Bey^��T�ι�|�t�b�� �3T���
�/P5���� Y��<nje�=� �Y��Yk�RzlfĞ��$�^�]Ґ��?�(	��S��;����Y��&���_��2>��y��"ŌRP�쳕�'�=��DFs��b��@���.����y�%n�����d�3
yall7.JN�)��]�?��<�34B�oA��q2,�c��e�����-#�KL�e��L�_Э�5�4D�5�|At�t�e�ݠ+Zp��(5WH�l?&Wb1�\�ZQ�t����ɿcM��w��3��X4L���>�H�7���XaG��WϏ��A�ݯoO��kB5ć�:�R�U+9��nڮYg���pM��_��y죮�]��:>l���������v��w�炎�u�ҋ$�z�p$~����Ae�m�υ��BPM��N�x��Jf���J�����9R������,��� �hy23�]��0h��.
�T�&��uL�B|2�D�x"O*1����<R�#�8�X�Y��Մ ��%�ŧ�f��5f��ťr��kI���3�^pL�08�DS;��d��`��$؈���4���׶X�L��"��{�'��Fd!�W���o�#j�02���<>d������K��3w#_�$�+�L�"a=}l�[s߾�d�dWM��p��D������#u"���3iI���I�q�$NwW�υ�����`��e����5���.݌��*�%�n�S"�|���`�#��}���j�.�ґ\B�&���G)��i��>��Sf���o��6����p��*�Q� ���l^��S��Q�?��#ov��yNj(��(ks�X������ɦ�v�wC������X�Ţ��qZE�;Cx��|Eo�<�t�2JX�`�2���s����/��	���@���;�S��v���� �&ث�uFl�YN�v]�XoLbg ����������F�c�[.qSYc��kX�<�I-��=9��Vڏ��bF�^� ������;�c��y��ۏWq]�H�� ]�d�+@� }T񆘝��`���i���z}dQ�7�2���s�5�r�ᥜ�bȜg����z�X��±�0`)Ή��x߭���fZ+�Wb��F?rC�@!o�S���HV�0o�<+���$����Ѥ����E����7/����8�a@�j�t�� �Iq	�:j3��h��X���y��#r�	�{m`��%_"5mB�BW���\����O��SXza���4��Ä娥��`�qY��9�
��3�w����Ѧ��,����c�}�� ���0�yZn�[��;�N�eq���Q�Y�$����cP\.R]2`-�g������x�dD�d�8��Z�Om���M������n��y�0\�V�Q��;�:�;B���*ߍ_�!o�txgd�D�ڇ�9^F���X����t�jE�?����Ƃخ�2�n?;���<A��V�F#J�{z�t��P>���{���,6h ��j�W��� V��^��@M���泗�>����"?�Xѳ!Sh�If���N���]�j0U�cZɄ��
�"8��N?,� �9���r���n�IQk<��tLq�#�>��l�� _���e5u;�&����Ohj�h���s?a	����>���A���O5�Z��=�y�Sr!�gp�`�#,�ܲ��g$�*��7�/ �%:b�6G�#��J$$	�)�S���\(���\��LH�zH�
��7�%g��SF�=I.�zy֦�c��?�+c��~�.����O�7/46����F�Y�:IY��2'el[h�7ȷ|$�F/8��^��`�b�˂6�B�ސ�EOf�
T��܋Dq���5��>M#6�C�̅�\��xtE+~B��q0��dJE���RX�#z�.v�� s�$�#�XE�ʻp ��Q?kH�x'i=���B���?kԩ��y�&ݣe�G������
)�6G���e^��I��6K��-N(�������4��ݤ��5��ҿ��N�>���ZlGE\� *���c ���]Ny� l�hy��R*�!-��&�H��������J��)A�["z��e9U'��J'^����k��O�;��1K%]��s!�u�C��:8u��@��+j+>P�E��#4��c��*''W� ��`FڜN+�촜,�����qMCWe2�_3�F񑓁��LBuo_6}G������$7����Q�i)�P��h������%>�oΫh�I��}�P�_w��E�2�Љ��JH3�4�Z����Pl�:B~�l@�&
��HNiT�(�-�q��.�.��^�*/���BȮ(��ՈJk�^����ʭ-�� d%�����S��*r��0���
��J��W�I/e:;h\ �s
t3�*Ld���~��Љ1F]���[:ЦҦ5=*͞�Sں~�}�y�=�y)yC�N��x�A��@�c�2?���~v��q�_��~�e})浂e>]f����z.�O@D[O~m�V^D���T�L���fd���'�c1Ⱦ����Q����%E]�?'�w>�7ɤ�,~��w�*b���S�OC=�Ш��rT�othş�w�\n�T��=/��.?PlG�<N��0�K�0���g�=�=J���g�=��³#)���eg�zT�I�w��[��\�^�hK'�O*I�af��yG�י9�B�qT8Z���a��^��v�}G��A(UB�%�� �Q���.��"+��W�A���_��c�0h�奸��S�f��!m��U����v���s�����HV,����܁�S�P�'F��1߇Ԯ.l�mA��P'r�>�R�ڔ=�Q��ׅj�h�`������Fχ�F����r�{�nR�	=_Z���8r>~а�],*'	��`�ٜ�86MCYQ0g����4;mL��\[R%���$"�0����E� ��G��k��٪ı$Mg���k$\}��kŧ�%f�ݟ)G�~��˲i���HX@ӿ�}�R��"�NƬ��jfn���Nsw�&W�5��@�`+;�3y�]����;(`����Q"]2iY8$��(�pG�>D'>\�S�x����$����ඖI�T�Ǹ�<e���nO�����hω���'�1��Htv�+#���L��Es��X�hH���:&FW/�s<Þ+.?v��]%aYv�����0��_�;C�`��p$��IJ��x�ᑎ%E!w'-jEr�<��i&�Tb$����E�]7�|� ��g���+ާ�Q��>C2�3pmT)���o��6�0���_�:���~
�JF���9Id?δ}�Z�Wj�:!�S{1U��iV}���9@@�]2n�����"��u� r]�&8�E ,�/�Yjȿ��8�Fs�>���b@�C���"@lP�D{�J؎J���F϶W�9�?���Mzs�.4�p������/=�5�ک�����Cڴ��y�����@/�u�����(`��S�+���v���[�ι"�$��}�I�-L���L4�A���&4S��p>���龋l o] ���%�ۉ�D{ӈO{�<W��A|�%��Y�Vr涿�k�d�� IW���1�a+a-���a&�!�~>���?�,��^p,��9(�E[9�e N64W�-`b����j��]���ģ�����]���ٔ�_��@Ks&JT�Ȃ�D��n���C������=۲�s^y��V�W���� �b�^�l}J��o"�Нp���̰�XK\ǄcӀP<K������/(���i����P�������NF�y�b���U�!8�$*����f� ̵�g��ʋ�ʫy���y���{l6,K��R���u0�O=�&�k���+��Ț����h���ІFE���m���Yc��NQ���1��c�ē4�$M����Xz���b��W�*��P��S���-6r|2}�8�_O�SYh����] �^�g%GS�b͏I��,���e��D���m8�Wk���B׆(�BV�E�EU`�.ǌ��"�˦��__��o�Oq� "�Ҟ4���ݡ�띴X3�%ڎ�%o����	[\�2=��j#�,T�+���R*�h��
y��{L�� ո���4��)�e��n����B%���S�G,�[%c�4�p�3A:z����" '�j��WĽm{@_����w�7yIZ��7kz�4M��՗	�\�1"k�W�������^G_��@�2����G��0���-(+e�xl��c�l�^��S,�|�D�_K�Sw��T���]r���PW��D���V��,��<&��ߧ]��0�Ol1�bW@�uu�Q*��cyF�_ĕ>���_��>g�Vu2*��#��)[Mq�i�H0p�at��l�Y�,�s��˪t�,�������p�!	�z�=Cל�Ν��,<E.t���9\P�����!g藆��G�.5�ZϮ�ۻ�) d�E���]\Q�w�Jk�4;�D͍L��T*��-l���XY�g;%� �5<]�:����^£����gV�)n<S�xK��� �S��$Br�I�%Q���D$�Å��h,��:�Y����Ρ�r^F[0ŭ)��L�aӿuP/>[��28�r��o��8�K/�0%�U��8F(y�����qn���P�I׻�$0o�'c�Ò��O�+��ܣ�탷�1��c�C|6j��e����|^K�mKT
�����g����
m
����f���I؟pj�k(B Ƌ;ig�r��vgIeC~N��s�A�����������2�!SA3��jT�_Yƫ��-���ӗw�K˸�?�c��~~2��8���X�Ù'-L��̃��ouQH%&�C��-d촆V1Pẉ)c�´�kiE�pK`}�.��v?�r����y�/��,�5yd��	�6g���d�Z�;d�� �i���LN�S��+�b.t��p��d�'��aU��قV�K�mf �*�̝{�O��o��%ALZM/�ף�y���mC�㴍	2ā 7PWӆ�������*�|���=S��Xx�PMk�Ŵ@�d[%J���p�$tV4�3��~%�qƺoUgo��dXp��(�fʈ�H���ɤk@J�S|l��9F�����2p��]ǜ�,EB�=���P���R�<��������B�ot����u�aR&�:ո���y=&\����'{>!
DD� ';�W=�S�u�,��~�{w��Y-x���V�*���-�7GG��.&,ư�5���S
�zTp����?҈7��v|�T��G$�9T
�e�c�7���ڊ��;O�P۱�B{�ᖈ�PQܿ������)��y�q����=�r��idg%Gr��{'�sއ�^v���?�#`a$t6�t�M���5�eo�/�)�R���웱�L�-r�����[&ίMT.�D޽�Jӽ_l�/H/;����h�c1n�J�ټMQ c%(=g��E� �Pu.�eݺU<?3�x)!Zo��7��ym����3�C��1u�(�ǶPm���~wd\�!B�Ǻ6R��U���� �`�,2���o���t�c�Y�>��������{<<��=�S����5 �Z��&P��ɖË4%��X��ޟ7���;^�m-o��h�^8ܮ���4�,O��+YT't���0��k0����DK�U���a>��ux�����P�.V��pf�Y��C�ʵHĦ�MT0�	�ͬ��@����g2��e�+{y��wj�i��X1]�o���&�;��.%�2g��y�{��--j7bf��k�b��7kV՜m,����AP*?��v:�ā���4���{:o�E�����C���E!�b�4l0��(���D+fG%|rC+���&�$鯙淁ȯ H�y���%�m���?���y&9Lν}��)F̱�V��	A���u���t���-���������jٷ�
�����|��ׯzTIi�k��kQba�3D�r�f7�2U��=L�_�q����9 ��E�J2ǍQЍ� c��מ�:~%L1ؑ��Cς��4~�r��F��J����*l�ړ���YB1�$mHDQ��4���:����x���B<�����
R԰�B�@[?�jUTҍ��:�점��Ҫ�[u$�����׵Jx#��[ׯ�Y_��R�`��V�P"x�j�Z4ΐ��V�}E1�4����x���8X�� �l���Ƙ%�gǰ<�n9�\�_�4u��6����n�@Yd�Y�Z�*;$���f4͎�v`{�6�O���~"��t����s��6������0�T̒�G����{29l�L��
Խ]�����3o0�r{�]�~t���)�������(��L@^J�]�^��a|�D��b�B�������SK�
n�P��.'Z��Z>�IQ�z��%Ah�#�LQ�ꫛs��y�W@ԴE�=����'z�ʷ��E�|N��r&�����E�?-����6mk��P�e�j��Ƥ�{�L�V�C����!d������C�ś�,�q/�9]�9�<l�9p���/o�>�>���Sf�h�h7lvr������q��Od�p�5h�Ng��>�0��0z&�l|�`ś�� ��]~aX$f|��qsƏ� �!�\�t�{m�{o�4��)~���Ͱ[��B�@�qO�~�_�}|�A�Q�W����}�0{Q]�z�N$O�8�;��*9g4��T��bzF�i�W����sk�+��Z�13��&Z��|���Ϝq�[�H� O��<{�G9ۊ��Y�1ӻ�lླ��Ř�Gگ8!�X�#��`=]ͨR}���k.�T5�h�����*"��</�)���*�ȕ��:���ºp5K�wmW>�L$h,�4b�e~�@�_��*.�$*�R&U�����Nl�:��<j(�D��N�P�!Nu�v$!d�ҹق#{:��d����}#�[p�"m�~^|1A���k�}�.��q�/�A�I37
{*�?Y�����p�~����s�ħA��&U��T���Dܣ'h�j�;���'?Ȟ�K�wE*����������׸eic��hk��7�i	�><�?��cw��	a�49M-��|�iL
7$Vu���ң�ϙ��-F���-L�z� W���gx1�B).C����!��{�P��W�z��[P4ρ� �>=���&#�m6��J���[r�I<<卻4}h�c�N�)א�G"ӱ��P�q���.����?��f���P�m�d&��G���@��3���f��?�&���1���<ýcr�=*wR�᠁d_���0�I�%��|>xQ��#Ï�<�ti``5����կ?[�,��V����9�.�U���Dl�`�z��'23�B�HK��L�@V?�to�7�$K��*0e-�ÇhvdH�n�����h�=�]�%|�3D�L�4��n�����q�L��";��h�h�(h���)�I'�=�M{[w���������񋱧y�r��V�ӽ���qr���7jOgj��z��x�Wk(�[?8��:�+J���E�?���^�=��P�Ő}d�R��E���&P<���4Ν�I$]{��u�zۺ��k*5w�4~��������L��ū3N^����S�+<�I��Uw��6����%�����~�Ш�H��ۮb�l������ �J��!�PD/0��i��KX4�3M���{��,1���le�o^��i�	�[)�摒��'9�]	d/�c#��Q�+mjO��之f�n�->����#{Ϗ^�f�乛6��Y��!]�f	�K�-t�78��,y[�)2�(w�W�}$�`TVE��P1Ɯ�*��{���C�l}oT>J��Mo�sqO�0���?,ߖZL+0URh�mu�����u5AFS�Q*��zw ��`Ez�%&��h�(+���\O�S+w7��b�.T�ĉ���@�(ۺ7�jd^>���x�D}u)���)�2��d��nХgPi!�h��#.�̉2kY73��&|(�T�_��P��fC��Ӵ��FZ�')��+��)��F�\�F#��۵�f�;����=:�$�/9�I��p�*�6[�/<oX����f�7p'�xݚ�	(4<��D1�_�+ y��	���a��~�>��zz>yJ���2vq!6�ҡ�_P�T�����:]e��(ӈAX�5͡�%�ɤ�8�^^��ݳ	w�O�O,��M�ϺBdz\W0��&HB�Yʞm���@ ,�[J=��n�vq�����q��v�ˌ������ب����6���u��3���e�����3%��BbDƧ�Ap"������╇w�e�p��{���9�:� �����B��2Ըg[��ꔽ
C��m�l���Fގ>G�\|eg~�r��w�U@r~G�� �a�OРi-�Χ�m��n��Q�H�+�B�&Ҋ�лkZ��j/�6��g#�8T��>�<Zॽ��:h���Bw;kV/��uA�q��Ø� �4�D)����'���\ ��SW`��<Y)�f�8�����l�v�("ѧ8�ut��n�* ��jW���l�����w�F@��g"�a�=��sU(Ӷߓz�9_�O�'Ly��0<ړ�mh��<ۨ	��:��x���^g���Z���Il���-*%�p�j��h/�`7Pnn-����#b�F��ѡ���i�no���E�TˏP�]��b����鮬��a=Q|J3�u�_}���D�=� 
�|d��U$�����f�D=9��C�ȶyK\B�(�|�aב����#�N�|���3�^������,��@�''v�k���W����[�JU]�^����#ŵ���R���Сā�����>��Z�L�_�J[�}��I�~CՈ���Д��jvRs/ F�v̼�/�'�����Kj� f�6�Th_9�nE �r�j��C�%d��0���Y�d���]k/�9����-�g�Č]�R�RK4<�uлSu��Cr���5�ך߃�+4V�%��C�e�ϖޯ�_���ؤ�T�.�ڦ��@�)�@���9ȥ��'��\�
��ƹm��Vث퀄������}��\I�^�=sg�Nq,�řikp�\?͏��w֧H�) �ށC�}pk�p�LK��-��
�>'Y7���� ۈ�
��_��4�r��M��)w��SM�e������{��4�������x��]ig1�����X�ѩ-��;���P6�_rε�A�T����_*�SqLR���<���G�nL���u癩A�WZ�O�1U��-R ԭ���Z�n�'\;��%4<��.�Ǭ�@u�ȵ�eUH'DE�S���ߋ�ޒ�$2�DƝ���4l��y�w��w� >��XYwP��Q�'_�_\ ĕB����FKNk�j��3�ճxR�C'�LkG
3"��QC3¬��G'>�9�= 5�!�]9��mS��xD��`%�Q����M�5��U.+�:
{S�Q�m�C�{5��i��r��*�dv_���ް]k��}?)\����	m�V�ک�<R��t�/�D@z�� �p�$��!�`M���ے"��H�o��/�|�w^�@�ld�1Km���3a0J�E�m�Y�[�Y��We�� 1<\E6�[���Pm]>=����4�Xw =T�adi�ST<��1��l��K�H�@=s�q�.�r�s;�a�"�<im��k8������E^A�ZR���5��BN~�KS
��K�͞B�5��S�w�sU��kˁ���<4'�R<ʠZޮ�qO��@waA������
5��'
1P��V='������Z"�P��H3��=���6%iS�vJ���w���H{�)�~YP��e��!�p���kΆ,�5\0/����n��/�ԏ�^�!�7��=t]np��NH!D���6�.ޖ-������ct���5������ǔ�s�#K+H��c�0�X����5zv:1 V�>`E�=a.����������h�[7`���J()C��G�+ȵ�����&?��[.�u�h�eՖ��j��a��6E�@o*y�	г���1� _��ꔟ]e�"��A�������s�;f�#�(��X�z6�j1ΝM3�;5�\U�G28J���ی��.�)U|�(aI|B�{���8�>� =�K�E�_i�Y<�@[�&=]�+�����7Q�C��������V�MJ$��N ��@8����Ѫ;�a%Z3D�`�H6�u> �<{�T$�W��"Qm����׼QA��D���A6+[xt'�βQ ��ɬ����D��o�Ac�)�V"{c�:�0䳸И�j#��H�p�\�8��ǱAaʂ��FP��M�+
{��iU2��L{C�&�\$9�fR��c5&��L�%+��z8i���}�Л�׊T�{��r
En�Ye�x��X���c����$��SЪh��YrD����S����]�M9S�ը��b��(�ˢ�������_�
D����%D�o������cnnm������VM��,:�>�T0C�Z��|�G/S���,FQtw��w1����F/9��e�'E��o�%Q���ҭ�zMu1�M��`�SA��.i��r^��~5�Q\2�{��k�]�����כG�2��THi�؁���A�e�]z���Q�Kq]$�f0����	�_�*��"��C�x΋�ppr��ܽD��M#��Z����� ���x�"{�J*�wP��_�+�>�az4{���%��]>�B@����b�z�%в���]/<�9�0?Q����ߕ`1���W��&�ff���8U.��l_)sl�fʦ���<�@9WU�ң~G'h�k\���u�$�Eߋ�v����K@�A�+0��t�%��ƳNXAs�8RX5��}ZQ�yF�w����H�z�./@��f�*��3U�-��}�@�hm�r�f����Ca���mvw.����:�H�e��&߯-�t�ėk^5�Ѭ����X��[e���JC�r�!y��'�!��xC��7eB�J i���LI�O��9I0��i^!�r���dl]$��~¦δH�gqr\C���n�uZ�/>/���C>H�N���� �20��������j�Q�ܬ�$/�*��/�� ��BL��T�א�1{��@��#�1��Zy��,�"^��Z�(�<EL���B�f�>���h�������t���X�R]#S���<Y	�?�W�t��W0k��q\�>��d6�}�~���q� ������ߦ��B�H�_�Kr��ya!�L������A��y��$t�:�Tl�M�StsU�5�V[�P�7.��[�Z%�������f���8=�N�;ቍ#�S���!U�e�'�����9t4�C������yV{(�{����H�cPX{�%��V_q~J�G#v�J�t�Uʿ"�DJw|R8i5'�\���-��m'������=�dTO箋j��"�m	���������@�z����'5�V�8��Ӛ�dwDz�y}��x�O�z�=��f���x��
��G�5��*Y12�n�j�O���'e�n���.�(,��dm0�n �p���nBY{ɤ�1�q�C��v-�x��g���t>����_��X|��fc���	]�UF@y� ͆��ժ$?k��1�svo\˙0*"�>
)>�:��g�%^T��&��Cr�-TT��wF�v��Q[G��lx��rt�/��v���TGK������T�7rD9�G$��������<2M'�H��3;)����~(ʞ}��� '��5����	LX��$��s�!3TB�W�v��K��	<2+�r_T��x�Z��S���{�}˖J�������J���I!��Q+�K�u[�0
y]ƴ0�����^r��6�V���0I���o^!�ˏ�61S!�<py�J�誧���*#�"	�I�KI���µ�=3
f����(�y�T�M���Pp�dR�>��ne�`���'*Ϧ�1����"�Qkov{Xi�����K��::(er�!�%�8�K?�jO$����\�>�)�/��������-B��L�m�D}
�a�),FI=c�t�T�Yʑ����:۰6fU�l�=L�Сx����d���Bk�ݚ����TuxT��prh�7�v��޴]�Zy��ŋ�ݔ"4�W��9�5H�7��o�#�T����o���Sc'��o����4���tS[.r�)���ٙ��-Y��W��/�Ӛ��)����LtW{�x�Ѯ:籨�8����]��"y3�����y����m��I6�&���92����b���������o;���e��s�H֖r!�r æ�<�
=�zf����p��$�ܰ"I:����Ɛ��H����!W��;� _~:Q�|��{�-����2ʻ�,�>�H@9�OV�!&<��!Q�ן�2ƇbYKK�8vl���,�0 �0nWf���B߄�Z�;�h���Oy�2=)n`(>%0��A��&�9&����3�ߋ��J$t肶���Z����?�|l��^� N؞�2���g���׉����Y>0-��qu�VP�i���v
��D9��w�U\gƏ�a�;;_H&�-���#������T�%IH�����TB`4<�v��$�� J5�����^�N�*r�"�NN��+���0�Z�#�k����/��O��5Rʶ�y+��=]G��?�sJ���.po�F�����fv2�J���h0��m3��c}sQI�=��4�|i|d������!S��Ȼ~jP��C���d����c�lE�[�vť����3�x�(�K!�O����.�Q��<�/ݦ�C���faOV`��?R9������z�-P��1m�^gA^�2��m�a&��Qp	7���1x-t�>>��&�����b�����W�J���	�VX�y3�«���_��Ezߖ�#�sX�yA���oA�F��!!�m^�:���F�O<@k�^�����(9����N��� �z���%��T�AƎ�'��P��涪���	pz��ֽD�rԆQ����U�7_%eɴ��V��lL�,�멹����ZQ J�R�3�!T}�����o������(7<��ҍ�9�&дrD�R���]'�@�:z5D����*tr�,�X���iU~�u�N��bל��f��|��Ei���+��5�_Z�Bm�+�Y7���6(]�qXk7�-&�1ذ�wH-%���Hp�*W:���~a��BU.�rC�h�c$nL �F�/)��5n6����E�ߦ�ĉ���x�2*���d�����,����|g���tک#}�������O�"���f�
n�k	�����`|���.�����7O���(՗ �=�9��z��[��~�I?k����tZ�FZּ+��x��ø�x���o��^�8�m�NR��c>YI2~<�O���'�BR��_6���z��C"@�+�*�9fT��`
}�u��@����V����v��{��9��n[1P��[ї2a \UX�B]'yCʒ�73S���M�ߖ	���<~NSqx~4{�m\`O�<L�p��М̮�smb�
n��W�C��XTl�I��EN����5g���l&��N��(���HD�c"��f�ѡ�"���/"|���mK@hqq��wg� l��C�-���atF+E�n#1�T
D�Uy�����-(5=��;��2CBUe��T�t��Ǣ�_-��Q{l���B��<��cϱ�e���MK�qC�,�Vj߄։���L��qbk����ǿ�W�v�i7-ɱ��J�Z�!��͙��W�%4 ?�0�|H�\z�H����I�'��2JE䱿�Y�LH���u�2��������f���/`�F|cfS��"��۬����$�<��C$ī>��:�BUJMW-v����l�c?��H�����ħklfZ �J���hA�rt!cV�(.P�E*����+��Z�M�Ԡ�^c���T�s:��1yl6I����Y@�Q�g���57OC~�lV�KTS�_��l�l;�u{���Fs��u�ގ�re̡�sw�C!+��I�bP�w�C����|�Â離��0X>��?s����э��1���y�5��(�B�ы*�@�v�rt�9����^�<=�a����ؿ��S���H���% mB�i�� >���)q�Ab�T	2l�����Y:9ng�=�8DrOC�c>�MPD�9ۖtnv (�B��`����d��ۉrFp�4�gk�����E���k�R� �fP~�ZEk'���t\3��i/������"_nk?� �<C�	��YE�j�wzWq���sh�$�t�"�β&(C��F`����|�q
w�iA�hۀ�`�	O�]�u#ׁ��o>���P�l�����R��Է�|�hO"^aws�Y��>]!�������j��
M@�����q:��K��2Ɩ�+�K�Q�b������X �:���W���`0,���K�����TO����ȍK��*��/	���蠝 �I�<��_W!x�s�>�s�Tٞ��|h&3vȫ`��^q9'��vb0����G�2iO���2ٌג�1����*~�#R�@`/�`�*ɗ���*55i@�aUy~��S�"�m��	��<Q�L8%�1�(^�.w��_��/�0ţ ��JD�otB�A�+�.^��g��֘�tU9h۽X+*f|*T�&�mz��U���!�/N7?�q#B��Ү��T`�x��U�T���\m�B#�~�Ɇ���[�����h�J�+�8~� q����׿S_���Hv"'���A+�?�p�l�U�|��Q'k���Xu�b�H���}��6,�_ U��A8ŵ�[�+Ux��H���'%�_;I�,�D9=��6 �]����ƲU��Sx��Y��_;���*����$�(��lJ��%�v^���%�iQ��Dc��!Km���ݬ))�k�r�z:uc0���+.	���,�Ԩ#*��V[����T�l�����%��;�&�c�G|.A�&�����{8>���8�6�$���Дe�9�{�>�]���窊��	��;��?7�:��R�J�=T����1�1�ۥ��j��S?j�`��W)-c��ug���O����`I�(	��� ������_��1SO��3�ux<��5�f)�0�KY~�P��d*�B+�c�c/'��/nF9��Q��2���0Z'����$Ѷܹ���zM�-�Z��q���D�������i��˳-%Q�-�;�+��ù-�8�O�J\���[��c��}
�ͣ�X��;�)R����"^!�^�e�JF�t;��ҠC|��e���a�$���-2��)�4�i�z�Bڇ$md�uE�,̚ȸ.�ʊf���lA�^�2(�N��!?I��1e�/<邓���{�$���!|y&���{�� {��Pz��WUu�Y��'��Nr7��W:�}<F�Q�K3����Jp���������j��q��ul���oM�<��0lNiS�����J)xr�w�|��Y̖����� پ���25�s�G�ew/]끪�X�<4HQ'�z<Y�<��!՚^��v�c��V�����o"�wL����wCc�KWc8EL9}6G޳z�xh*
�?n��$�@�����{�L�RГ�0;j���k�)R�������mQ�����I�n6��.^'��$cb4��>6b�᫾�������Ѯ/>�\���O$��.�+��o�)���E_�I�2��˹�i�vvlm��r�g��P�I��\��� ݓmS����R�)�N78=z�߯�� PN�B����~ ���En��In�C�(��ϗU���2(}}��lZ��B4����@Z%�2���W���4����Cu4x�(oD�l��2r��&y�3����3B���_���zFiAΏ6��o���I	ˡ���=�L�1m��m���@,^PO�{���rgK�N:HT�bx�k�L�Rdq�]sd֒�.Z���]����c�n�E��#�8�%ܾ��@9Cfշ�Dxߘ�O�{�R�پg�{ޅׇ�����a�=�BR����}�Gs't f�O+[�9�����~W!�e��ϬT��bv9ݵ5QXLVҥ�К�v[_�~����hb�V��V �ǍMh�n��ΥN�#�~�>����������cY8��}�@�V>�ܕ�&;�?a��P�-�w]�_�N��������#?�]�zۤ7=$����1֕�H��e���I3�"{Ϫ����c!߾?����Tw���R]J+(�qi�مmQt�v���Q�Ǥ��F�`l퍻̺�136�VU�Qs��[â����7l*�G��kU[-��.Ӣ+��
�y��-���Ů��vK��c �����߆;�# �R�5iA�*���)qŹL���d>��m]��*s�+l2~��K��-��9x�A��V�����gF{Waخb�'|�.u#B�݃Z�%���Y�i!]V���o��t��a��vo@�`O�#����I���� ��L_^7���mm��3��M?-�Sm�`f��(b��Q#{� ��#�����a��"�ꨜ�J���H`�!�g	f�s�=2� �3>qH���rc�p��S<��(N-��?��&.c�P�H���q$h?ѝ}	��D�*�?����U�sP��"�� m?�_������4C;/z,�/g(W�Ni��o#,<q��҅�X�r�Β5	j�Qx�%_�R^���Q-t��{�����X���cU�:g�	����Y�����Z�T��U�c������#Z���ú4�y���ܲ�̓l"�O"���8�9�2��X���F�&��x6�m
2�%�1uIg�� p�N���}�dxr��o������Pa��'-o~�
���\Й����j�o%'�Z�n�UOZh�9���q�t�['iа����$oބz>X���T�R���C�c�2%����PA�M��gB%��-�k
�`�{�8f�b�Z3���(�X��z�G�\��X"!�f��V�T$<��$\?M}� ��%�
��"�țU5�tXų�����s �f=�Q�A>��U���g��g����#�;�|��^4�w�ܷ���CȔ��hM�r�W��qa_D�~THA�
��{�K��Ϟ���p'&̓���e�GѤ.�)��m��,U�E���n>K��j�c��[Ǭ�s�/��t7��O��^�jYהd��k��F��uǩ�u�3��dG`7�U_4��3I�h���D�O�S�1��	���RZ�P��m�R�@؇�����l�3-岆�N�����[�flZ���W��<��W�e�
�Y�z�=��f�~�^�b=䑼���PC�9��ޯ��q��;��wE��]�#K	Hq���YA��i��n$����4jQ2oc���K8N��i�a�c�Xu9�]J S.�g���Ì?"����>��g�'&|p��J~W[�F� �2�B���J�T]Ivp������؟�?3zZWn{�&�3��S���|�஝ޙ�9pح����wD4�>�c�Y�N��F�E8qX�x�	�"��4h\���rX)�[�]��� �5�_v�ܶ�i;l*���.�؜,���nGe�Z�=Bn�VGK'Y�5���g
|�ۄuv+2;G$ϡ���e���W��.��T�U�<0��{��|�,�&���ٺg�9@s��F��}:0�V%��8��}Az��W�	nXa��ږ1�|��a��u6Ƨ@��d���b�*�p[e�VAV�dB�}D2=��р�]Y������O������n��/�H��Ta��Y�X�����s���Y�K��c����Iv
�� �p�q:|gwŘճ�p�S�����~w�r���B.��TS�[q�#�_�P���/r�`ev�1���B<�ý���y��� }w˫7�_oqf�D����F�L^0�����?]=��ꆢf?*���W�A/���	�m�n'�a�Ȑ��=�U(������Í���~�]{�j����nyc���+b,6=&Xͽ#SXC�נ�A���L��Hנ��0gnglW�����@�
Z]<k�S�$=�P���>�2 �_t"X�$��Aָzs0gAUz>g�O�	��Ҷ�1-r�x�PHf!���.��3Ԋ�nJw�)^g�N;*�t@p(6~{TӇ�=��$`kɬ�����p�c�o��CO )���-J2��t��k��݉/���I��r�?�h� ��~Ҭ�6%�E?3~���=�7�-���ښ�v����4��p�6(�AJK �7�sx�OTBy����{��EA?�c�\��فD3pn�y��6���p�{��^x��j�Ԫ�hl�)5�-N���I�q�Hx�`���Q׆�!����ݲu#7 ��<ە�|D'�����Hix6\�}m\��G�66��׹�o��u�3V��'%?�V����s.ޜ�#�_qfM�FJhS/rp���t�t�㻼e�����US��}yF�,,a��c��(<��xe�`I�[��:���Vg_�.��廆��2�ʼ�\Ly� ~!�y�8�y=0��!c�ՈRmi��ռU��-Ϭ��=����l�y�c6��6��i��\�Ls]�u�����(֝��ؤ�G�qb٫'��Xn�|�d6��������~��Fкh�;���{�N9y��	!�C�oo/ƨ����`/�kEi�����pK���X�]kLD�&��	D5*��Tog�l��O����
�lЍd3@|�q0�7��R3���_LWL�[F�Q��T��ѱn���q?�V���:���pU���'t�U},�G8�N^ fEE�ݎ�6glˁ� _�If�34��wx���m>�l>�F-�K0'C�{��Z7��@��B���˚T��h㻑�*�g8�1[��fHltl��W��-P��D���"* s>�/5�v��� d�R��m�����gF�i�ZbU,�����[�v�A���Hg ��;,�_�2jW��|,�0_��]�p�YR��,��;Т�_qpJȤ�:���AF�U&�R���Y�#�q�gT�O�w��$`�7em�`! ��)6 E��3\݃�#���:���JW�Hc�P�@��|�H_A{�a�Ӓ�^�׿��@�S������R��^�_�cJ׳�!oB�6n��`]������r�>A</��T�-ۯ͙�G'`JD�%�=6C.A���� m�*�u��)+a�{*{�ڀt�EB�q�&�V��#�(ȓ2,J�d?V��R�(�h��lߎ5.�?
�����
_��	³w`��'elg�#W�VTn� �V�P�y4��^�����Oc��M^�(s�S��44eo�"�o��QN\��x�MBU=QX�M���p���$���ڀ����٢��H���jw'�i��l<��B#��ս{,�����Ӻd������u��y��S�|zw���|�q��g oM�J(JegїI��gᰑ�농�1WB���l<����Q����O�6O�^��/�^Ll�H;Mbhul�7���io���~��8J�F���!���4��Ļ!u���C/�(z�_4^�sE;�ġ7D�<%�}i*����#�g�7ep�Ƈ����}$����J�߳�Z���,r���f �_?\��K�Z2�d����� ~w��4����S<
�qz�	F������� �w\�
�c�bi��&�M3<S~LM~X^^��v��w�p?r�V��uV>������2�rb�7�VE>[å,����nv�7���-��բ��Eȡ��MSB�1) 3�Xcfu*O�_��������-�a�r���>e0>�>Şgw������h�<Oݒ
bmpZ�i�:����v��X�0d���.ۏ��,�A��)��CK�4�3;�}uV.����@�:/rC?g����V��VRo�`Ɔx��T��-�qB�$9	�)?�����,n�U$DWR���=����L���E��t���Q�i����_^�<���L�`�] �U��o��Bu���
�Z���� �ӳ����z8#�ߖ��|�@I���wGr�� /������h~Ev��R}Q��h���.JzGM�(VQP�j��ո�s"�c��w7#�I��7۳me�S��`��|(��툐��e1�#��7b%���]|����u/�.e��\G���%-2�@�M���������+<<���\�Z�O�������拶��.�9<H�4.�0B?��F��b��C�v��?�� ����H+~����(v0���^䂋<g��~���+3�J�B��|���U��\��L}�Cx@GG�v=��]0�N:�f�f�fҊ@��>�*����-�A��i�Z��.x&A��~1�9�8��w��[� k-FI�t�x@PU����wZ�o�R£��P#f8��īéen��Q_t��s�c�L�R� NM�[Sj�&�}���Uk����n���}��m���ɡ��?Bp'?QR9U�w�7�(�K���Iǌ�"�Ju�$�����6���[��<��Y�~PR2�-��nȩk��M>�ַ®�`�p,��l��Ϧ���o[l�tVy&��k�2��3���;U2\����g�9]��l�����ثZm��BL E���?��A�ki��؂`���u���[��Մ@#���O����!���xܴd�	5���ju6(�N1�\��k�&`���%��?�,~,5)���L��Z�~�r$k?ڻ���w�|�jÞ��%[���Xf���.$�Kޱ*Rz�ԇ,��Mu��965"���%TJ��ۈ��jl�35�g�u_���i%	c��Ŝc�:ѿo#��Ӊ��d,�U�~3���ш�E��?���W�����4$���Y�z�?��
�CjҨ�S5�01��&w}�!�! �(�{�.�7ڶ`��7��D��^T��e9^�l/8�9����� ��R���a��N&K��^(k��d}q�ɸU�6Z�n��s��`�{�hsKOD$�;Hz�#��rd�Un	���{�;z?Ft�CU�m?KoD&��#)���|�sk��B���
C��P!��Y�s����y�\�1K��К]�1��9�u)b�1�X�;�tx�ܥ/	R����l&�&T<�L?�Sh���/h`pQ����L4���?Ȉ����zR-�!��?�8��bd]���/�2���~7�nF�3G��T!q~���U�Y�]eN��u2�'k�g�`=$A�&�RO��ĮaQzIN�BU�h�yz���V��ڐgn��V ���M�� f����ٸA��X@ ����ڮ�4'[����Ǜ���ъ�c����Kt��;�����p"?o�^/�� �Y�&�,Ri?y�SQFk�F��/��Y�"|�(�"�.���-���sө�}��Q��6� 8L�e�'~�(��7���/D�L㗝�b3
i��o_l�=&�,L#4y(�psAM���w��t9vKՏ��G�C�a�O@O_?'f�5画����R��U�{s��w��"��pM�X�xk�$W9�uzh�2~�.�rZ���L�~FE+8�k�{�E��ǡv�9p��wW��m��Y�w�� 5"�M|N5�!<MÓ@�߬i�����BpBEo8O�#�$~����4�F�a8p������'_�M���K��>��*M���0�nR�I�Q�.(9�4o�}���I
r5�tu���~GOy�i�m���'�����)t���tC�,�7xE�8��-Ё����2�%8��D{��i��G���$���`\����<������b�v:"�w��+!8�ΉAX�j�+ 6�!:2�MG%������5����+�>�'$�<;
�����H��N|������f�"�~�	+��5m©��8���H.����>��K���D����q,��/��F��`�ʜL.-�	*�f��d�(��5�;)�ܷ�;1p���B6�G��w�Γ�����F}�C�c#��F�#4e��A3֥ޣ*��)���������W����Q�e�9�����u/�%��:N�ä������Wxi�����	��_C��C�a���3l��իT�Cuf��##Cm��J�!��%������Γ���-��a�=��n{�˂RYL�(:Z����(�'�8uu(xQʩ�),o��͛��8�2�'쒭'VxS�������"m@ȸ��hR����e�@��8D�x"|�= �OsjX�֮���]	��E7:�h����,�I�X�W&|&�*G�5ɵO�����J��>�do���)0s�h/Nf�ҿ�-�$��Q�@�c���/���0�Q�"MC�e0T$���b�M"���@^��{F�G���>8��m��BG��YQ�]'r�{F��6�bk�������K_�����������=�g��W�V�*�7�"z4���&��_�����,R8��V����E&���xQ	C2��X�2M�:�a��X���avD����أ�f�T�a,��s��\���xF~?&M�N���?���)�M������t��Pa��Oq��o U��W����@b_��2D�Qz�:�Y���Ɏ��
`�,z��*�+O��C�xJ��w�S��'#.�(L����H��rf^2��cڟ��Q�}����ZDyE��& t���lT?�e���*�2Yd������-+:�&�z�z�5i1�����yp�#ֈx)ȘX!��b�v]8ptm��
�a�~d����̲��~�Q`� ,K�`�Y	�%��'��\��k�����B��y�	�aR�W$,A,S��K�	�&�!�i�6��z9ў�$�$��t:��v!l�xk3�+�J���%�H�n
�Cr�?<�l��6�����<�q�1��<��	�>ճ��4��Ĺpώ3%�{(������7f`V�K�=Y�uo�˰�u���6F��b#�XAOb�m��j����<y�g�m�f�T��o�*{Ӵ�VC?��f?ʕ����G��z(E����q�!�'��8�@UA�ڦ]/?�̆��"ES�exi�V�WtbPz
*���C�K�������42��/Ы�[�R�0i9D�T�
h�}G��HJ�� J���w�	F��r��#9 �w95�Yy�H,� ͤ���#l5��Z���X�Ȥ^�5��S�zpix��1�Rsa���[ `N�Ii�I�&Y;*��bb����%�3r���I����A��S��<-�Q��YZ���a$��&,�����}X�Ņ�˭�G�H$F�^p`�O��!B�5]�}eK�>�Q}^�3Q?U�K�&��R����׶�C�˧��9���Y�}���|H:u�ſ�|�F�J�
�U�&+n�/���s�/̏B:��\)�A)�T8��P�.a^����>��*>�W����'�s�YeZ��P^�xcp�%�,�!v ���LL�cq\��}
�҄�:)��R����ǰە���kB�/�+!7ـ4����A�������c����?ZHϥ_X��sI��PD��1�G�.-s��0�[��L�Ϛ���M�V� CRo�wUM&4 V�ֵ2+�=� ������� �3�	,'���������O�S����E�K'���߼;�XM~�	��!=&߀!4�F��{!�z7��Y��|��`6^+ލ��M�K;i�-$G�F��(�Z0�ShÙ�0B��ǽቂ��"���5�$5�i
kr�q�x�$��4eめ,�a,����$H��"P)���+]@�LF���\9h�Vn��B��+(����Ի�|��\�zģ��π�D��# ��;�5}v�5F%O������Fm��p�,�����y�G�O�i�8�k��}��SW�H�SS�K�(4�A"۴��(��8;YC���܁n��ȡ�]c���� ���E_V�/�=��f	Ϛe�)�W�׮ŪJcFP�)!�z\OaA�T%<	�}�qwL�0O(�6�+�}y�+�ʆ�"D��a�5d�aWPV���MPgQ�b �aK�̂��p��\('�9><5X~�Lz���i,2�K�b�S����`�m0���4�"<�_Z���%Ө�+(a��}�O=��7\Y�G�s�T�\a�BB8�~��k�m��_���9)IM�R'�T��^O���g	�2*�=��Ca3;>�U�Eg奅Vئ\! �$��[�<�tb����p�/�1L�2��f��~O�ۀ���q�zE�Cw�-h4�J�Z��C�w����h�-�t7�0����1�тò;���S���5�����E3/uO-�zl������]��q�n$��M/EGm��є3����]�kv��(�#)m� ��:+�����!��[�D�z	p��@"��on�G;�a�Œ@_�
}ʸ�L\�4<i�s�'�^-�H-�k�7 �؃&B�Ӫ.�ffa�<6cy�$,%O1v}�\N~��;�}�Q���S_E�LN��B�HI��"t\�mũ|���:���?��t,eǗ�� ���@�᪙��,���6�]ai������dp��/�xc�O%wܬ� H�]������kG%9��&|,E�ˊ�� Q�]�\�t�E۩R��ȵ��\-x:5:�S���u(X�����jd�ϯ�A�� w��x����r�B,/�a����u�m��!��gƺ��-��\D��B޺�\�,��:�?�p�Œ�ߏ�ug���,;a2�8�9&4w@� �غ&tx����ط�G����+D"�0��u[���Y~j�A�Ɵt^�\,Cy�ɇ�h�w=矍���x����2��f�U��9F����>��~��CґA�|�����uY.<��V�2�o����w���1�P\��W�fV���4�]��q�����:aJ��Bґk�N�r�����,:?m�3�o����{�8�/Y���]�&��"�
]��ۭ�X7�-qE�RQ��(n���; �ϡ5�ޝW���x�z2�ЪP44�&3-L�[������٘�m��;��Ԩ��~G�0���4#�`ִ9�}ѝ)�=H4wOWU^�{P�mk��P�b�����&�(�=L�;����B����s�=Y�v�R����Z����ҹ�wH���vwW������@H�^���1�&�����\�1�Lz����Ϗ�ip9j�֜~�D�Q/�<��$���%�=RS�u��� �AFh��MHRk��wr���kH/�[�Kj�Kpօ��	9�h�r��Q0�ف��ޜ)67�c+����K�tE��nŹM1K�\?o@8��.ꗉ�]���h��}�d�ع���,����^��[{�{$�`{�a��;�y4�<2HH�Cm5��%��q��.��oִg�^m��l?u85��hUo3�
/ឧ�<W�S,��$7.�d���F����]eǷ�?��Ƥ0��7�V�e
�`m���f�[e��˘�e'��+dcP�&���69��a�c���y8���2�0H�j��	e��_J��%(��._���>����鐞8�O�����sқw7$�JBu'!�i�G5�u�{2��9X�H��9�m���Nr�x���s�q�m��;�Cq�e�RTAj�Ψ�?�I��`����R�SUH'is��SB�e"ԧ9�_ ��^�O��^��?��*��( ��*��M�r�}Dxֶg��}��14����m9OH��F�Tu ݑ9���|4�� ���Q�+�&L����%k��N����>�7R^�v�*c^��t��'%BL��]e��Or���Zf���^ `v@M%�	~O�%.5��Y*�?g�se�,��r��{�kO��?	�����[�N�|��4��R��Ŭ��q��ь��Sa�b4�E!F�2c���y�z����3YX�������3*]��k?S����ں_a��4.e/���ÜŻ+�h�D��_����$�q�U�~w>>ֆ��ZT9Ľ>�W\x�C�=WD/0�b�8C,o��U�+�$;,󀡰*T����I���}��xb;�!i�n��4=����*߿F��7���JX!�J�<����C���vV�&�V�s_-��t�8� ���5�\t��9΃+h���A6��N���`�e�:{��:4��u1�+�f��YX��a�q��Pz��`�;�Y�8����d��%�y9�D	��5̧���ek��o����<_��l�Ҁ
��d��+�л�����'���d*��Y�jT0wik�jz|�KjL�֫.P#���Yj�:(��mҾn�|����Y��L�V^\ eͰH��Q1�pH�V�J��WN�Ej �G�9��k�2杵�rب�f�S��"i�]TF�Z�4$R��`�[��Ͻ��T	��e�]��W�1���.�ǋ���?�L,@ЄA"�c�9��>Q4H��3�*=5IHm!�)�~u�aȅN��T!=����~���i����lR������	���8���K��_�mp�i���k�8�S̏����,C�/#Z���2�!K'�kБ���,�&"	���Vߝ�eo�����Ԍ%����ƨv�C*�X0 ~n�=h��21t�����͞��Ũu�Vs���L��vŨՆR)�!�Y�ܗ���������m��9^F����k��c��o )23��Q�[E�xruj���7h�8(�Py�9� ����ͷL�`	DQѻX�ETF�B䕿����d�D�ђ��t)^i)�,��-ȠgB)ʟ���¸� d-�Y\;7R��{o��L ~z1�I
61��1;TO��*��X��n���I���	P�dE�{:���F�8f��[�'�Q��F=s��[1�n�v@�ɂ��2���aTĘ�
���
(pK�1,�<�P$qj��\�/�W�EM��nr��L:편�*h߁�Φ�@ �W�^���A���^]����	��'���5�X�踀�:�N:��Ě�B�a92h���Dt���=����T5�f��}ͧ�&�9z��	
�%Vx�Rj+L�%�����a(ED�a�G�\��䘌���QWC��xq'ӭ��z�4>�*����V*,1��;�`B�O�6a��͉pcU.�w�we�����S{��`Ї9Aʹ�E��H?n�@��U.��/��*�w����[�n$����c��6��%���U�@��&�y��"D�&BĹ���t&�+p��J`ҵH��.��������W�-aH�|�Ux-n�<��&e`�����fU��N�qqQ�_�˪ �YBq���)xyL�x���+�b<i}W﷤�Y�8ublNẀ�������-�ik�Ż�:�+���;����=��+,�?���<�3��X�� Idf�]��0J�#���:Ï�h�X=�7nk���yM���G\�i�N�2�Ɣ'��{Fe��Dc͘����t��z��9�r�X�|�*�	R��Qo�OB��-Cγ�����M����$�GM�q�� &���5���^]��EV;%$)Āׇ�7���2	�\$��������z�af�Y�i�h��?��z�u�f7��@_�K���B�ӗ�%@%��&qx�j���߿S�Fe�+��pZ�=�=b�����0��1H&ٿENn�Di|B�l��	�L^�L�v���M�)���f+�(����ߴ�)hK�Hof�����4y:�E$_�"��Qi��|BV�n_o`\�%�\���S�Jj�0d�_���a�ȚPl���*]bΜ 7�{�}�k鋓�C�ʓ��U�"��N�ǖ(�W]��tN9Eb4-ܓ���H�#dS.M��4<v!���ۯ#���	��޻fa1?P�3H�o*_�����H}�Sr3B_�qFN �r���-x㭏�v�UKg`J֓�s�Ҡ�a��@
��������v���œ�����sh�� <I���:}�f�2�[p�6rwtm_H�1jR$JQ���l?����������_�v�^`�a��u�S��P3*�g�߇ �$9�]�^U@��PcۖA����n_�����I%8g;�`��)L��ѧ&x!<��B2��g�BDt6��$�זK�ڕ��8WI����Թ�c�S�S��C9s�]��PF^d��o ��PT�D��}7�p\z
��_��E�S�
Q�0���CA�O�jpF��Q~�d���,[��yYh��`��cqO������C���#�N�F���%��QéuQ�7� ��U��0��6�2�K%�\y@%�5�>p"Iu6�[�1vn���/���َ2v��9��<�>�8��s����j?�<2jaӹ�Θ���	T~�L*�s��Y�
�o:Г>$ [�V�2�w��,_�	pR����L��2q��ɉ�|0����|Y\��C������m|9&!ԧ�a7��Z�9��Җc��q���̚�+>��7
���1�{V��&M��}�rJ����#�D�C
�Pw9���R�KAcֆ��?!��0�b��#I��E&��*m���-f~�i����T�VP
{��g�
IA�!8�,z��X/�$���1��3�k�Q!�%��j�P�e��#������!�s�EU�LHq�BV>��]	�?4��aU�*' �I�z�~|X��9��'N)42���_ ���.e����&� 8T"�ܾ>�_�ѕ�!�г��A����K����|p�(�H%��Ɛ�jt�|��Q�ip��Q�l܍����B�Dv���g����{�@E@�k�J>dYX ���~�M�
�ԘX��V��y;L�k��
�ط^$��9O-�e������ �����h��Zm�����~���(&���i�G�gM1�;�"�|P�j�l�s-��5n3b�h$��Z������'�XrsP�^盳�'��eP��`�4��M����g��өn�B{9ݠ`~�\���Y�ZAc5�&��,��d�>o֕3��I��;�W K��]�Fj�$lj.�4���j��cPU5�F?�m"����H���6���K�j�_�|X�J��Bާ��\ִfp�ݿ�މ�_:���� �"y�S!6�����^���4�wݏ���q����c+RT�>g��"?�s�C�r� $5<:X:��T"�5x"��R�o��O�}�vƴR����B)�O�'�[2T:��,��^�s��90�����-s�U�;���nd����L���+�'�oz)�ݏ�5�D��ڳ3o���e�K�E��j7��՞�����w*�&+�l��Ǝ��� �N�֕��K�#=1�qR�`����3,��QC%�(4ZM>X��)���
�C�!\�́�m=Z?�d���u��͒��W�'���k�})�^5 �V�kyX./N��gp�N�Or��V�"�C��wV��#��?Z0���F��I#��b&\A�ý�o�ߵ��!�م�*׍V�$��?�Kx[�m�1O��P)<dE ӊ��k�k�ˑ�hu�{�G@O48X䨮j�>����j�|���b��uS�c1ef>�x�?��ˁ̤�w�H�$�WJ�΋��Ҡ�@n�����g$��h��h;D�I���@����&��JЬ ��B4q���X�\��s�k��V�)�*�b�>=������/, ^���Ӵ���MZ�?�?2�e��`�X��n��&U�w�Q�^Ӊ|��y�v/_w���v�W;�@�?E? o�������iTA\�4�5�M�1<�8ňWq�� ���PA���;TT�D)�6ۦ��Ĩ��2�g0�M�'�!�a�LxkY|_�}�����s�@�q�.'j9�� q6%#�/.Ⱦ+)�,��%�P�Z�jj7H1�B��6�c�AL^�բpk�9ҫ�I2K�[���l�	�AgJ��r�$�n4�^�`�H��'i���x�r��"�}���Ⱦh����n�����gSu���^᳅���nf�h��5q.��H�Y�PW��%H;e_	]!Iل*�H_�����u[9�o��恂�q/��(����uS���	7ڬjZ=##�;3�f��xz_��+�^A���	z`N�
]JP�8r9��}�G.�V�H-s��m�^��yX��RJ����iA��/4+MCMK�Dv~�eqb��ado.�R�G<��D���2��i��k�ʟ���� 3�cG|)Q�v���<К6)�䅟¿����S9іLO��1�~j)-��a:r����$gs�FGe��kCT�d�T��?"�m�'�G�=�)�;G���%e�h��8�5Gõ4��R��kI�"'8�҇k�{�	����K�ܑJO|`!���Wm�/)Ep�fD��l.8_s!qeT���6���Wx8?����bմ/}��n�������I*����G�F���{�X� �>~����ð�,�0H� ��
����DC*?`ZHDr^LϦ�v��~]�������k*ȃ���@ �X�.����H+��l7�=!�;�aef��Ѥ����m�fl�#=��6�M���TʸZ�m��P��:�~�cd��֝6��G4AK3��x�C�(��Tw]q�����I�J����=���4��2�#�2\�ֈ�8^�]�l���!���~�Cx��t�<�"�j Ȏ���/&�N��0�,ܥ��X�+,`ZH9�r��S���1�ýn��u��3��#��8��a���і/�7��I!�qKG�7'n�b�Y&���J���}Ѹ��&��/��;�tR��N�~��ϔ����hHmdy[�I��6x�A}.g�Ƒ���'o	������D�r>5ZH�z���1]HB��v�#�6~������jS�#����w��'���|X�ս�) �c4��Α4��a.����V����V�$7�eƉ.�r�p�DB,����]y�t�e��$S�[70���Tg)]���Q^)��!3��A/n|x������b(Σt�,َ�ܧ2��K������fʧ��ك����wK?���mt��#c%��#���K�Z9+!�m"�~�?�����ǆE�H�Ji n]�WU�2��+5h�zc�e�5�1"�~��TU���p&3E��Z�r(�(��R%��" Jt�Mh�_PHJ<�6��y�?��x�Ui0O��0�-�Չ��w-���pܢuq�nv��1׋O�^���{{���\��#��h]u쎹��f���fO��d�&~깉�a�|���o�_!�
CO���=�Q��R�=�.`�1C�1�f�$F|�ج�a,�LĈ�"r߰v�������sw;b��l���[���ͮ���Z &	���O�yR���D��%1r�}�N����+����e�]<��3%�mF,<&nU���T���G�Ζ���g�{�8�Gt"wm��-3��І'�-��ݩc���7��\	������Q"�v���v���i��(Q/�5g��^}��`?i��^!g�y}� \�q ��υ�?��|rŖ!���j*-~���-��."60�ȴ���Z&����GԿH=��I��8�Mqz#:o��n�	HMrc5c~�-�m��{>y����?R�쵄 ǿ�9�D&�OV�]�24*��5���tDE�z��`�D!9=�6�9��\� :M�O�>�q��FB�j���ZJ���x�L;���Fo3��C�aYR���ݨ�j��N=Å�`e��|I���
}Y�/��L�X8ȯ�"�����Fo��`C�0%e�0��d�r��-p��pԷ�1�2�c���Db��.9���l-��DS��8�kt�S3T*/��s&$Q(��s�i����<\�pM:��mG��x���/w�S'))Z��gKCh:[ӚF���\���)e� �7���a�Z�Yxݜ��@Q_�s�os2�'�n���*�Ihh��p~@f��@OK`��sW+�C�L� ������r;k����y�S�U��P�ktU!c5����bz#�`,u�m�| w�q���E��Tʆ�
���l��x���5��&�׻�p�Ȉ�ZY_6/VA�8�:�B_��M�hA��ڇaJ@�<rHN04�x�����*����g����r]S�V�����������P����"��MY6O������ü��'v� y�,��nC��z�p7�ڀ���ۊg�Ljr�#Y��v���jFFwF,�̌�@>w�aFB����C{7j�O(l����Tz�`�3#�ƻ�_��==s���Țr����;RڽM�<M�Ji�'J�G,t�Bx����_�_d�:q}�*����f��3*�m����KQ��b�^M6>�.<j�gQ��g}��25.�H��>Y��D����&�dG��2o���!	����R�*F0��KzP���=�*s�|J���ͺ�<:����7�*Kۼ$�-gݬ$��&V�]��uyg��կ5�L^�g>$�;�,��q�3�	㒲�3*�X���ï�i:�ټ���v�m�mԇ/�u����i&���AD��.$�s�#͸�(Ӓ
�GME� b=�!B��x	����S����XKt������p�)��!�u�,�ߘ�
Uw	2�Ͼ�?w�*B��|M��O�Q����G����1q�� |�Deh���9�Tt��v��E$$؜�g@�iu>��#LAC��X�e���7t�D�D92u�W*}[`6�R5��r.h���h��)�!��݆�E�/Lj����w�9��	7p-�kT#�4�֣��c���A���0vj�%ΐX�l)M`'ụz��^����EW�E6�h��^j5+��A|��x�W���?�ͧ����x�=K�x)8�Ĩ�E�Bf3�!�p��]�}\_�[�4��
�ªl&\�3�AG�^Bk���7����(E��wZ���x��q� ͬ5�Zs�%#����V�%j9�b��&�tX���rMJ=gA�#�)�醈�?����u2�(����<����5Wn�K��w�޽%�\�������8�s�F���+{	�8��s����뾮�˽ӣ$"����,5;;<��h���5�b3�ةh.|hGAj�Q�B;c)�n��R�z썫�F�3<�ٴ�{��=���,�\HU�KG�h0�E�U&��NL[��{J �Ql�A�L�&�j�r���Hи�F���>�X	[H~h)f�B�9�I������kF����"���T��q��O�"TC�4Ag�]�Ӫv�$�x�矊��ᮖF`�*[;mu�`C�e�A��4]3~z�f�K������/�څ�ӊ��7`ν%����������]�q�����뇯K�tD74%�6h�����1��>�u�M��j�¶6�x#������H@�m$�;���'	�b���W"C`�r��Ȋ7hJG����jߘ���Q�ĻDO˭�@&�{~5�.����4A�e�g�w="^.@�m��ɡ0w�-��.���Yur;Ɖ����Z��w{fE%�$�L��*�-$<��&����.-/������%���C
�+6�Ɍ�+|G�׵���(�K�<������(.|�ʚ-޹�&�:�?A��<�ۿ��2��^����k��(;�]K���(+e��"��q26�Ygep�VЈ�(�D��S l����H�A��΃,@Nt��AL]��gѮk%�;�3MfcV#|�r$�� 2��㒟x�x6D�+�^������hs��ҡ8߰���zi%w��fTxaL+�ď�Y�uy�F3��j�D����֥X:գ ���0'�iW�\(���/o:\����	W��z�`��
���u��
}�LA�:N\S�8�M:������������Q،�4'��!"�ICW��ՈsZ7�/�0]�.������Y��~x�A�{���τI(3O��1�+za�^��fU�5i��T͂ȝ͇�@�p�p���F���V��!�6C�6_$\S���-�W� ����>y�M�/�����S�^� s@Ge@���<&�n ��(e���S,�b��� 	���
71vŭ0��դr�?y����b7�ˆ=K ��p�C�L"����m(Jqε~��0�u_ؒ��.�u�Ǿ	F��2|~�W�9���-��+�a��)/�uT����ͮ5���%PV�D��K��R�O�����MK�[��2���.��5Gp���q"ן{�M�Cw�钭Lqެvʕhb*%<����y�NI�3�w�������|2�"Y�|�WR�X��m2�9���/�#l�������`?\;��Vd�M7�ޞ��We� ������I榙"Mb�)�}Qg_TU����M�	dn���fTM���c�yoR#^z8Vf��}ڳ�2�V�d�B���"�B
��h<y���#�5�L�*ر�P�
�R�C�)ӂ���Z
~��Fx0,�a�Z�s	�H��[���1�c��qҏ2:�h��f�:q�)��ּ��������B�*�b�2���.v1ڛ���)��>i�;�]i0�{�TR/�%����5�*T��Ջ��is��Q�1q2$�?'�L���&��'4�]�)x��uY4��R>�q�,K�3�	�iB^�/�����:�G�iK]�����`�y��F�����!q0F�Q�]�To��
��H�p\�XAj���� O�� <�����/�+*����&U0%ʆX�8�,Q�u����D+6A"h����s}O��(b 1���4�m6��U�M�˽��h�i��{��Q��|�͍W� �L��@�+4U��F�b;����ݰ��&=��}8��Z|c-0���+h��9�-<�"�I/������%��q��ӌar ��/��q�;�5R�y�e�M�\m�D�=����t4m�S#j�;[1�����X�����;���a�K���ͥ���������6��6�g1�D��۫{<����K�t������xV��w1%]BI��녜)��M���c���;Y�Yl�<���5�O�6>�qM��e���*��ϲ�Jr�>�[m
=�f��@i���j � �_��X���`��_�CG���*�u����<@�Gpw�s�"r�:�ۖ�Q�]�}���$d�|�[�*�h�L�V�Þ�#����ҥ$A�06�� �*_�t�q&�f�
/v�$HM���"t^ά�-�	�5������p߰��`��L��!�cɓ����%%�t���1چ��Z6,����ʥ�4��E�*�)o�`���E ���^��*ߋ��[�rO�y�g��1�� `������b^DG-
�S�E~���%�I�z0�G�q=]��5*�L����=wE\KS�譆)�]I#�H����+�d闊����lS���5���+�x�|�9��@���<�t #��Ύ���}�����.���*/(l��҇����h�>��է!++Kr�u����3\&U��:��,^����p�%Q?��/k�l��D�@4@�t^��(�8�Ӧ��H΁ސ�2A���h�}������rF�)tDКy�%����� �!u���ɐ���EsQu�F�QX��{H�S��c��⢍�2�zM��;>ͅշܿ�3����]ȟDC?����e���� �f@�@���u�=n����ĩ�Lj���_8B�H~���2��讋,�"j�w1��w^�v�t�w%���J	(����F�L�ܣ����������v�~�]yf��!��6Oyl]�~�_Tx�`��5�h�P1�Aڪf��a�����)P��>��X��W�큆��`��5�}��0b��T��ٙ����q��\���k�:�N/!M���"p g�3Ռ5��F����	Q4� �!kb`!+e�.�BP%YPDA���Eu2&�V�����}�1D�X=���Gk��&���MlG�^GØ�G�'%�����^_ٰ�y?�����])'i`y9�12߷�B1�y	�l�wI�shN�pT'{�1��Ӝ�C�uOt��r"�&�' `�o<���U���=l�� �V^�)�/c��N`�l\��
]��E�1]53�K��ɲ��(����L<�ex��Jx�G�f��a.Vo`M��L{��� J� ����FC��^= ��}�cր�}tr���&���oO����Һ��(�*vc����H�:��}C�g$��s��''z|=G�g��@��#-�����p��xQ3;�%���V	��K�<r�|����']��B?����Gq�d�W�r�(l^��	���S9�)La�g�;�Gf<F��*%������M��B���Y����?H�i�u���W��S�!zo�T�~՟!�E	���h��$H� �υ�W������G��Ш���&�V�zz`�P�0m��C�)K�J�5��sm����y���Qc���Ro��Ϗ�`��4��&�������T�@�X�"AJ�첻Lj��Dg�����|���ʑ)m�-įv9ч�<f_)�e�0toW^��H��E�U�H�^�Y��ƒČ�N��g����6�����o7��].����2Jo6.������f4�t���J�s�>�Mf2|����ƽN�kv覷�P`=s�K� ��.	djG�;6>�Ǧ*�s�*��6m=S%{�~>��H9�5t����({�rui/R4��D*�`w�����:L|�G+�o�Ģ�,���"0�>`�$���V9a3h���w�厯f鋔+S��z�S�*=��1GR�8]��W��5��g벿8�|'Lf�H'�M�S���(k=y�p�C��6
��msG.fb^�oyW�4��aZCT��[6���0a래���:$��"���7�af���;/ԣ�P�#��p�$H�C�J��W7w�o���C�5r��h�]�#4؊L`�D�ԑ�?�g�� �	�KjV�緩��*������|�Bt��+����G��C��9���Sx�$R�[�l���<��l�RT��<�Nۿ
ՓipޮiY���Mivj�ȵ��1�6X��`G�Yc�@��3��;!��O��6/��ep嚴<�c� �EmA��<��,$�~�I�F�����1�+5�YJ�LF��M��$�!1��{��tr)�ir_�qN���ڵ��ܱ��%�.	˪��
�h�� ���P�쏣�o5	��N��ίP�x*�6�V�g��`$�2�M�*�q���������J�컪p4��2I����K�m�*��v��u_F[a�0ܥt�ӗa}��&ء�kNه{�y��h�����K��xIyCTo�F֓�σ
<�yw>A���;�
���y�#!��ړ|�p�Ϊ*L�
�r׾���Ym�7��^�Z�Z��Z��q�.E��P, �V�^��_"g���^sq��Ǵ���$�vu�����9�{�u�1C-]��%�P`r���=��t^�0,�)7o�B:�Em�s��JG��j����O��WUS�������O��{(D��]G�������V(�fy�nea�w'��n..>�<����/��� E̟3��I���lQ�nؓ��-��M�t6���xeu�#�sߧ�wA��
(��X�"���i�Z���9M�7�ܐ�E����\�=p�m��v"`0 �>��A�p+y6����7��P���Q�dn�3�D4@���u$�q���Z���r�$���n�:^վ C��e��		V9��6B��W�"�jF���|RDͣ~?T0�����:㧐��뒄�~n|N�X���ͩ�񻊝�G����=�����w�A?P�FEŜ�t�@�����d���cJ<<�0D.�������t��
�� }ߩ�<w��t��0%b��[=��GD>���y�^N�����#�?�!������oS�P�w��z�7���2� ��D�솋'���ٮ�?�GZ%��H14�O����
�l�{߯�๜��Om�"NKsΟ�ъ0���#S�$�1	�˩�ny�f�Lc#骲�=�P�J��#��(�^HMf���C��X���,��»6��Wd�b1���&�C��{��� ��,%�0�� ���)�M:hc׻v��-M2�&�n�P��d߆�;��oP��A���_�z��ȸ\���������gT%Rŝ���y���vc$�>���"ѿ�S��Y<���F�����t�ߏ���t9B ���Y$�@�Cro�݃�7�ef�N����b;�y�`�P'��/X��Pw�3��(i�u�&��GXT#%����85�H�?X�n�	�m�W��	E��z�%�E�̽��F�;i5ԗB�wxt���2ƫ�$����\��t��0ah ��T���Jv�(n��u�q'���� ���
=86��LHb�4�Y	�q��X�H'@h(��H��6�-��	�˭�i�s�#XA�L.�����m7l3�s]�Fp��.��{wDLe�W ���t�������*�O�|H��e1�3��tu��+t���8�0z?䡲�流@���n���2`:��I�Ǧ�h��TQaL�t
��u�!|α_:�q�>�����5��/#�20���?�c�cAݲ���H��������B�܌q�{�{��>Y���+�j`����J��wt4~�m+���W����rU7�8���k�q��=Z��\����I���z	* ջ��㕓p�v4�#aw�6l�5����h/�;�
)"7q�>E݊>'��޺X����߉����3Nx�L �.Ua�m������Lm2yvT���9T_=w�f�?�P����k�Oa� �Z���P(�X-�:z��K;bF�$ ��'e�I��n���.��qH�)I�:�#少%«���uH��,2̂r��5�)4�V����i���;��Ҁ�K(�*�.���;ʸl�s�c���(���Ԙ���/&�H\������������}D��x�]b���	Eǧ�,2pԧF��Mj��,�`�YK��74�M�܌KP�t�		j��	Ǔ��*�A�,�mp���%J<�6�.���:W�e��d�;[^����鲑p���Q@˭�7+7�;l"�g�{<���KuqRe�Û2���7��cE�}ނ�O�t��ƪ�.���}�׼�Q=���Wa���G�0{����}T7��]>c5��O8;B�テ�d��:��y�u�~>`�Ń�����\�c�@�闘&��
�i����h�L���{1��ߊ9|3U�!Y��p���ů��=����:Wts\We�S�m���d���?���r�֡ld*�@��x��P����y�F��N	ʬ�O|�����ǭ�T�?�����-1o&I��`�$����:�ԫ�F�u��A+$�xm{�8Z؝Ϣ8-�i�f�&��&�.�=���>Y����b�Y�)2�X���t62h�3O5U�S�s��Z��W3򿦨�щm�}
����El��L9�a�m#��X�ޡ����t=��.'T��HO-�3�7O#��5�mf�4��U8߾!_�jO0�`��Ln��u%�P��s��
H�N%��؉O��0�>}@�ۯJ���Y�u2���Z��T7��M�:���Y����s���s�a�#k $��@��G�'b��I����f����ˎdڧ����zG�h�)Ƙ�9��9�Y0nT\�����^/I����sĴQf�}jc�"�q;	��l�"�M����֕��#e��J��&�x�F����Iї���"��9��$\�jx�d��&쏮p �X�f=3�9Հ�ES�`x^�p�2>3r[���{��UƝ�*/h�Q���1y!,��}�1M��n���Y~��$���Y�u:�2�-H������D��b����������O�ń�Yn�i�:�>�I1EqYnй'�/���n2�pd�F~p�oB���Ợ��%Ң��0�J�K��>Y��,1�������ڌ��'����8u��t�fDQ��&��$2��u%��8�f_�S���O��h�H/� 60�x\�;��#�U*xe�X�䴨�y�nk�-��eF����7�&�SJ����ྚ�݄V^��(%Sr�O�lz��k�� �5��B]B�4s �Z)�߶"�qp�AO��ͧA�����*�����11�U<�=�T$�ut�T:���s||0�&�,�ʞ��hyM��R�}�lz���:�G��G��!�e\[�{���v��M�*)`75v:p���ɔ���H��V�C�UX�3�?����.��ʱ>q݀&B�eL5R��X��:�����;���A{Z�9u�D�Ɂ �����t�%��O%Gb��ԏ��v]�!����DͿgf�/��G�x���v���_EP��t��CW���Z9?ȏ���e�p̺�he)W������&�yJM����f�z�3�m�-��T�$�(?�a4l�F�È���*Z�#���R"�5i�΢*�'Y��
�E��{J���8]���Ǎ�Nצ#l��\g�����{�II��
�e�:v�&����o�Pj��㮏�mQ �
�>\+ȉ�f*�P�f���A�nG�.������)E��)�܍������M|�H�{/��KIM��vf2����%ؕb��0!7{Y2��&p�j�C1"�c�[�+9�}'HZ� �"pz�M_B;�6���[��z���c�3N�O
�R+s&]9���I����� ��E�9bg��#2��a�����ڇȳdf�,RZ� �ӟY@<��4ިo���w��]�A�~���Ky��l���SoE��CJT	Y"#Y�-���N�Kx��)ō	*��f}����_�$s�ئ�. �,���l�D4mt5]4Չ7��%~�q[$��9���E���e�lnH�N����俒����c����8�����1.�ֆ�,�)�&��Ҷ�]�+����Zl�4�"/Ɇ�����)U�����ot�������|<й=��v)�qg1$F7�x=�0�-���6�����htA� ,7��.I�+��"Hh�Q���`���{�g����!��=��o�k��|l���5Gg��";�6�	�J��ȸ�G�~iA�����ud���Ur���;#je"r.�	b��f��"�Ih!z���L�Q������ApX:��s�2��9�[}Q�#�Sin�G������N�7��r�ğIk7U"��r��
�����fb�Z�鹵��q^���k?�`�&�uS?oi�wR�mVhy�{z
鵺L,W��I�+͂w'Q"u �����1�J�b�FZJ�`x���;���{=?D^��[�PN7:3b���%b*�(��ZTXf�n�m�@,E�p����{M��u��]�^ò�����3uu�ot�=eN��x�7˓�V�����PC��$�������N
�LM�,���A��*Wdͨ��w�O���E/lq%\؁���a��!C+M��ń�% t�g���.��w�%����v�ݭ9���G�B��u]@�D�;�4b׮F^=hx�_�p�_£a�NAk��?1x:o�wmw"����a�
TUg T@Gx�3-%H����b�D4i����b�t��΍�N�U7�SH)����X�v"=r=8�<�̾�FG�����a)Nt�Zŷ�H_�0�x��p�%�o���?��}~s)s���p�gk�a��Ũ�ͺF)Z��lM J�S��5<z�˞-���3���7>�RN�hUc���n|b͕ɒ7��������-��.~�%��)�g1��v��q�#�=׆Z�{��7�t�"���=sb\���G6�]���j�	�l�^��-TdoW�3'�I3Vov���O�����8-!p.�J����5AjG��AR�Ԓ��B��}��n����i��Vw)?=;�|UP������.Wl�2��hJoK!�e�,9C!��㥯�^j�{��`�^I�?�q�bWk$7P��7Iv^��;�z∯ܹ�eg�Xb�G�N��׮S�v�	����������,�L������q:�J�^N��ũ�v��y|����-��۰��W
�'D��w���@��غ��ܝ�9�B�HW\:�Vv[
��e�������h�sc�~��gE�d�:��w��9!��goѷs��}��`�\���r�č����2�r��s�i���7�l�}'묛���6kt|4��@֢$����)&�Ջ��^vi)��1r�z�d���A�'-A$ͦ�|4{V&L��Z�I���v�%���׆�A^�-�ũ�ܨ;�:0��{��u@�j����C"&����i_d��)��)���&oQxV�O2�X����Y{��j��¶^�:~����Q��uP^5Xl����l��E�ꩱ}r�0��w�eW?a���G]"����@���*�PN���ɷ��s|aRV��<?{ꕪh1�2x� 5˗�W�1iL���0���2��ʜ���g�'�}u:�v�2�j.�E^�v�5D9�Nj������R�|�$�t�6�i�E�L�q�s=^~�K�X���%3
�&{��݅7C�ќ܀t�H��,@��a�I7f�:4�&q���H"���i�3�(Y��@dp+����l;Tl����p������P��f��Ǌyru���H|��
��"��J��k�T	K���̷����<��T6��@E���ư�iqЖ��o��֡v��!#�R+.F�D�C��F0$�JCȻ���;W��&�d���kad��e���V	�u�^��i��M�!�¼ƨ�1tN6�m����3_���#�+aM� �����6B�o�G�ݥ@��)s��!��i#�z-��~GR���0���;��.��;.��Fl��Sɛ��'ɀ��##_Dmz�N{�7;�m��s�`a�槙��SvO�&Ւ@�k;�� {4��y��4�	��2p��-.�˹T19@��:GZ������t������ ~ɔF&̒��S=�����״�S?f|k�˧;ʂ�=�B�_Q&��fph���إS=E�=)�ޑso�]~q����$�ߓɨ�Sg=�Ԇ�A|�G�A�����nk�xۈ g(�S=3�!E�z�*��I�;�۹A0B���±���	6-~I�`�C�\�
�����?p��ش������N��n�{��кx6��M�^�L�N�)߼��`�`c���e�[^R��S%@mӻ���'q8�H�^.7��#�S��vY�������R���9���yK�a��j�����\�+�G�͛�Ǥz4T,�yl����l��J�Mɺ_�,��P��	���K����!6(%Ϝ����+�Y�:'�h��yF,�#��.o�,&:�VpR>�N�xլ�<S��E{��"Ɓ�\�s�ݼ��h��6�\:p�x��c8��,���Ww�]��qT�gA� 4~3ܵ��Uk����5f%J�ޢ*ӹ�#5[B����9�bbk�G%�	�!o�H5��7�w�ڭ��-�q�{竄�Þ���T�jWs�WKx��>�q�nfU"��F�	��s,�b��2�f�ִW�:�#d�� �"y1xNr���#)�]�2�"H^P�N��wYO���^0ÕI��gAH�uni���P���E��H4���a�Cj$�? ^�VƄ6V�3��k]�J�&�)p	�ct=5n�8��m�t�8G���o@8��^E]*x���V���T�T��5��dnm �U�O���zۑ�}����t��B�:2���E��1��h�g�v[SB�n�"_�K1����`Lcn�3�E�FU4EJ㭮�����)���p��1��GZn ������ȭBZط�.��nP艨�J���Y|Y�i�@ ��b�a���Ox�����~�x��:�����뎠U:g�|5j���Oh24�0��g��a�~py>�6c�N��G�Wk��Ǝ�p���_Sf�teS!�m�|�dT��2���Cq�C܉d���U�<������ͥ�m���N�S� �-��lw�V(����au�U�9��o��[�g��R`:�Ң��b�o{�A��ʰ�����?��~ɋ`��а����.��:t�S� ':��MǍ#�ͳ��#R�ԏFҸQ=�3A���9xj�8*�ٷ��ڰ��To0Nd�*ds��%����;�HTfH��9c�Uv��h���?��T��5��l.�8UU˗-���I/	7u?�'�Z�	~�'��?q��S��Z��g�B�O�i�/%��,-4h����)A����e0�urf:�����v���|�B�����]'�����DY��eO*砙�Wk���m���"!�{ʵW�����)�������2c[y��"}'٩j�Xj�q-�C�7�*�z�Bz�d�������ɯOC<[KzI���F��HP⍟Ӡ#�Ԟ���G�������bxJ�\<]jz�'��EDm�-��g�,��p���@��|�ʮE�XM�7��0�i2[%��%���]0m��vX���!��M��<��w-?5>Q>0�#x��=0G�?��L�|F;y����������Jj��,������Hp���4�Q���G�<�ӎ���({Z�E�uq�H-��+�4�o��r�"S��P-�f���l�r(�H��6����+�L���<	dM]j,>��U�p{+��(!�d5�A	��*�\-�d̘i�i}9��"zڠ6x׶˽��^����o�J��iFE���������/&#%�����s���?%xx�%�-}U��E��"�r�Xy"?���GV��TmLO&��~Z�T��s�.�&4b���Ax�ՙ¥����9���J	P�|�a�ñ���j}6&ܽ�I@H������V������`1�օ��ξߕ���ڷoi1���������ߥ�%`�	�Q[DX��x�?I�N���Y�Pc� �#H��؂>��Y��8��(�&�Ԙ���Y�Sw-57���4#���YA�W]V��DB`*?Y����s�
O�8 $/�a��L =��whn`�_
vm�5k��N�p(����7B1�duk�k���x��^�͏`$w��+�=Ж�q� ��P���c���#��I[�!/D�$%<�1B�Z����@�!,�ag�G�N �ތ�������(Ռ$�YWjCq��n��Py����M%��*��H�z���x�g�A�S�(��
\�^�yU���^�[t�0�������l��V ެ���uj�gNB:y�%����4��#���/����:���z�Sﱢ�=R�ߐ�y�_�-<���fX�G�b0�f��ia�Ur�5�{���=��94rî�r��I8�q��m$���$E-�m	1��7����1x_.���mܓ���M�W���l 6��'p��h�Ϋ+H������v�K�mfj�Xu	�|,�B���k��B
>Ig�M]�s`�:��
W���Z$x韒��XӟĬo��bw���훿Ә,�Y��tߟA��,6�|�J%wmbK9�h���F �w/���b��0n��Fy���Z��k�o�!|;��T�W�9�q:��-��E��f6D3'5�"@I�!H���bͪ8�7��'�;٨L�|.��tċH$�t� Ǳ,ď�eJ7�S�6D
Sb˼�������h�f)���7_K,�
QvG��Gh�������2��!��-��N Y�9�+�V�}E��D��:÷9��p�����L��K-��ףz��-vMV��~	�;��$���r�R�*d��D�#4%[�6��ʏA K�=�l$�_��xI�k�D;���\3$w��(��R�̚Q��.�#?�|O�����k�Id�Ybpgv��A�+�+��2�e�U#���b`�������
e����K��|-�T�+wI��k�o�frD�#G�5�)�<�fL��o��-�Ag����&8M��
���ż��f]
l�n��	��o�l���˫���� �6W<Jd���.N��G�-�K;M�Hϥ���I���:�e�[�G���$��␑'M�f��|:�K�T
�������H��-��Zp:��~ws-)n$1�!��J����m�'3G <x����r�~�����%��t)A���A�I��{�۪]ɩ�&�����֭c��<��4�&7!JXes�2�b5M�T�_y���LAI f0��讶(���o�eF(���pP`yI���q(}1<Ŕ���'ɈJvv�I�Y��񷢎v����_�|,q�S\�}�^�6]	�dK?0%[,��qE�ݶ�7�+�5���O�Qc�F���ʮwz���ӮH ~��LG��Ю��T�����Df�������
�t6s.Ǩ�=lV���Ai۳Nh��n�<��>@�Ϙbi򈃇�&]��7����>��K,|���~.7�D)���E�U���4mGv�����	�&�I�+��V�i3S:�2d����Π�X�U�� �?)��>�*��ITk����w�kl�E:�n�vŚ\;eP�^
�sC���.yLߤ�2�@p�S��J��-�RP��2�O���D�.o����VUM�N�X�pc�AZ�b,�8,窳8�Ij�S6Z���C��D6H6���'�w?�sb������� k�>� S����#r� ��~c�"�\=�����)�d
@� �ܭ��>����)�R��<��z�
�~���X�|5��z��;�P��nA����[�.�=g���l_��<6w?��k��ڽ,-f�@|D�z(�!�J0:#�K,�Rc�M3�� �Ӫ�O�p����UF[�7� �תƪ���	<j-(]�bK�R�t��L�Q�#w�P�\)iBT�g�I^U��R��*�AC`à_k�����&)��霊1(�V�<Z�A&��%7��W��נ��Y��@m�����a�c5k�cɚPA�:�X�\WFr��w��7�z�"n�����SY]P+��e��r"``k�zj� ����Hg��O�!����R�}#��0BPAfZ�����{�pָx��B�΁����Hǵe��5= |c�7>�o��2ŀ%{��+�em�D�T\�x5Aj>���c�:�3��+�>z��a�_7��� ��Dc3h|!�"�v8\Y���~����"�z�#G���j�=>��fn����<N��Z��-;ۂ�ݺM���FM3�r�,��b�},����(���.�6 K���X�n>��-)��ᇑ�e�N���
�Ϝ��� ��f�r���l��B�4���J�E>No2�η����]��J�����f�*�����-�ɇ˩J��nC�!~�l�}5��n��?0/�9�p?��z嫪U�W}��A��b=K[0�s��B3��!�����CG`Y��ҟ4+y[�o�J�>é�TA�1M�J��)�/��	�bv�^�j��NjZ����[2FĐ�Bp�\1�<���-&�A�7k֏d V� 6�$7׵C�:��F�F�_�Z.���{�P��Q'��. �!�:����w�+VV_�Z��#c��r53>�y���tv�����������UO���J�N�Ks���f�X�@{qty��+9H�L6Zd��_�\J��t^j�w\d�Jú�݄,�^�eG�:o��s�>���n�M ���.�vhc��Ll��ٓs<�t}�-H�;#p���l�)4��ϥ��h�ʓ�\((�����!%�oy����R����P�6���\����7@�;lgЛv�M��ā9����K�~�.�n7ztn	�C�g�����"�8G�)p�S�PFsg��濤F�r�C2��%�0g��O�s܆�.���LQ"��A�4��bb��}���)�^%Yo r�����<tӭ"P�_��L��\�L��{� �U�u�b, 5��0P��O��)u��̉&�~����X<�݀7T^u���&�V��~B�S,#��5�q*�ψ/����엿l*/��\J��9�6M2��}T����MתaY�!�!�0%u�'����{��a�Ad��{��p�RKd}�ޚ�ұiߪS�ס�m���Y��<�\M�x��SX��%�A��W�����D�m�{���v�A2G� �6�Tu�E�V�>~3�l*�Fk_kH������(|S�xB/Q��%E/��Z!�DV�:j8���� 5�Ƞ�x�|��8p.kksr4�^����vT�&>�;��N�4��0���rd�
C5��xW�UK��P�	�s���{Sh���4w��k0���Ll4�[�.�.B�h73�\���Z�R`掩a?�=˨s���,j�.��{Q�+���ok�mj � 2+��������P��l#1	ۑ�1�o����e[7jĩ��Y	u����6�Q��U�����i��:�	t�� ����#oj����V�JꞀ��ۡ�ۄU�<���ޕ�4�d���^b�a ����ֲ�gz2F��n|�:�d�=R����ddW��Q9�6�I�N�S1᳛Gi�6T��r��`��0d�O�
m��m?�MϢ��쪝���s,�.�[�����~[��Gt�wB�S^�&f֓�~u��Ez�aI����$�;,Dė����+\�0]
�[����`F�����b���J� �<��.����B���7h�%�1���|p2x$	��O�m]ԏCӻ��z�3<�V�{n�t^�x���V�I��J���iտ,]��"s�,Q�D��a��}� �7�h��������Zb������h/sz��`�J��b��W���^�G=�m�f?�u�B>�i�?�ӌ�1N���XSQ����nc�����bY#������`����N���E�� пI\���U�ܒO$&s�`�Ŀ�i �t��V`eC�bA�d~����=d�Uػ�q�Z�)����>�'}����W�i�6�&��T�f"
63���h����b������Я9>0����ǂ�/&!f�Q��d����-�6��j�9H�6��d#��Ynƹ=fx���>��uI��@ۏO��T��}��p'St�1 �s�D��K�,�ɻ�0/�����X�\�gI�@�� MxVT�^c˯�
yq��-����Iy
�_�g�9K�,��tw<\�\�>��F�Ni��H�^��c��х	c_���8y)���������!���ɵ���aw|��w�	S耱U�eǹX�,����=��`8�t�@��ʜ��nT 7�+��f����V��:�����Y���	T��;�^A˾��
7Ʋ�8P&�L�:_z�bȄ`EL�Q�H�Ax�21EL�u��Id�	��yf��w��n�7$1�f�'O¦��y��� A���L�q�|÷��a~:��~����Uif�j��`�f �����6��c��mCcΑ'�o��j9�m�c����l����D)��&���1�mS�O�8�(z]�"��
vf��5W���a4킷�mz��&4<kHe�e�����!h�C��s@��(���l�ʑ'���:����.B
�p�"�s� ���SDO�r΀U��p˿a#XX�И� -���Ǉ^!I;՚R{�ָ�Ӯ��yDE��KK`bWxym�^1;^*����%Z�>�_a��Yl.[{b���*�`�������K�f	�@��R��*J�"�d��I�&���a�����K���#�I�uHЫժ��qT�T�W�i����ك��J�IY7A��p�I�9�g����k�jaD�*�i� I���jk��wW�M"���~?#1���g�� ���x�|��v��'񝴅cN���OA�P�����<Mf���C��ar�ܶP�)���(.~�\�!)�Ѡ}Ϸu-��i�*����������lW���CjU\(�"��{C�9�d��2%>���!-�����#Ց$�zV�E���s�s"�~@-I�R���%�u2!�a�v��(Ov����'@��&?�F��m�K2��h�ZE"B$B��� RΖ��v͝���f�X[5v�9�x�z<����J ����2�ZO0Է>g����NO�Wd��v���5BpW�%�:t�H�9cS#xZ��nX��Q��W�ric��|3��8KJ��R�,�Z̽W)Ί���D�\�Tai��,Z�Кˎ>p��Y�?�4��Y���L��Eܿ���Sz��Diȶ
���zݑ=M�Gx��be�V��[���o�]	���z/~T������j���ǈ�G9�q�����0��}�f,���<_�?h�J?T�0Zlju_�Z�PߵM^g�C�7O-b��eE֖�8�%�;���x����	����򜬫�t��󶃺��MDk�����7N�ч��>/I���8p���g������ˬ��n�׶�x]}<�������٢^�c��p3�b:�#���<�>^������g�!>PE;>;��u}Z;vǵbFK�����g�=@�E�x]�p3��X�V�C���|�d2P�pO��q�E�� CL�{�z��RDdpS}��M�|��8P�+��赩H�q���Vv\�݋�圮�l6I>K?U*}��H��(���/D�![&���3#3a��yQV���0Y1�뮲Ei�ʇ9	K��%x^��"��<�vPZkG%>H�O$�h��<�����w�/��(hY[����@p����Po�4�M)�K�ʿ^�tH&�V
���֥�>v�zgנ�Sg�U�]-moJ�]fr1���lY�'�,=�T���6����ҏ��e�M��!#0���`����,`��0H0��+3�����4��>S\��r�b7��yJmR��uG���X8�f��r<x	#�!I(��J9��#��Sy%�@�����������kt8��Z>�teK4� 4�,�d#w������E�B���z4��L�@�t`�֊��Q[�� �Pǘ�����a����ߏ�.����=�Ys{_����#��_��@�O��M]�V;�
�(�e!&v$ߘa5P��S�̂�<�!d��d��:���+@���l�̣7�?��?�|����>(ᖴf�٭�j�,`���;,��I� ���J<�l�v�#���1�'XT�7��:W��mA�;5S�����=�"�ŭ�\ex�:�&�@�M��BE����d�2��yݠѵ �Zls5o��I�.�i�cS���~2�'B����j 7/�϶��a芑#��c╼��Lr2(��Rz�7j&���z�Y�p��BDs��}�}R��4a}�qH��˾~=/��S��gy@�#V���傺Е�"���y��E�b��?`/��������"�V�[�Vc;��/�^{�eI�V�M�T�$^���s@]�w<��ZE�
�0b���jP*�M����RT����(8C������gޙ>�~ءCހ���cZ���7��T�`T[�+��������)r�FR�;���!z�@���X)�L�be���n	��Y�*���%� 2�s�>���&I�A�0�6!L[l�H��*3��5.���JlT;lbf�5J������qA
P�y'���l��h{M;���qUH��v���4>���Xܱz�%<l��[�s��T�n�#ĺ�NE悉����6��ǳi�G�1Ы���
�
�#��|��ƹJ��uT��G��B�	3�3l4Sq�����G�q����1tШD>u����,��ozA�>X_mQ�!6a�B��07�H���:WŢ�D��ei��sGY�"#���},��^�i�K"��#;��0R��0&8���n�!�0.<��	��)�_B�
�Z�N��pmW��"aO�v�"��_@� l��;r��A��e���f���M�^I#�y���z���'�d��v�����R�����S)?7#��
wu�<�`/���E7�i?p9�F�~������(�Z�k;.��]{n_�Ir��6��d�ǉ��m�B1�1�����j7��\ד� ���I؎~��tTx�'t>1)�,�����+�A�8�4(d��H����,U�cbo���pkS�ep���BNj�+�ˠ�.�|��l?������9�3����1��|lJs�[�Q�Ȟ��#^`�����~�G����kA����4�=F�˖�p�N@ɣG�%�wRp��y\���&��DKB�7�;ڸ,]�� �V[r���^���#Ͼ��1�2Y� �f��$���H>=�Q�
fӿ�"�|��}s�����Cޚ�1q�h��q�<o��� Y�:�Ê,��&���D �1��Ur����� �k~2l��$�Q��!:�҉����1���xCz�ǻ�{�E<dD���9�\�y�%� �����gYG��T��^�2h��Il��Í��wGt�X��geGܒ�7e�׸�@�Zչ���?򚧴���:6@���=��S3�ԅ�9��@v�����K�*1�`6C���"�o7bgű�#K�M��a�f�rP�7N���5����<<h�|����oF�}�$	��߽~��n��-��^���2&K�"�On�0��u�C�ۇ�_����4�w�>�LX4\w�Hz��j-ZZm��X���ڕ��\~�hyE��bs��7n/HL��i���T E�*/�/���#�#F����K��紅VǶ
8He����W#�өR���T�-�sD�6�g)��@ ��}q�S-%X���ρ2 O�F�"�Z}�iČ�{Ee������'|)�p�n K7ܔ�Ă�ՓW���)�iEװ�����U� ��yT�F�m��u�m��р��=���q>�M�uc\�p�L�M��x����sƊ\�K+���I�T@׎���0�~�)���� k�#�t`�^W�}Z��3�k�$�}���V�����S��%d��g��9ӣ5��%T#��s��I�~V���3H�=x�IT鬓vQ_8}"V/[	u �MlAʈd��WkY���HK�TI}L�\�؁ǒ�VG�������=��*��>�n���;�๬�@2p���������h�[-2��pd��^��(?]�z���q��G�xX�jZr����� �w�Ɣ��}�$�ã��������i썒a��R�ѣ6^Ŷ�������iQ�T�v��0#eQ��� �d���tB�o���ҍsj�וN�t	G���z�.��
G����s�Kf��F1�U4+$G��z^��Ȳ�Ʒ^����ea�:���y���_��S-�+upb�:�����$xnm��	����2gf)T���KZ�� �Rn�y��b�{.�['�2jж�4<}��3�R(��Q��n��l��7���O�p�?	���_�C	��}@Y!�'���M�o���ߠ@R&�����؏q���A�]�gN.9��N�m	�6��m��	�n�b��k����e��[��+���"w_���ڷ�u��H�t��eφ����� Q�mk�.��p�~������pP	?�V_|�\��k�b�p�&�|H����^+�6Nt�lk���~Y2
}�����=O�AH�ײX���_�EF02�v��O�|)<ߚ���k^#*��3��y��\�f	�(�� �U]�����ڋ�1��0:�x���!���z�����Շ�^�'���gl!���y,2�#&l�Cda�Og?��-�N[���A۔��x�Ǹ�z��i�%� ��pZ���1`/�Q��ɂ��^1����e ~�wE�*��!�=$\��*���E�����E��HC�s����OJ.pXQ�ӊOZy�]����>G�8�.4���5�%x�G�Ńu�^x��7E~n:�W�6�5<�P�d6m'6X���v����ԕ�,P^�?���'�K:�{]���3i��Ϣ�a�<�n��2�aD���pR��
N8�(dzQ�)@��!��XD��1 �d���F<���� 2��& I'0ٖzW}������; �㾊�<4�3��Kz�E��.��=�.�2��y�\&"z�b�@� $uhA�s��"������-P,Z*��&�����,��~�N�W|ǄW�8� {ĈiX��W�Ӝ�<J�ɕledi")�Kic� s���CZ��15����HT��P�r�;�6|)zk �m�2ޮ�B��x����1R����>�vr�{7����'�B���	�5����o�$JT_zfOP�S�D�JP�����b�v)	�V�w �X�ˇ�C����T�#��;+ߐr���)N~��bX"�U�[QH��+v����㠜�WG���G�XM�=��7E����[q��ܝ�-���.��W�%�á�\�$����l��m0OiОnh�X�λ+-
g:P��c�2ݐ�Ǝ�AA�Pbm�H �%s7��!ٞ�Ȣ�YR	�$��eMrUϏ��M�}���e���1�̋�X'(�R s�g��H=�B�K���6]�p��x(J}��C�A�z�yº�������VH�H%�s�@�+hewuj�|w�S~v�_��d�
���Ӂ��&�TO�������}�u�<��ꆏ�u(>��n�ER{1�cx��+�����j�2��t4�]�X,����n&X�m\�P ��*O��;�]�'�w��E(|(� L��)1�:	� �|u�� ���>r���Hc��ݯ�����=����@�?y�v��@;��9��(i{� Yshl�9���{Q?`�E���p��}�w��h obp�!֢��xVK�_X&�e��|-�%��CA���1#:�͸aͲ� Q�"c	��̗N��WyY��L�^���t�2��6������OĞ�X��]AU5�}k��������E�蹽��1ߏ=J��g�w?!:���}�r��qo�y$1Tp����6�u���#	�O�b�Pz���H�����ٸ�Zґ9��e�#��>zs��#���f3,�Ha��dJ�ף%L_�Nm����{��%��F�[+K+l:C��j�?��A�z��4�n/=Kc�k�g�2s�l�.}7_DF�Q���s��v�����e-�l��L�����M	�WO��k)�(�%�7��h�A'��S?/���C(�� K���y�����b�L�Q��S�NTgݢ���y��-��|h�>�̯զ�Ǝ{�� �Hp��w��92UΥp�7�c5�^���F�-wS�d��l�v�]<
��Q>�X���ொ�Vq{���:��T
]0�K�e#.�z��O���ٛFpiܦC�	$�I�h����D�@���q]L箞�3 ����+�$�ҨT3=�D�sNA�xƤhd�?M�ȼ�����>c,�����(��#AWǁk���p�l��1��^�� %�gWx�w�8�Fl��Nb &�v��c!�5������gи�SL�KI_���?�E�xz�狔�
��%�G�fNŷ��������,tD�\���S����3��W��32�b�i��e]d���bS��aG�7��q���)�R����3��7�m�5�� :�5�88�gLp��^�؅���¿Frl+�B���$���A�~	�5c�XZ*�%4�=9�����<U�2�l�(���rH������Wլ=�q�Fc4.BJ\��fʤ��9�c �4���`Js�#y�jR~�j�?>����5�T aWp6ƥP/J-v4��U��7[�<m���d���Rf��~���_N*��L�:��=�d����Jn��W���;o2!�d��C�}�g���h�w҇�Q��+��VfrW�ξ�BBɃ����t�;}'j��$��K��q������>U&͵*��t�������8+�c4���<9r�^^z�+h�O�iY=��~&�;�z.q���q�u�����)H��s���|<�&�+�w��qۖ��_k�����.AŐerNJB�e��B@���k[����� ϸ#�v_�	Y��b���5�J��3g9�^��@P�D6��:�c�(<�Z�H�2�=.e��r,���>T-I�¶��a���B�����|�߼q�O#��}cߎ�X��@�������j�K6�
�Bd~���|�ݦi0@0o��*"�)�7�i�F��^F�ܞg�e@m�VQFOE�U�{���UJ�z�����$O�(�1�l:�%3�!��t	8NuJ�etmH:���#�)Ќ�ċF��Ą��������
�㘙hNW�6��8�ә�V�I���	^G�0�`���N��-'7yI����F8��ۜ��ZT~�Q����Ȗ�fP���ö)�I�y�{�uۋ����{�~�5	A%|6���[�+1� ����b��C��f�����!�:'��4kE�&����h��+�˫��~)M{hp�2[Z�(��*�N��R�U (i<�I=o� ��	�FϤH��c%L�~
�).�:�;DPPk�`7�ǅ@�b: {���C� �
�-RC4�����I�@(*�L>~aQ��[P�N-��X�� K���Uͮɏ�QsQ�0����e30�{^*�v2�
'�ٺ�g�yǱ˷N ���mtQMXǴ(�2u�����n%7~�=_e�٠��=W�~L��wX؞��w�Ɏ�p�H�h���fZZ�
�4�ÀhTP�%�j�p,�ω���xI�u�JZT~���܃+:���O�V)_Y��"�V�;D�S����^o<��j|�/z���ܪ��8-�z�^�qE3R� ^�F�roϟ//���'����Z��{[��H�f:(|8�?���Jw!�5� r�#�G�q��nj��n�D�:'��	ZnS� ���VBޥ%��9��p��b���`M)_Rc��m�=+��ԅ����1!��C3oI��-:�D'��4�����oY��K��bd��j������܏hMkb���;)Kґ �7�L�.�%A��alժ��8c�H���tj���{K��J�Щ��3���V��<�|����ơureEo߅BE�S�!��b�t�G���F|��!x�t\zj1��-�~ut^3@��k����`�Rwz�q�!%�ߐڶ����vv0!e�f�k��Z��/�W+�QJ���A>�f��
s�-�i[��m5����ri�OЖCy�ɷ����J������Got�I^CP����W�#���}%���t�
곦�˼���7�w#�^��T�할}�W*q�Hp0>U6�ĭ`5-�ۈ��˲�d�h�.Z,�FVrwD�i
W��O�ֆp=��`�ZqoO���>���ϻ��a�u�U?�U���vj�nm\���yP+23��ST����L�F��f���F�!����8^
�D�6�/��g��/�]�	\���Db���$R>����2���Swo�V_�@-��q����ŦȠ��u�.e�"p�<�Ռ9��Dp��F}3�I�@�=Eԇ��9�O�	2K��w���Ė�-(���\t�K��M�]�P�� �4��Zivǃ,D&v����[j�R�B��t�Y��hoq ��l!�[Bx�Ť"�?��1���%`���^ ̍��h0õ��)����1S�F_��/��|� �Z&Y�!V	����w�0m�v*1��(H���ϒcE��1�N�kߚU���	.#�"Y	s^���K�qmNg��ŏd���#Cc�ԉ0����Gɱb�7CBTe�������l�4ӿ���< >���o��A���m��R4�ޡ���1�Bt�<��L����}���|Z�֗m������3��vd�4r���nTH�(�D�(V�N�A���v��^��٨9���8�j�`�����:�埲p���-�y�'�Z�7*GAaE�#Ś2���F��x'c��7�I�+�pT��S�O�L�҂_g��\���i�O�E,��s�����^�X!�_:�q�|��5B!�3[���T9����J�N��`�Y�E�e�sZ`@�gY�?�:Nw�˗t7�D%n��U��e��R��-�W���h��o�G=����k��;��X�ٺ,�Y`KT���b�;R9{q>c1��ހ�{d���_j+f�O�1Rs�����o��5ٓ*#DM����p9��8R2�H?'���!�n�(Z4a�7em����<բ��*�~�PXg)?�Nj.9����f�-��;3�K���J���`�5	[��@�)����1���6���M瞝�!���~��{Hq7o�o���C9
�T%�����l�׺��%1��`u\�0?��T�\4i1��l����'!�~,����͘�NN�
Tw���ς�Q ��eɶ��'��.g��I�r�w��\m�����1�/jX���D�'���܏%X��r�N��&�mPb�V�~�3�P��!�x
t]����=����Ϝ�SP������k're�E�w;��m{{�	�twrz��ym�B�ftn)�{���P�X�o����1/���`v�7L^6ea���Nu9LJ;uҙ @�u��a�Tec̜3�c�&̈́�a�]�W�l��oK����p�v���?�4�w}ϧ��Z����u��.� e�޼��h�^��e��22�SbJg����^y}�<���9oGr����3������dƔ��2�v�8��82!����|���8�E�)�`��{����"L�B�d20�s�1!_�/�?MA�x��1�:�/o͑�-c�<�Z���;�|��F�y;�,�C��6�JL4�?G_7O�V��Wsz����
g�6qBԋ�l������]�̉����{����(-��� k���g[}�>�м�o'���;:��iخ��"��#��M�t%"�+�<㴧G4����+�f�E�X��.�xk���)[���!U����L��˷�<]4��K�y��t�����5�m1��%U� �EחY}�e����2p'����`�dfJ�'�6�A�-�2Dk`g������^/*]4�6h��	ܒ�`D�b(�)3q�3:��oN��@u[μƔ�2���*=�D_̫W<��f;o:�<�#̵u�8;OT5!��:�wx4:�Wa`wf ��cA /�(�!2�˃U$������XE%.��ӄ�n�]�?���c��Q:�zH�3��nd�i[,�E����{�;)����)\xS�IU<�,J*'�y՝�
7@W��s�2�)* y�i���3�7�I��������@��M;g�&�N�SBj�`�#�S���:b`\ 0_[�����;Q+(F� 0�"��;��79��/�����{W]9�C�1aGq�!��y�ƁL~C��k�/&���~0�zS�_�o%� Q����Mk݋�6r���`�w�.���1�W����$���Ul�������u��X�DPSʕ�.䑮N���lЂ`�����A<����B��hF�@��<{e[qY�m�Y�B�y4�o�LY�I��rݖ�^�Cܮނ���U�[4�!��TUp�2��I9�e��Q��i�ɸ�ăD���ڢ�ar���EO�(���D��*v��j��/(qO��G Ħ��c%�вJ��T���ٸ^ �d�����̺��~�mg��!X���s�#�~�?�m���L"�M=�zၠg�0������9c!���S:%�=�A߻��@�3$��繘��]x�C�v�j����6�-�m}A�盛��	�x��H�v�"�ph���yj�4��H��/�΀NJ�0v`GQM�9#Rc�|�[>���Ζ�!�'n�K���}�y��Cܭv����,�r����"������-A����(������*=�Lj�sm�NC/'���7[�����9p����	eC��aej��#u�̄lĬ�&���C�N
�5o�h}��;&>�z������ֈ"=����q)�s��2'����d+F��:3	�5#�Q������*�U}JF�ϸ9@����{s��(�]�����W�������9���RC����8]���Uޢ6���82���Wq~�����"�Lr��G 6���ZV�l�e(ڹ�k��&��F^v��z_�O��Ç��M_A����E��E�F V�p����l��oć��MY�5+�6s2Nk�W�4��.��2���\fy� C`�YNSJq�C���������u�A���o�1�fzf](-�'f�GB�׃HSj�L�a�p1j�@�/�S��2����Ś�u�F��~Vk=BFa��<%$�T7�?b=�~v�n�T�H��l��XV���g|w^$V�r��|ASF*�Qjs��Yn3�Jߡ	"��Пt��_�?���z 	6�;1�āy�%��Q�rF��g���u/U�AOj��iɠ��(&�)2r��G���y�}%{�t>S�j� ��] �wbJ�;.!������sjQ:��vYT"'a�I�J����i|]OV���������v���6��n��U_�rm���rHO�ĸ����o��/����[� ���T�cU�!>�ʗ==ÆȘR�U���)��cw�Ф�n���'
1�]F�0�ǰ�c�"y _so�
�RmZ|�f��r*���Z�;c�҇���l�P�rj��;hY�=��{��'��_��4\�`�8��9�&���"n^����	��R��.��3e�C�}g6j�~�ŏ���(,^�!��_�]���U�g�%�)\r(��Հ�ZOW�\�(���Oh��	G����P�]F��p"=E��<3�����Yuދ��#�O�V˃\���4���Bm����X)�Sr��4{GM�$��WG�y������G�գH��p��|��`��=_�c��'���B�en�A&�0>���آ.�1�r��ȗ!x�P��-^� J2t��%\�;n��x<�X�6�j�s���"u�}��A����g�f-.��|:��&����(!�����Z���XT�l/@���F�u,� ._�|jQLZ�K�ʖ� խ�-�z�s�Q��q�VJ֬�?���󛜕\;5�X��-+e�*آ�߾�����/}<]�1�z�$��k�+]��S:�9�Rp��6h��c�~��no�Q�wa���2Klm�N+�,��*���n�V.�ZFӳe!g�,6ژ��&ׂW�C~���HI�68�`�P-�nj��3�2�MJg���}���jƇ�!�.9s��L�&4Rmi�A�
ɓ�B�;Bu��y]T��n]k_8#T#j�E����;me���Hb�BЙ�z.�y"���<9�r>�1!,������YD�ɍ3���$��89ėn��V�7�P�j��,;�ڴ|���P(9��d桠d�f ��H?y9R�5j�vq��0�.<6����f��}�*�]:F���M��#<��>-�q/s!�T	�o�tM0{ӿ�)(eI����0�s��������Z�d��-�r��(�I.���7׸�0q
a;c��֑/�@�1_l��6�Q@��y�޼��������n $��'~�,�'ɉ>� ��J	���Z�v�)�@��(;�p��=K�-�x-����ުJ�g��ɦC�˂lj\�,�F:$�����upI�S�՝GP�sk���!�u�v�!Oڅ$k����q�g-�XD��M���;$��A�T������/5����x�'ϳ�;�Pi�6t�w)��ǆ8p��S���z�d�be�c�����A���Y����6B�-|X�o�a�S�rA�c����BRe5�È��V�]����'*�p�-8uq��QC��sW�����Q�Naq�oT�		�7J=99�"� n�R��[)8��۬YI~�2*|gJ�D��/֊T��X�7�LS����ԗ�m��P5�-g�/�����6ɾ�P�Fi���\D�0@éYXp݋��d`�y^��[i1����Jf�q���$U$�u�BP�&�lߪ��Af,��+�o(�6����)�DS�Wԇ9)|�&�跞&�x����n�ǎ:s�yF�B�xO�~(�� �`��+�=sƊ_�9��$c�Ή��� �Z��N�)�7��<��배��P�<ӈ��kGb�	��܀�;�)=?"����	�P�=x�[�I����}szb����!F���[9�H��u]�}�ZB8L���ݭ�Ӂ��۵�V��
hۛEa6���w�P����8�n;D�)1��p��HV��&�O��%-CƟ���������ܠ
X�p���ez4���A�Pw����v"`{�3�|��/��L��J{X��$�!G?bz��M�7����]��~�z�ρ�+`)����9��l�3'��x��[:ƥ!I�t�}3�$�7p����}j�����B��i��)��vOC�H<��*� B�V�5;]��jM��H5`� 2��	�=P��s+���KP?����z/}� L̩��|���T�*�U��%/"�;M���>�fye�-�|���%�b�͛�u�T�;p�w�L�:SHW]��q�:�X@�m	���Q�B\������:hZ�薧�%�g�>r1�����	��Ð���:/x�7e^hi��R�֠���A���S��1�K:���_T�ܥw��󲜃�ֽ�,�+��FsOu��"��%G��%��,���-�\�H��'�[VP�� ��\u�:?�0!��M�����|\�V:ar~��%]��@̮LWǘq�Z�WZxr�<��Е�P��8�J��]!��DG-��l���+��4&Mr��6$:��4��O�&n��x`BBY�7z���a�à�Ih�v|h��a���%FJs��C�Q��_nc��$.��BF@J�z=rW��>*��3�̱��a��/1H^���jsz�\F�<D���E^q�0D�����q�fĩ�-�o<�N�S�O�Fg������?P�\�r�8�m��F��쉅�C"9K�9Փ�]�I(�_�bL�F�$�X���	�H���J7ޗ�pvp�����~9����KR��۴���a�%G���mG5��������:��4QD$Hf���=iT�\c�>�V�z�,���Y�����C�.�V�H�+�P�� �Q௥J!�q��7���Ț�:���(��19[�����i���d��|�O�T\��JN� �i�eg](6BТ��@IK�5�@ZЊ+rm-k:��� W�ʤ�)�r�a��`k���m���SG6U��\x��� υ�&YC�������������-YHG�=Z�۳��?�]��\?��V��݇�z�/�~���Lχ�$�W���b���~�bz��PcDr�ę�r�ͮ�"�t�<�fƃ�#�S"�F}�)�������J �������0���&&ŧ|�c�N+\��U��k���A����JZPb8���"/_jxX꠽?��n��!%G�̀�L�5c���a�
���g��?�rG�$M5�Nw���&u��s
��iDA�HZ�$�+*a#�����2.�D��8��$�����${�aN�Χ�wM[�p�,�Dp��h<��G�.۱ؼ{�c� ��D�,3%.����4��P�p�����KX[�����lS2{n*돚^��$��s1<�����X�`Sv�I7d���I�-�Q�,Ju+��z�z��O��Si�3Z��uMB�����Γ�}>M.q'qQ��}�$'��N�,]��䷑��՛�Ǿ�+���3�cӜ|��ں�N�9[�)4U���g�>�ԊO0���zͲq���m�Tj�$LH��/�w!U��lg%�7�c�]G~0�)g�ig��-~}\�ϕ�8��+j1pOj���*D ��N< �3n�i�B�!!�m��W�\� ��WC4�������[��Z:���60N_��B�y7����iM�d7A9�9��V�e�.���'px�?W�n�X�d�C�(��g�}�*R=�%/3w�-מ1�3���Q�]����݈5d��9�4c_�$FC�g����S_,8�ڞ!0�6.m��VK�@ ���A�]����	��{��*欉��^9͞`Z�0~UOh�<��6I}�|ǉt��br�c��+�D�`�N{��D$șm�$p�%i.��ĝ
���6�3վVr��p"F҆���tDQ�$<[Y 1h�.˕VP�V�46D}=8g>b~�9�w�A� K&W	N��i��F[����z|{�/yT�oM΍�˨��E��Ԝ�w/�҉L`2\�Y���&��$VD'��8%I�(�X���#�7�O�*lG��ك2�z��6d(�^�#��ęiJ\�G̻b����޹쳂�d�p����^�UO�||j�>�f=��cp���a��4u�`���8��l�>(I=&���\��0:T�'��	��n��6�B�=��`�E*7�%�>���wJ�)��?�u9�tF�8�OuBh��D�N�S���������z�ERr��:��������P���~�S@�\��m)�+��=� +!�}�"o�yJ��"t�sCOcj���&��u���;ɽ��(�0�6�à�f�w��rP��V�迹�:wT�oG�����E���#�����:n�{�_�Djǯ�X��Y2-�Tn�����}%���W�6%�#����Uw������PDA�yظ��Z�;�K�(Y��@�baw��J�%f�B9�Nl���&`$�z����;�Ag�US?�ֳA����?��<_�gC����|ϑ�B�UG��!��s���&�y��E6/�+f�칡Nw4���m���b�eW��H\:�7�����iG����	+J-
�_w�)��.�L�����R����M�qn?�u�XS!�G�MpV����y�@i趛׼=�ISө�ݺ�A6���ĳ�/Zi�=ū�L�gm.�rAGT*K�#�5!����+>��Ru~�i2swF��2��'Q�`��v��������%����ve�|��w�6u_dF�yr�C�â���y#�*��~a��A�L�5v�(�$5�(-���Ku�w-]�].4�*���w�| ��:`�`�עw�q{��˺��s�A��,��Y�dؔ�ֱ�hϓx�h���I�B74U��;)�:i:0�F��MS�W��?�-Ԇ7� Hn!�� |�J��d�P�q��i�|�ι�(Z�K���+���!��S����:�rC&���H��q��kO�P�I��H�u,6��+C�)�Y��\}�[�^@pz[�%���x4�2 �Q����,����@�l�7���)�čajU�������GŪ<�7�n	�>X\���x��w���h�_���~Z�Q��k��"I.��ks�>
�5�O��yJ�7�&޹,>�7���j$&�^Y�����/0�PlƝa�����NУ-N#���w,�.7�do_���ǵ�=�J!3!�;-/<�
�X?xx��z�;fl޿�1GR�M�P����E1t�==7$;S�Y��_�C" (|�F��dn@���+Vr%�� B�cQ阻�E�w��Hr*?�O���8�T�d}d�c��3�*�U�����O%�6�r�׵Sa��m���!"�e�rQ���OMV�8��ա$�P��.N�����Aoq/�8�nu͓�����x7��퓨��c�9����c 7������X�>9E^D�aZ���E2w�rp��7X���s3H�W�Y�rz���b䋀��������'K��q�165N���L�an�6��V��M����k����UJ�JM1�&�y�fP��I.by��}k2���]7�#����V���z�sm[�6X]����'��p���q�j������6�GSͤ^+�/�L��JvNM��_���vYf"�j��ZW�q�Q� �|�D[X��ҿ|}	A`>Oq䀻�H�r��!`Cp��W1�_��Z(	���S��
��i��%k�^չ�����2+(u�n����㑬�'���L�q�i8j̑��������&�{X�zˏ��^9| ��sșn]���>�w�'ͳfh4��)
�iu�,�W{�"���J��ޡ ������Yaut�f;��[`��va�7���uc �Ƽx�Czi	�%���mCV�eF��C����Gy������
���BI�E������0�]������v4��83	�%����8a F&�2OM�����薠���~ƨ�1l�\e��0ઢ�i#�N�ի&Wq���Uq�U۟��3U�u5���L��|7�l�ؤo��A�f��\�od.Ύ�BI_���nk�5��;������~Qa�+uq���*�3��O���� [���p��>�<"��`>脼"v[��/�_#uy0(cCL���3�d��a�tԀ�Њ��8�?�"�i���ҴЀH��AV'��և͞y�Q���G�[�i�$!rmh�j���,҈<�s\z�쟃ʅ�gb�����i$<YǴ��2�$��p���gq��{G��^J����X�U��V�-��ma�!q���F]��)p�
�N�c�/��O�v�>���*R�J?H�����W�8�yyU��i���-�u�뭅��5Hj���/n�.TO��B/��a>&��w_��c�v�Xl���ΧKI+�i��sb��u��(Z�]�I�p�ƛ{���o�F�:��!��z�:8�3��/�[0����9(U��%s��	۟c���m��� i�hW
����(ĭy�5�+n���_Dr�F�vw-ʐq!�E�ª�9 ��N��n�<��:�{�����Y�}_u�Ԥ� �����~7X	 ��޿U��K±:@��͊��,�w�,ʽzd�����N��r��(cAi���a�p5�x"�4N2�4"+Y�^�l����Qz9�5Q(nSZ�ぐ4}�:1�ˆ@*k(G~�R�Dª!�me	)`�kCE_p2Kw"���p�0��r�H��%��?s�Cد��%f�VwO�|w�U��e�H��4}��6[;�����J�P�O�b��3϶CB���r��[;"}Z��Tq��}�5�gnr��3LC�6��U�X�϶�*7z�u����/�;��jU*Kť�[��ES����sg[m�$�?w�̿�:19�Te���h��95Y���
C�$����H[� ��=�����e���R?��h�������6���lwD�U/x+:�"��5�ᥨJ��G���5�Y�Q�~�m�c��V���ɀ�OK8�3�,�_��R^����)v��gd$��g������ �������h�H�:~���e9o����5��~��/� ��Ј׬5]��j�&ӎ8K���`7cГwOʕ�e޳�:�q!��.�r������qV�~�� C����IE��&��g՗��5	q2�)w��M#\}&<�����U?���i뢛|�."�b�H���;U�X�S��x�hy���tz)���Q%H��	������W�jzȳ�3_�-G��^�p���A]�� i��p�U�����J�n�v�J�W�Rl����a��%u3�+����g�J(���P/�T2�=�u��{�=+��W^G���Uir]�ۿ���E��
�h��L�8r�
"o����a�z�}��jv{�V#������2-دE}�������Z�!�*� �:��Fc�Ǣa~�!�i~�3Y���,�%ݑI ^n)䌻�D���!M1��GnG����8�ڻ���R�-?���$�Q�{b��c���S��,~
�t�˚ �N��ņ���E3=KI7q6���N��4�H{����I.�V9ts�t�����G���x'D򃵸�K_!�<��Un�����	�Vy%��}����`�{	_:���:d���A��g�<s�=�R8��s�y`�A��%�(�0Q��V���-߲/i�3`�Sf�B��������Ab̭���t�������Bu3=�����J�(4����?����{J��!��i�U��(#��h��
�Ԝ�"Y�t����b����f�� �Ҽ�p�{� ��do��7f�n\��� _����-\=Y[f��(>�<X���Fދ�ɂ?��d~�C$a�ȗ���5~��7��s��_v���F�Qt���m�Q�7yh�����:�Q�\��F5�RJ��nY�H�h���(B�ם�%S�Q�ǚ�,x;��W -C��嚪e-��Ma��(�YDA2����Gtk�*���&g�,'\�Gg�sBi��g�ш���Z$B�
	+�i4��C�M~�͊���d?�[Z�k�H���!@nsO�DwD��=_�3U$�K�+�M��m�]��7���I��(�	�!a@ҸN�)�kZ��1������\���3�N�!��~����F��Chnb�E��-�\8}Y煿�s	Y�_>����_&�����
iI-B%�
7]w��ү�nIe6�vM�IP�� �xc�W��z*���$Z<�=Ǚ_[4�*mg)����.�A��.g�,���z�6�x��H�%��r�l�[}s�X���h GP��|h'&t��X�Eq��SK�`��.Gu��?�j��
3J܎Uܲa)�QF2�𪲼f�\��r��;K�D���d8 y%�	5�u�`v]�Yz�ĺi�L壀0V�q}�\O�R=�
}>�5�`�M�WGXd���0���3z��/�]@1�����D�zo��ط�Z�	�Wn5����;`�w@��
k��g���iZ	
���'��@{��c	���b�]��Rԥ�?�5r�\*o��6gM�N�E6���H�8�:)8��D6�������i��[<Y�]	fM�2��@���.ڴn�;?p�!m�O�u��JËZI�q7��g��{۔2�z${Z��b�8������d��8�q �C@�c�~BC�����yz�RM*x	���@����+>L���V�I-�����tV�v@��X��B\�(��g3� Q' �#B�T��aC��ElgG �Ȧ#�!�Vo�M���h�R���{�+ӊ��^!C�	ŵr�Z��7����s��vk����!�H��=f4c�4V`B�3@�+�2yF��N�O�s��ct��)-�c��b�8j;0M,p�F'��o,ɚ����^�՚-Iw;�����:�wn��,�����C������X���.,��a\��cV�'�[�<;��6zȉ��|t�������w���wra�B������=6FSϻ�H^'G�l�����,��*��������VԻf;��� *[�	�eDM�^4�����B���/)9�	�u�:��b�f&����ŤI$�5�>���bŭH������z,��������DX��G"N�֤X&���qp�Y��#��ĸ���J���(����&�Ai]���y�m���J�<K�GD|*Q�Mh!��� ޔ��d����$�ɳwG�3�D�S]3Ip�A6x��6H�Kj�#<x��1jU�M�w�<�za+�Z��7���<h�{V�[%j��I=�*(�Z�onL7/�9dA9�z9�k�#jJ�E�|�i�8� C��C� �@ρz?��%�A��8=�L�R�T�FL�t�q8߮ϛ<�S��kSv-�X�Փ���Ò]��[0���5�� :Q!X����Nn�S	�P�N�9�=S���1
��6ۙp��ɕ�A���)[ē~_���F�G,\�C�-贡�b@�� ���iЅ;e��/�t3/M����X�p.���#S����X�s8wo�PJ�s
F@�C^�v��Ǐ�����<U�no���#áΝ��6�7<	��ĸ��K�?eْ����kM�-�S#j��;�{���:��Pe�3���h��aj��9���$���������%2��CR���/I�w}jtc�-��a@��p]@���� x�8��c��ay��k����
LZ�G;���=3��6�̗b�����dc�OG^����4�Ag�c ���R�e����(�-�<ܒ_1ȁ��AI�h�i�i�1	V�-�G���V־n�c�y��z�[��Q��Rȴ�F] 8l���4�p�8 )�^�N�@�d�?~}2���e�1i̩S�����6��t�GrK>
���E$��=��P���>ߺ�A���}�^�����ޠk�/I� �j��F�a�v�����yIqg-D�Oa
�p�H�fm�2x̐&o�UpҤEE����8�/w ��"�8?u���芭����I+
��*��ho��Ai}��#4l�6�u�)ܸ�z#Oގ\^���{/�X���f�g��,?�G{�ŭ�Ta/O�3��c�B!�����i��4z�ko�� )vW�C������S�}������k�����S�E�������*=7��uM	ܷ��]� ��ߣ�ut�*�5vF��~w���Ő�����c@a@%��l��0�m�$��&��5)9>"��_����,C������ >u��lx���=��}�%)T�KR+���E3�qk[� ��s�u�w=�Ij<U4]��A*��q(L����}���d��IЖ����h�{�b&z˾L��d7�e�x�����dT��ސ�M��KRD��B�\
��Ӽ�äH��^Xڨ痤��@�P�v �B� D�Ԥ�_3��O�b[〈�(�{*}���ß .�/�p{�AWd�P;t��M� x���`��Z����9��u �V^���Q��s}p��c�]�fIwaKa|"��ϵ�O62��ze~��ʳ$���-5�,P��@w�+`KCZu����¢����o�O�ε��(	T={{Ɲ�AS��f̧�~퓌���W8����t3��&O9�4a�����1�h\*�4�GՓn�1���z{�!:w����<��d6�x��ɏ�����z*"����l��܉�B뭖;<h�&�*pC頲߇�#�R���y8��C������3�!Y���cU�s߸fvN(D��$�1Y3�ə����I���<Q9�|�Ͳ�ƴ";/��i!����"޻EL�M퓰̰������qV��G��t��V�!i��2� {E���<�PbRy�4��1��$ �?���*P�|�_�>��R'��*wއ����2$�X�����y(�����F)w���6�F�ɧ�$������)�Y��Hc���򧙵g��V��r�I�*��^nv-IXc�ܜ����P�ؾ���XExy�����JF� ���,�N���O�W�����fNAw)GM�a�s���Bt@*��s8A�se�+H�?��?GJ����V/���2�I��s|�����BK~y�z3(�Y��w�ס��D������6�;�Lf�@��^��|�t�+�Wʴf�u*�0�oXV�UjRK�]C��Шqؿ�
����@n|�y[e��c��`�xp&v�Y�wJ5�EV���S��q�w�@P��&��ߒ�?L�=e;P>�|�Wc���X��L�Rg���pgO��lG�C������X���YIZ��N��w	�Hw�>�.��P�І%��q��|�07f�[�`1��l㋙i�4�FH�r�=��8O����_����3B]��j8�N�眶0�!O�{�~B�d=�T�y#�x���i�cGg��Kʭ.��_We��
�h2E/��uN��Ph���$U�Ҕ��w�ge��`���iٖ�+ؓ�	�|�T����U�[SY���"e�ɺSa���w�eA@��Ic^m��sv���Y���l'�@�� �E�^y+U�p2f��Ot�vl%}ԥ�b��������{��L�b#eq$,�M��m��aj��F�(Â�[�=5���yZtfׯL^��N}_㡏
WJ~m�3`�M�w%�fR�����BܗO.u(\��N3���m3��au�V�`� A�:�����X�h�gu�r�/s��L%��A!b}�ۈ���!�%e�X1]~{��7�
�Ǩ?� /X�[j�&ٌh�����p�[N~;�Q�4��Ʉ������(�#��_x�&VCO��P4�H3�Sj�,�Ύ�vN��˛��T�R�j��<VZ]�����!s���N�C�����w����$��v@�{�c,-����X�j�a�@.���@�I�J�{�"&�<?UF��=��c��7_��P4֔��H�%eC/��D�B���7o�Le> dL�t�[���[
l�'�b����K�9)�ofԺӠ#����9���P�d1��4hN��ּ&�oͻ���V��G��[�lQ �̷}k�oIxJ;�ֽ����8�Ё�H>�H3�4��g~�UB���+c��|p�
�e�f��غ�S����?VfN���2���~��z7���.�#�!!�
ZG%��|�F� ��E߀�Q8U�fM�뚙�	�3_R��S�+R��L���k��Ea=й��aͼ��>����;Uc��N�,� 6��7�K�t��B��O�S"I����|�����GS�o�L��#^��BrOl�h��B�a�����sl��ML92�X��}�҃yj��]�t� �������w�1�VS��Q���'�:e��Q����)�h�����kA��5^Fb�� ��|������8�tm�Sb�九�-�q0��w�iD��nO�(b��0!&"�6$ W�qj�<m���5s O�:{ ᳣k{s�EIXl�|_�U����}V�����&�f5�h�gӡA�U.(���ֳ��qgM'�We�]͑��P`z`���5.�1[yu�L@5oO�Ԅ�B4�g�|"?���W�=�"(��V�rk0����[f��

��_AF�SS��m<(H��ݏ!)L���Ip�^���}�C��U;=���[�!Lw����*����2&M;�����3etu�Q����>J�@0��.�6S��O�+G:�]��R�/�[�;#�B�:,\+\�`Ӕ�(�ܤƘS�����]�U���0���.�΀6�~�7�=L�l�G�y7�3I�k�</.,`]|�Z�!!0YL]����E�8��ֳ��Ё�}���ľM���;W	m��a[��3y?�lР����7�7G�����,-b�CQc����;�3�{��u�{��ɏ�:�e��hH���ύ[.�FB�Z։Ю+�또�^p���˜Ƞ�hp�[n�-��>^I�Y�]�#�K;�*+�?��m��&��^6n;G� �d1ۯ�Wk���s�Y��}"�_�s�o<=���[_�BI����#'�s�ԒsVݘ,6��S��5Lɥ%o� -t�I�E�@�Z�ؔg�|�
�C͔b�dU/Ӕ{�Y7l��0�~�PU��):?G�9�v�ˬ1��䖥ifV�^���-T��U�.ajtӿA(0�ϊ�3�u�ʊA<zӓM�������j^��]�������^�0�E�;ZȔ�S�&��&o��Nl�>r)�d�{��^f��� ?qu�5`����T��L��y5
�3��z��������c8��^��h^�kI�Sr�zfX�M)/܇�KB����'I7��6��UPr�F�G�^̋�#ؗ��'������Ŗ���$��O�]��Ebz:9xB�Au���&�!y�T��^]��< �*k7�?GƬ%E-��%zՓ��<�4��c�#NТ��y����'��z�S�1�Ƿ��5N��W�yz��eE�E|4�D�`2����x� ���,�w|�Y�f������*'m�3�ٶ���>_��ZH�L1\�-b� ��l��WA�y/��+اWG����\w������T��&�s��� \�:�6h��D�ϧ<���	����H�Z�q�I� �v�a�B�S�<[$�z4�5K��dl�:��Y�����L��8��C)�b[߶��$����*��j��cG���]��l�X/���H֯|	��iihm��җ�w['�� �Ch��mȕ����z|�{�T?v�{�R�/��D�9$ �;�ڽ���I:�<&uko���!MF{f�4A���^��I�U=�c�L&�W�ګh�}��Z�F��؝��Y��7�&՜N���;L��YE�e�r�~I�����~ڤ�^�T�lԅ�F�D�O�O��5཰1�D6�㐊HԿz*���~\W��Y��;R.��N	�Q������x�+3��S$u�p�=d����-C�q�i��R�]:*I`|��Yt�==����H;C,-I���Vͦ�y.qå���>t��r��F��{�-��U}����\��� T�p���;\e?��\��,Tp3p�J|c�h[iL΍�<�ӗ27O�=�d����F:��4u�k��������UD������a��]J�x�\�u�uȡg�J��5��py�Hj� Q�р�Z�]��3����������J�㠀R����Ƭ��
YӛӉ|C�d��^��r�Rf?�o:
{���Β�������b}��~�omq���y�QRRWhMy��&y���.H>4��j���Q��'�.6x���+�})^��@]jP�&��-��3n��,���w:�-�P���R"��?�� bLi�iW�|��v�(W��h�Z������J��p��fƶ�9�r�㷳y�5�>ƺ��r/J�)3�Be<�F���3�!��� ku���_%��zx�C��]�W��-�}���5������?ݛ��;O���Op��wo��1.�sa�+���+���W�ݍq��Y�Q���j��&�1���ag�[���a�a��	_�k�F|5�3<��3�,�#7I�B��|s��M��>�v�/M���j�>���+E�$d�U�0@�h���B����0)�T��`���"ap#�0�ɵ��2%A��H�?w�Բ�(䉐r���<�����\}8�������Ktr4Ԝ�PBjt(xn�����J�L�������AĜ�\#�_�s�3��hP���:��H7���;J��mVH)2�a2-G��˱�c-W0GqvR�8�@b�|�f���mS {�����C���pβ�?���A���*�Jզb�������=Y���G�����|H_շ i������_��擃�K��dO��CI��r6Z�3�K0!����*e�q�6v@�唊'��mmN��F?�ے��FNx�ɪ��3�t������#�vz�}a0`�f��:�#� غr��<+���4��7,�\�/���u��Z����Y��=O�UME'6�>0��%x��%b0Q�s��B�
K���5�$,�*���Z���P2}��@��I�����8R*�cm�RֺjeE$с�Q%��O��c�2�=q��q����ർ���:�}~�#-;�'=s��ng�'��I�2y}�?S���W�\D�٨�j]��X�z�c��/9���9�*�M���<��F�H�1��%�3=K�C��J����D_ɸ���,�������7yl�ݡ��V�E��OyB��|�)���AbH�l@?����RA�G��ఋ~-�!�����A����[�B�K�ҋ���½�`"��%Ȓy������w��e���8TU�>��@�BhF�юG�K��-,ة6�N{��둡��"0��|��Ʊ+��hm]
�:R�*Q����Z��6����B6��&���¸��V�6��h$�]�N=�B�XJi"1���_��.������X��hL�?��8�|j�*Y�qh���	�<!����D��o�E���P3 ���B�T�x�˲�C��HLݵ��ɻ�@W����4U����Q�(��9���y�j<1�s�Ɍ뗔(8ϤS�-8[p��*TA��B|��˚�@GyǨ^S2
S���F�q�*F���u$E���g��޻�H�4�|:d�W����M�i���8�y�d��p��ca-�����|�SP(��UwɢO���9@N<��ܥJ!��L)����u�:36� �v��Y@�`ݩP��)�!�b+�H��4M�U�<�������6zb2��B���-а4�jѲ�'���eQ��W_^�f��;x��������ɨ��"(����3��TḢ?��.�1%��Zؕ���Y�jK4_U�������:M�UӋ1Âg4���ƛG.&E�,sv����_��ōY�{�D�gP8�~ʐ��޳(�2E��M�WdS"}I�A��.�k�_�E�����\.dA��D��*@;��L�\h�������/ȗ��Cs�Y�C(�;��^�&@���/��l�i�Yv�k�-s�$m���"�==m왾t����5q�f�M�n}��kٍ�������;�������2h��İ�����g/;�{E1H1i-"�; PGg��X`��b*�G�A2�����H[����-�����CHܝ��h�g����[ӽh@�P����,OGWZD0յ/0�X'���1<*�,�Z���yiC΍-,��J$�֧���E;�o:y�H�r�r���X-����vc�i
���8ki�}6Z��DvG���f��8�ԁH�Me�`��
UW�K���yqr�Vl31��r���?S�Rx]m�d;&�c�ձP���C/j2�S����e=Ԟ;�<IY��X7ʬFd�F.?�Wu��-�3F��5�*�u�'e��|���i:��jk%jC٣���_O�����-:фɔ)3wWX>�vY+��w�t��.��4�/��}f�'����g)���4û��#�|K��kkx�����(^�����)���;�`��1+,�,F���-�wPЋ^}GM!*>n��]a�P��Qp��[7i��D"'1Yxw �!�2��E�}&2E}o�zu������}|�܎Z�OM��!��ܚ��s3I��F+G��x���O��5�p����'F�K�j�fNR��1y록�8������:���O�7 ������#6j㖐�����U��-�Ch4�*����I貝���j���!�ι��_X15�$�i���U�Ê~r��!�+|�<5�
���M'8����_Q+m5�}��i��2p.\6\�,V�5k
�N
���N.9e,Hy���Y�B!���o�:��SqW�`R�t�[5uL0�x̼���$`�������үwRw�n0�Cj--���a�(z��-!��n�qEщ�y�<�>Ş���" ¯g�x�ڄ)_����1�՚"0�
Vީv�	��u`q�p��Ɉ�f�N�"E��g��\� �k�/߭��
7�Na3J<�a������ʦ[�D�4�tgur
{@���#KXԑ�$vϭ�/{�f�j�ߓ60����b�'���H��n��2�k[)1ү�ߡY����//A�2���۩N�ٕ%P\��i�QUsb��e� �=�b,W�_E��	ֽ��u���j�Tx!�5~_�������캬���{ir�#������T��0q��Wmf&����a������־�R��"�I\H
���_� � �M��>���xO��}! ]H�M#9^K�3CI�4�D\
����9v�-3��F�Co��?ӓ-���p�iq�]?�C��QO�ǰ��&�����&�"�p��I�������ߜows�$������E���a��q�5w[�xF����[~xAU{Q�U��)�v�%8�����99K56�ݎ�$ɕ�����F��6�af	`���%[��l��o���~�^�1��U������Ӡi@rbR�:m��%j���H�	�6�����=�5�W\f�[(=��'難e��2+*_�ʕ`�B_�y�]Y7+�F�^N&�C��ؓ�\�A�&�����&4�w%�[�$���[Н����1:E��#�哳�c�_���>�S5��݇ �X<�gܞ�>_,�ji�h5�L����=����N4D�7�����0��0���¶�K�������8���� 9݋d���P� Z�$O�p*v� 	�!�'A�X�� 1=W̸�7�R9�׺N+^�-�) !�����zg��@�t�Y�[xȲrV������g�Fh�Эc��Y�o�3�K>��Rʫ��߹�K� ��rW>JL.������|}��t�$�
Br&H�"dV�g�b��p�"�҆��hxKR�BG�N�@
NS;.�}�|y<�K��D;�dHm�?1��]�X��Lhq.'%���x0�4����7��_��|�fm�4?�4Ȗ���k�6�K�~#��=ω��sIlc�z,��G�Re�./~ �;C�6�u��x�7L�~�7p↛�v��9A��`#q�đ]LO�k�p�����~aH�HYZ-/���D�y�4Pm�y�ި)�q����cA&�[��HJ�'���D�y]}�o��`<xB�k�i���^�t��~�T��7�E�A�a]l��鋌��?���~6[v���:z+Y,=D;aG���a�����G'<(Q��v����Ke���h&j�	:�X����'����0�:j���Y�ǜ�|�v���X2K��w�u�%��6���\���%�L�|@��8:Gu��4`o!���K�t<� ;�l"�l�tN��QL�t�Z+�N�A����/��EC�J�o�pk�܌ꥃ3�E7�;���7�7�1M$����P���Tq�ʁ����˜~{"��z�:�b+��� ����$���[�׈�\E�Djg6�ݙ yG���G�}ە��+Uw�^4>��D��������}^���ª�N�CI'��f���?/���%߃GV�#W{g�Qۊ���D|a����K�+ϲ�#��3ѐ�����(G�� ���$� Y�
��K�����%�����T۽v��+:~������^�+�!�}�`-Y�����.�Kp��D��jd
�-2LӋ'��HCA������Ȳ��e���&��ϸ�njb�Yo�&��K�9#6�"��WA��>5~%��M�<���ZJ:!��~3���d����>oC�R�:����IEN1����Hyݕ���Aw��U'w��<V���[�2�N�Y�r�7���K=�'q̂_S��5�Z`eվc�
�D�g9�t�~J8ś�2)��ԑ�,�#~Y�� �%�{9e��m���mT�Ͽ��Ȧ�L}�o#Ў*K5{�qG���H{R���N?�a-�w��6��<��b�7�\�]�/���h�e�����ȳ�'��^����cgO��2^�x�K)�G�υ����s�H�p��n��D-Ӯ��JAZ]�go}�KR=�r�-�9����m�l�Q����iε���4� ��i�K2��}�hK�����X���M�5Z��t��j;�['�C�լ�|��
9��!�v?+��=4@� ��d�叀-Zoˠ#'3^V��AK'RZu���b6���e�..2�s�F�d|�$�`�r3��xpH�&��q��% ��h 	������)�j��̓��+��{P
���ʮƀ�YiN�����\p���<;t��G��5��6V�ZN�����ڠ��K��l�?�P�1�'���CP��,J%���n�����B��dl=�k�����_�1ٵ;-8��(c�ǪDi�.��?�&e���s�}����;�A�GS�
̬Q�ͪ�9���C b�<fΟs��C�L+�ė�J�[K�j��=�����w��-?�^���@\Q��"�����s[�@��d��#}Xa5�[Ү��b�gsJc3�"k�@{�C3:[����x%m�ַ��C2|�>/o�����Q8��6�y.���(J�bj��T��IN���nLe��DZ�;��X�� ��@9�2/���K���Z=��:@�D%ݓ������A�.���7�����cvP^���%x�t�рeQί����m$y����~�u%�"3Im�s}��Y,:�`>$S��٥b��ܞVi��z�7����
V~���7Ú����v=�\dr���x�C���&��'Xj�v���̀�L����\n�o`��;`>2�z&��o��P��>~#��<W😕s_�ʗyfI����;[|'���=�~���ެճe�Zh��"�	n7��L-��i�0%\ˬ�������2ō[vL�V�#�xG��Ug}`<�>�7PP�Dj��4(@��,p0��R[ M��(�E��*hF�C���˄�\^���q{�#e�Nw�CȺ�z :���C�ռ��j�^?���&p�U}�G�Pֈ�W���H�U���>�쮙�7fU���»s��d=���ʰ3 �E�_����G�BZ��?��+���c����`�>�l�=�)>��gH����=� byu��~����_(��3"3!�zLv���wA�Ǜ���zY������]��>l����Z�v��O̾����Ae/f���|���3N(=1�;Y2Fe���ū���N�C�(�m��
��Ǣ�[+_d�/��I]j���0=᪕,-;\��&�ba�u�u���XŽ�!5��h��V�-���hQ�ۚ�s��Q�i����nw��b�=�y�۪KDk\\���R�O���.�8��>H*�/*���+Oc�A��E�ֺ�ݶ�fq"=�W�r!4�5}�q!���؋$Fݦ�k`l&�&���L#�.���� TNy�H(+Vt�7�߈<ş��C{�3oX����9�{n0v���;Ʌ��,�E���e`�J�k�w�\,��4O�H�_�}2H�9=�z�N�|?lP� AY"v;�෯��C���5xnQ���Ю���ЍZ�����T2և!$�/�����?AB\*�s���P�r���n��~<�މ�Kram��%���@�в���t� ���h:�k��G-�M�.GY@M�j��y���-ΊUj��Հ\=VsG|
��/���Wď���P�����N���r�2��,����L�h#ī�Wy�5�1�8_4T��Wh���'Mv�|��C]��/�0�.T���9�&��s*w�`^1����0����B"�d�T�υ(Lԉ���}S���>�	��@�i۹*��%�*�3�?�vQKy��6���֬�6�3y ���4���xz	a�Ցv�x��Qm���A�'*W�+&HI��� b�\��Q�N*!�FF&x	H��v��fRIC�SJb��CjB}�6�_�T}����r���V�����C?�c%є�%iW
�.��X}�[ ~���	���k�ypM�"��R%x�ڧ�ˎ��g�+�ga�y�g��t�.}���P~M�X��y'��_09x.-P r3�!�)�7�-�ׅ��e�Aܰ�1��iP�[s��W�7��ot�?C�Q�&���Vd5���^>s���["���oD�6�����淽�	@�I�-����$�y�in��d/�x��=���X�B/ل���׌�YS�?�uR��'����z�g%\�O�������D��t��Z��w�w�����9ϯ��U��.5�˝%�N���X�oQ����HO�{5�H����@%�;&��+���eۯB[�ˬ�]�${<X��/d���Hw��!S�;v�M(.9~�<�Ͳnw4vk�Ԕ����0�%P�Z)�E�8T��kO����	�t�ny�-��T82���,��#u[��<�+'t��3�4'�������	�.&U�۩t�E��pI�&�mh�'�bO%OiD� �  ����B�8���~�Uk�<�"�uF9�a:T�4]�iJ�C�kMw�9򆰿�3a5���e�~p`rA�i��!jy
����`#���+��#V��FX"(	[sLL����f͊3���69���^�bv�m\@n�OTN�Zx��@0֮	�}��w��7>G�
�pĦt5����o2`L���)�l�������Ǹ��W�s4��/m��:;+�O��Lj�W�`G�F�'_���?&�Y5h���1 ��]���4�Rӊj�y*NG���ˈ��)�2�л�/�#:y(+'Ͻ1�0��\�^7?�G���[�<W��5�w�#�CH!�tw�Q�N:�����f�z�7b�S��i'�+�F��[�<�K"/��}���k{l4q{�;_&�����?��,I�A��gŖ�����վ�;DO���UEܗ��e���3��f2����a.^4�jh��p�&v���).����p��S$�*�Z�"/@jϾW�G�܇N�x|��@�1�J�xs�"�qgl2���|�z�
�F��è^�_<SuXU��$U��a����R�ᚦ�-`��Q��{d�k��h�z� ϝ�#C#��\�<Yְ�'H��;�^�yd�I��vO�Y�ygL�������g�U;��zOey�#�Q:nώ�	�u�Z*Y@�w�P���Q_�8�����&��8g�d�hlЉ�>�UFÊݕb-�!HX�4���.�>B��յ �xQ&�7�M�h�T3���^��!��+�|�!�ak�������ǲ1��&�f�-�4i��<� �bխ�T�bt�$���;����
�p�}j�4|�f����q�@C����0�����J��ˁٚ���s/�+ɑ����pp��������GI��?7 ���E�B��M*�4���]�x)M
!Сdի�d��yt&�� <��<__�^7��ph�Ԕ����7�1
đ,����^T�j�}�?�W_���WxN*���t�d����&X���\�c��y`0x��`2�K�2ds�\}��lۧ����$Qmu��Ƒi�$�c^��7�֒�+��u*/�������}`�p4/y!�CM�BD���o7��՛�,�'$���'��r�>����]��3S?^��T�7��l���ۛ��#� #���M�Z���t�k^m����jY��@rR*�A����07F�kM-�?,�qB�Y��L�'a��p���k��&.�[G���n6M�R����h�˦���떂-��]�����'D���"Or������=j�e(��_9�6J����E�v{K����#��%9���N�Z�E�5]�s�����8g��	&=��\Z!H"�'����.a����Lk��
��WD<���Dv�L�R�TjWB�����~��H�ZN!���UB̞��{	�k�ZkH���7P@8��hfI
��̅.��ɀ� ��;���p����6q��Y3�D*i�(�k�t��Q�O�̉��q�%F͍
G>��.\(~>��st$ﴖaD�c�	k�I�`���w�y]\�El(hB�@�gϮ�MT�J`�L�$�/�o��m+5�Xr����\�o�!��g;�l�[k��3�����Ї��{e�\BU��9��F$+�-&�wuxyi{y�GbK��x'4��ye�d;��$���1ZR�)>���ޤ�>F�1!���&':���AF��1�%����H���F�m~�<�g81D�1�.V/��/f�޶G�%מInI<�4�pA�H��n���a�`cV_���՚�M̟�a�$P����#���B���3���Lh���`R�Y�2螃�wL@�ˉc�rȼNq��L���:�%�G2TP�b��O�> !@`�+c#���7n�U�MP޿���놥9�`#��{��{0�x�^kf�4�b��o��Bb,dC�^?�!�����m�@�T���ȯ(�
�O��f��b��3�̢6ͮ�`��O��j��y��8��/['\v(� 2��OG2x�G�� r~Ʀ\'��'Z~�V<.?���JȘ�� �-�3YR�z���o�V��׳t(�ҳ��kV夗D���f4yz�1�_�)���%`�O^gd��3����o�8L��]�I���wp����g�3��;O*���^�eY4#燒곍t��*�q蒰j�B�6�*����x�6Q�U���¶7ZXIr�m�6�ȅ��SN����	%�s֤���DUׯR�f�a_u��LZ�f�#��L�,@��>n�΢���N�iO��ͽ�!�8K�^��7�,�$e�B�l��a�S-���tZ��X'�	t�.N��Y�1�`bUx�I��O�P������.q�(�V�:��_��r�N�[@�Ij�4e�{iN���m]%S��M�Eyjs�����Er��״����.߷��ևuR�v��6;�a�����Xnc�
�|����`o�1�p�P}L�W۱�H ��iJ�=�&��]B����e�QV�/��//��.��o�� �|����ҥ>�:�B	T.j�[X�>%[=�ـ�cP��>�/�k�i�W����9|lw�Ԫ�JM����叾�|��6t	[�? �+��I�y�׭��'f4k�h��
&0�N��	�>��7̺2�-~k��:}GJ=�Kd�ߤ�dh\r���pח"qzSQ�YDU�cG�ƱD��T �E�IG�r�7��Cn_2(�z2��Ր`�rT�C�j��$�^��W���i'��(��*5�d����c���E��<�X���RH{���kh	Ka���V $�l�ؔ�gГ�2�ÈIUZe���	��e�_ϓ��5�U������������9%#�Κ>=��gI����� ���B�`�qԟ�*b���r��Y�+��#��["�/J�UW#SF�m���e���f{h�,�<O�V%x����L�
W�JBD^�A�xGq��B�j�I�E^��p׏_[G�F������/YGB�q˚0	V07l?�8ۂ��zÀ�S��vQB��A�0ZM��k��O\F?Q���=��1�^��(�ܚ|b���1U��M�<�`%��)���	"Z�m��;�vKt�Tp-N/s�/���!�\(w����U���&0#�o��=�C�델p6�4|1R^ԝ~��z�Q����×�yIEY�Ѩ������8�K(�Q ��/�N��ɞ�D�w�p���L����;@�6���o�a�o˺8ŧ��\W��)�`Q �&h�����M����B4���p�o��&=��06�WL5ʎ6����f[�A��<馦b�'���@�Sz��\薁����X�a�C�+P�l�:�M�!����ޞ����� (�����/�]��;~;|�Z���l��y�T�]	mY���m��7��-	Ƅ�;�b����0�|��|o��ȭ����C��f9����m��cz�mE���;e�Z&A= ���d�V#��(-9$��S�w��<Ew^}OE��ɹ/��������M�����ф����X"	|������4[�QO�
�����۳l���JP�G����B���b�d��<z<8�MI�Ô�u~e�%�<|�
6�����k��v8{�DB��P6�t�
9VB���.D���i�����GL����[NQu������&�����^Cd�x|!�T��|�7A��Y�7'���#W�˘�k�x����Mf��3�͇����5|��V`��#��⒬��)��g��6�!weO#
.iʊ���߽$��=��Az�m��4�;�~А��[0�-�u��<'�k�����y�����\��@HG��ģ�����rJS^���׵�@�M�P�t�s?�l�x9ݒ�*�#�Z��?+|lu� �%~��ID|�^!���S�=�Q�>���N��:�\�T2}
�LIM��.�����|���jQ�U�Q�m���ָ�!7zbk�2��n���`�sز��%Kj�ڸ��xiEQ��ܣ�ֹS���!�����ݾT��a������wxn�Y�l�ǝ<Y�H�Ue��F�29��b��_�����Uk�5�c�ryJ�,�8=)�e���'	΀�y�'�3w��I[�]�B��u���M_�yC�;�tI�}�0�	y�JҾD'����	�G��ٮG�%;æ&�?=S�|.N�4�X:dt{����h�ׁ.Ԯ�mF7�������@<�\�B������� J�<b�UG���`壠w�#h�p:�m�.̡�W��~�IJK�Oe8�z�Ak�mS���S��rJ�� �G��m}/��� ��AG�;y?�f0�ml����%gS()��_6��a���AEuGT����9�W�YqV��O`e�K�Z׺��t��˻�����+���:�`�U����Q��e��}��Y���Ъ[E�����&��˂�h+�d|��AU���v��6��7��`�L������&��|J3^M�挞��Q"ؚ�M-AJK���߈�vJL�����V� ������o,�]��6��Eǎ3�h&����� ���t��;�^��c�V�8��ŧ;�C4Ğ~E7�g|���.������C�|�U�Ef	�h_t��вJ*m ��^$l�I8rY��n��R�@�W���0���<��������cXO�_Lv��f��I�����x�/Jck��Gby����]'ɣo��!��2{n��WY!
��.���5�/��>��w�Q<1�6��Eu�뛑F��c�������{|G��}���t���X��]	ѱ2GS��S��F��Y
W������*��#�����(-Ͻ)GĽ��RI`�N�g��U#�~1�2�r��Kk낢�H�3����rjt �B��S�J�eIH��hyx�~�ĔH;��w�kd ��H
	�N麵����~t0XՊ��@�A<�2N��.O���׼�:�Y�mP7�D�(�Z�z��v �j����t��V�-��hZ�e� �u���xRl�S�֢�F�g��]~/�� ���h��Oa*�q�u/�0ݍl�"1ӹF���a��o�n�ޗ���ܦ2Qׁx`.с�J�S%��NQ��rg$ռ�,�v3Q���+��v���0�j߳{��q�0�ˇ�G���.����Z���F�����<G�>^�g9A�MD�L1�7�Wۮ�n۹
�a���/D�^ޛ�l�#����bz�1�D5��3q(*���W�t�N��ThYd{3H�p�D�$��&olF�m�<��n�-�£<Wa1��u�T�[��&	�Um���QSD?�G �Y㵣J�v	:qb�
��6҅G�>s��eڒ8�vX��o
!D�,��_cz:���9�F`{��/I�߼�C9ɭ��?%���qa����5!�{S��P/X� ����w�K��c�S�����V��aD����������d�2>p{�Kռd��a�(|.ί�1�c+���9 ��L.�]�� �,�[�N�c,nr.��ǂi1+Ύ������T'GE�*7���L���1�4a�w7�׭Pg��wR�F����8m�̅� zIh��=��w�Yh���m�n$�P�W�i*��<�4�>ߏm�D�A-�t%����0	o��H��T��r�u�>7R�3��m[NZՅ]�R�Y6�'L�]�:������U��L���@� 1!���p�@|?1����������CS�9 ��d�J��*��%����-P��&�S=��\��;D���3uc�$1��d14I������.bzz|�cu��$��O�s��� o�!;!�ٟ[O��q��Ω�-C.��Jd�G��Ni����
���G:���#��H/���Pw���#v��9$�Cw���YJogtg�=㕬��$^�E%4e�-a�GF���:�MY�/�%҃"Kff;:H9�z��`8۝�� �y�_� �d&���c�	(AH���y�\�^+�he\���`ܬ��V��a�kѴ�@�p��Y�e�_E6�0y�ӕ�2��"�8�ř��l0&�!2���*��ݹwe�+�<���h�e�9���U���ԓj�p�WO�,:���Qxz�}��}	"c#�' ����";�kv2���L߬����sQo�@�e�JK�~���m������Dr'+�\[��S��֫���o�'�Hy�����%�r�!��E�K�#���T9B�0J7ïҢ�q����"���II�2��|'�D?�)xC01�*��t,��0ku�au� tlM]�f�L߯�v��-��)�IS+t�@���uv�����t:� 4b�^4{��R�ɮ$�f�9'�:Ţ=�=�Э�0%a{M��i����9�k=m�N�e�����%q���f�fl��*Xb���*
�UX9 �����e)����"�[���d��2�p� xf�_�"�ɒ�9��u�TCx����.F�z���ϳ�&�~����`�������Z�@L�x�#69���Nyu�0P�,��>$[�ZFw�O���p48�b��}�^��r�:cMНL�'�h�0nr�-�*pj���A��[^�F\|��йf`ZIE��2�,�N>IR�V����2�1����d1i�qC��g��L��t	�(�5�V��y��E3���#��l6N��GguNKx�n�f�@�� �����#��,P���}`�Ͻ����6�h����Pٲ��J�C6j�މ˛�C�E���R��&È~C���� �	��@��B��A��G��y��Ґ��t�r�)I�	����5���	�8Z��Gy&�05̅�vOF��r��	��AHя�a�_Q�Mˉ�����L�/���؊rP��"zr�׃�;����p�ԙ�D%����K���)@n�1����.5��siy�X������d�(��P��L��ɿM���[�!#�T-��Kq*	�{\R̵3�~��u���Og�v��X��I"�+v`VY��TT#�G#�g��`��R��k\�R�c땚��O]��d]�^c�w��x���h4�]��|�"�Qu�i/p'ɮ]���޻�]`y��w�����������i����Π� �]U���or��Ư��h��� �}���f���}U����
�p���{��;���?�$�kh"˓�h�CO�r
Jl�R���R��_�3!9Ω�e2o�����/��M��}��"n�rѼmT����;T�̄ń�'��炎K7��y��{/ƇW,G�+�pD��"�a�������
�|e���������.�9�,u�. ���ad���X�@����h*�Ч�g��j�@o�D-�YY�}���;
����S��0t�v3�m����Mg�j���s���I��k���7�yL���w�6���ܤ|Ӷg��JK���U>1��f �~L6�����`��-I�~�k�@G�0>W�&�h�JZ�})X�HZ�@?��6'+���|�FO_)z��eƀ�%Z�wxO��`��-�F�2;��d�FӲjtAP%x�Z9�v�Z??�?MJ��s�޹�M3����
���۽C$�'E5�"�h��VFmŭ�c�%V������p�{Θ�8,%]h�r�D�}�1	z$=M��N�ؚ+�w�imFVe�ǡX�xa��T��#I��o�V��0�PE}q<=�}3�%��=������3Xa�J 7w^LWlEs����3|�Y��F�������;ÿ��CaNmuQ3�V?qnP�+ V`x�OX���Ī��"{;�2��H�����jgZ��Ů9����ʁX{�JhIjo���Rc���w���YWBEmvrx�R��ը�a̱�~�OB��F0&aFm�lH��j����!S�|5��n�>�(Χ%N�k��'��1"}�t@��7g�K� ז�hƬ�L�o�3�<и~I}�,O���p���s����1�e�Aջ
�{}�
Ĥ��R���(�s�C�R�p���md�PMeEBs�h��ӎ.йW�cFl�N��_�W>QG��פ��^n�<żj[e�&9��*�Z.h���.
u<'��^�,���������V��|/����ቝ��AA����I�8�;�4܂�$)AG��7qD����K�5J�*�J1 Jl	Ӭ�&�M;o�Y��t�g�BQ�t����ڬ-{I�q,�ԁ�
F��a�`�ս�ՄCs�����Z�$[���PZ�?��WG��>a7��m�[i��W�t����Te�d�|:_�Z����J������@�����8�iL�BJ�ԟ0��_z�w(T�##m�<[�M[���͒v/�g��z�*~�"��sr�Y��I<k����E2��C�n8>����L��=>x'N��sH���/��1�� %b93l�u�lA\,�s����;W���$�]��q�`�7W�aZ�F����16ⰲ}2⻩�������ͥ6��od���ˉ9�i�x����l�����u�H�E�Z`��<��m�smű�'|����jD�"L(����oCC����~�󺖴+�݆�`�Đ1\j�uK��\��7��,�1�>�e\�D���W�d���X��哵�L�5�*k�y,����s�ŔOnV@<����F:Bа�G�Ph��Eg.����b�?2�����y��E�#.⾧L1����X�]8�l�qX��������[�?�}���A6�z-/r�,�jO�Mjv�[ziu7���v��E����z\�;Ͱ��0�q�F�u�ЍPv1�M�sQ���zm��>_z)��������m�/� �z��qa2��)����6>�7��Ȳ�VMnӠ<{\��D׊��k-nk�R!��Bb �@�����3���t�qNϓ1!�I�>����u?/��P+�j������w��gD�g�T��74�0���s�L�.���X9'b/�B>��QZ]n

�K�!��S\��C�'�"����ҡ<+�]����ҪW��~{����%}}����t�ԁ��fcF_�4 5�����!��n5�Oa�C�Cbލ5\��nv��P�r�xiXǯ���W�K�tp��m��Kl�_�0���e�C@��𚬄��Wn�!��V��W�^*��7K(�۽)5^�`�t$`PoN�����ơ�O=T�C�~b���݀�):�����
���l��ajB���z� ��~���X�Xj�3kr����=�2�b8��Ec�$�4��ya�}k\gN�B������O/T���y;J�i^VV�ݱmk���֕�4���ؕ,����yC���$�D�^m$|�<��>�f�b.Nz	O=3�,�Y\��֖1������h��Ç�7�6���z;�bD)�#����R�WR��5vM_[��۝�kj�hiu*����)�97q5N�H�M��/��i��f���X������Xh:���d����;�YdfP�S2�#�y��`�*J/>D�t���ϝ�w�ʛ����Z�^�8әV�lgk��5�ߑN�k(���Fo�V�������fH�t���o�z��i�M��
�p����� �bP�,���1o#����I��#�R��?���t����Ω%������:TQ�"l�2�,a��a-�������֧����*H��2�bPk�#V����@�9���0�`(�o.?o)#?e.�B�16�=�(�
�5��!�ڳU�������WL�f�� <S.��Xh+"��� �]k�ۄ�r�5=_q ���*v�%k�"��j�%\�����::�C�F����.���"�X�:�
��"?�$�B4��<�!ut>U��;�ܐ�$�m�Tq��;?�Ti�'g;�l3�1#5�鋸�W�[^��J�����yPW'����bJ;��Quxd��W9�:g0&��R	QM��򆺅����b�$O�/��p*�`H�c�����D�Z�{�-,u3�?�rs��S��#�i;�^�[%�Ok��%�"�KBzGD���4F'9��L�ТXN�iF}�!�u���h�����-�*�AO�
���6ܠ���w�QI��X��a�7bq9r�_o+瑡��5�#��/J���fs����O	z雪��f0TE' �����-�Vuv+u��E_E��ܒ�w��%�d����/C0��#*����1[� 	Г6�{���8iY�6�T0��M��ǲW �Ö㙒��7G���t��޽��R��	���������K����?�y����:Ә 4i݁g��H�e:(G�a�W܋�FNES� �5��7�b�/ B��&�W���$e� �Nz��S�V�zkR$���5N+�A�8�k`p�~�4"�ښ_OW؀!���^��1���j�?�d��cW����ϓL�/������#�fb�g��d��m=�(�U��I��q���ba�6�1�i��AN7�o7�c�?N��4HW�jɻy��������ʅs�C �ג���u�_sho��?}��Z��W���O�ۼ	����L��H�I��f��z�J��i�F��gMKӏHy�;��w�Q�+?z����?�-�%�!��HYۊ$Ȉ�i��(�+�7�� ��K��֛��t*֒7�/p��xi�(�������8���D�]�'�(��������w ݲ݁���dIt��6�}���;C�r.�����8�Y��B�f�������ŀ2�&�Y�Ym�\��\f�/�3��7:��%fG�BED�@7��T�p�&j_�6����\e��-m��KvIz���M>}�f������M��k����p�����!,t��J����qB$P�9{���Wl]�v��
瓚ɒe����bh�O	�6��0l�~�R9��8A�a1�1�[�CR=˷\Y�jY���1��o��v����$��Od�<��1bb6�P�蓵�dk኏�ع]�c��-�hpC�v��\�Bk�`S���o���3�.X��H��f�C�%\�\@!��i4Qy�ֆC_�#k)9�����ph�l)@x2��*9��>a` �м�"�Moy*cH�Yl<�N躞��JMpo�7�U�% �4���3Xha:Ͽ���U���)`J�*Z�{��.j39�)��;)v|�i�Ѩ�21B�ۍJGW�R�_E�=u�y!�����e3�17>aq?��_S��43���@�b\�Q �pn	.�f��q�����Y�@��Ͽ�6Yb	Kg5�4����{wf^��R/_(N��c'~�N��U~.��Eq��s��@Z�\�O���a��A��&/R��W�JLX��В����[:T��Ȓ��(s���Sr�����K!y!�(4EQ�1�W`�ʕe�Nef�P���6���5Ͼ��;ΰ��T�$�;ܟ����05��{%O�/b���N����u���Y4�ɯ;�1�,��%r��=؎N�����G�\��:��C$����wD,�p�w���Ӣ/�`�v��2���t�t@�JI�+3���W�Q�L�mK���.��[1����NI�����3|�	u�$u��iQ�"�)�c^u5��������xb#��Ē��YSq��#�p��Í���8�S�n�0i��|���h�u�E?S	���%,�~���cy�'�_\�
�2X)!�n��������pWȽ���|l,KO2� ꓼ#�H��S��ؾŸ�hh�Y,�@�{-�Ѿ���sND�hkuwL�H�6�S.L��{�df�T4���bx���O��j��M�e���̆Ԝ�s�b��T2�,׌1�|y�=���u�-nD��C�t�\Q������0��7���Gq^Ev��_�J�I��Pj�Mq�t���X��~�)(�Y���sq��
�,�*���T �iJw6u%��{��)�m �ʨ�}9�Ixy*w;2��t���Կq��g�6>nP�m�k�ūg��j��;��Ŝ�ǵ˃QT=��γ���q��wO�#ef���+֨E{�B�PH����a�6�*��ԡ�0��J��iK�.'4n�z�D��Y�w;�R	 Qb}�D.���=���)����Y���%�ۇb�C-��ɼ�i����D�掊��]
��\�r����槺r�#��)�QC-�܀B>��-u�� L��o���!-���,'%��B
���L����.p���ϱ���D��kR�c�Hq\#3��`k�ӻ�H#X�8G���jH�M�+�͇���@շ�U�Qj���K��Ƕ����Cu�Ӌ24q���?NxM�HbS�	n��B������8�S�P��A�%�������<�j_��I���ͮֆx��%�������|B`��ɜM�s��9��b�~�S���~��Rw����l�͊�7���ν�b���8~�T��#�x���N��f���奾m��ȕ�0���no#�T�͘,q�7%�9{��+S�8J)+��������w�+^���0��Co�C�ן�J��y�Y�� O��ge'��No�7��S0�"M�f���G���5��2� <�( �p��U	���+19��A�,��Ji^�``�뀼dJ�qy��C�n�?���I�5^����]0����g�1쭻�{o����!�2p�{�--�Ї�Ίz��qy24#�d7.�ki�d��;��w�C��}���mB�> HY��{�)�q�~�+�ܔ�^����NǉB���s��+����x4f��s;�5��j�Y:�d{I���/SǰbV�#Β�}�+����d�@�Ö��t���p ��&�r縎1"�x3s9�!��e�2! 6yq⾮w5N�rC��x����������]��;Qs�o��h������\�ܝh+��P�vL�;!%(S��sڍ�JOT�7�ȹ��o�w45��I�lA��Ϣ1ZhXd���7�1M8���sQw��	ukH�e����V�lb0��τ&���$	��x�^�#g��	��[�K�����p~��5}��"���(,l�f-Ā#!��8~��t7)�UzW[�TtY�P�ぐc���2=zC�lH������
��Un��9+g�H����W��W�;T%i@͐]��6jqUt���L�q#z���vb�������t����9�#p�k:�YBv���c�T@v:8�t*�Yo�Y��y,�aF�y]4kV8%m������*��T*��X��o=�m���OZq�?<�,6g܇��K%�	�C	SgAS����$�Ą�J+G�藘ߦ�^q�l�ؖ��Vm�r���X��)��
1CfA���V	�u5Z4�q��<f�]�uǱ�[ƯR�VJ
��:�L^�l1cFӳs�~�Ϻg�:�s+�% ����4����DU���j_�3��X�"��T� ��ә+|���)=���w�\��4��
EfD�����:�j"��~:znw����>��?�q=hET1}>,�'p�-n�J��,ࢬ� �����ߩ�����=P�����^��"�I�d0Ɏ�C����@�Jk�˴+��Pʬ~�e��6:m8��̤�;�4���9ZT�=��mUȨ�+Y���$�D|�	.�o���N�e��2��n��J(~�Nj��W J�t��|	QA��9-Dĕ��Ur��-vZ��p�L�iW���t�&+W���#rv0ӟ2z��d�^<˸��<vXj�[��g��g7�uϏ�&��2A���4;7P�|z�k4�v�1��t�#Q�ViǾ���{\�.�G������j��%�k��*bm�&N=4���՝�gdh��� ��0�lZ��
6��[m����j��i#�@��P��PW�	�C��L������Ni_���fg�G�weL�݁��=�O7��.�b�u�3�t�"YUy�}[>Y{�  �O3 ��3�Z�'Rr�W��Q.p0��wg>7D�+?�fz(��X��V ��\[��������y`|�� ��ʊ^0���M��wU��x�n�����w{��GSg!)���=�RDy�Z O0�e�H�u	f��96]���H�����������2A�!�p��J�	�~�N�˩4s�c�_�z?�w���T�8͈^+��Cqy@�Z��ļ`�틱U�����}�S�0hu*�ۦ�R��yn�$5�Ql�p!~��f�Շ�h#cRfw4bCR.�F�p�Ro���`��2��ɇ�#
`��!-�v<���o�R��4y�T���ᰰhQ��vޔ��?�J2�m{����j,��mF���"�b�Wu���d;����
	�5�R�x�yՂ�-��~tj1���X?|,�[��5fK)|���P�M3~���	��OM=�Z��^��ğWy���r!U����:�?
�0���)$iռ�!1������P7#�v���� nEs��p�U~��V���o�'�@���;I;n�Gn��X���s�2�$}�pYP�t���z��!9���'��c�掎H9+���W��1a
�Y-���T�轴>�G��z��K(�)
��7m ���J���^v���C��	"q���"GG��Sl"������Fun�"b2�ن�&��m��3�53��@�|�{��
V��yB%��&�ۄj�������&��H���P��z����[:�B���G��a4�&I��#n�r?������.�����uAN.�m`�e��^wk�
~Si��A]�)=������5I5�o!^E>)���H���P��]x0]+5�ܙ�$����HW�bd����>�rFP\�/ ��e.
M2'�Gݜ�̜|1�J��XPV�ܪ�*�C�� )�XU��G���@��5�<6��/��e��@~���c����+�*�Nm��޴�����D���+��& 	��Ϻ��a�-�Y*۫�����6���A�����U�"0E@�}��l���x�`��BV��S݁yA���f��a���]����H$��ﺍɯ��_\*�����L���n)M�3�U�3��fpY2��5&WsF�
AcD0���x�cxӜz��Чtqy-a)���Ō�W4׵Q�4��	�:ؙ��;���c}���$!�����˵������q��e:����R�=����Ex��E�I
b1�2CV僖%Y���פ��FwY�>y�)����R�,��� ���' F��V�տ�f"���G���s�,�u�L�D��y��2\i�4���>��7}Lk��WZ�/�J�U�8�I1�����$�g��|���(C�ר����
u	��;p)�����"N̊�O� �O������@!�d�)K�g��6ʻX�4��^�a�!O��;9��e�JZLJ�5�A� ��9�a��	��.�� �D�i4���c3vn�᷇�#
T���( o%3�{ȳ�a�WH5}��Js�@���lg�$�"�;����:6r�¿�{��=	y��7�!yfbĤ;A�7O{6{g۴�	��g�0��Ϝt�y�nF�D��!ٝ����x��Vj(֙����[0ᦂ8�1줲u��c	����\7���|w;8��T�A8�3�@\�^k i���\r�"s���ޮ:q�n�Bcs�c >��.,� !���)c&��j��7��}��S�Ȟ(��k��=v��r�۩"m��2)�?��X{~
�!�d�rUˈч��*$A�y�m������Zv" <�M�����
�-;0fm;����|��ts�� ��\b~&*L*	��W��t�+<���g��Mâ���:�� ��;��3O��gU����^{󮎠�cYv�9*�(��!���7s��I���>e��RS��p��	��^��*h�cy���|J-fKD�j�L��>p\�)+D��o�E�ǃ�k�؟hhC��"��̡���)�r���0�����}0�h����,��B�P�l��N�'v�4?�U�.w�L5C��$�a�����ɚ� :K�+�������Rc���mf��
��0�cO��E�9 Ԝ�|�������sW ��F�l�Kcx���	��Ьw
X+��D��Vx�'�y�K�REp~)���-m
�<�P�����\¼�ey~(�+Kzˈ�BiW�� _Z(��&��WQQ�+�G.qݤ+a��10)=B�����D�(��.����9X�Q�O<�z�����%Ӳ��Sxs�*����┱*�_6��xs[S�^���7���s�7��Pk:�)�|�#o=��T����~/N�X�c���\�������a�Z�j=ۡQ����E���S�����.��.t���!KF?V+��!�������Mi�_8Z�,V�ZV���&%|�j��J��?6r
p���j[�!��ݒ#h/�,K)AM��A6������|��]<�&����uB�Sz��X-2雲��! ffRY�\ӄ��J��jh�ڃAg��+�;*������!WӀ�t���v��6kD��=��^�-+�����<[�X�X��L��[���b���=�b-Է����*~gM�"��R���w��V������'��p��.�e��l!�^Ql�����m$���F�x�F���.L���[�b��$�,w����be�ݼ�L��%�U�<�Z�9�}�
���gF?G�)8�'����/�\��|U�$�m�fM.���˗oz�,,�Պi}�_�##�����I_j(7?�эі��k�� �Hp �i�]��
�!��U�*�5�x	u��M��6¬O*�C���E�	�$>ފ�"cG��,4N¤��T����2B�N�����^�������8&��G'�]����r�GS^\ڀ�w-�T\t�?�A:':~9#���$�Ys铷"�lp���z��h>5�����X��f$�q7ګ�����"69��0[

���B�+g�����k�>�Gpɶ�7|�Op4{ٜo���4dX!���[d�݃�d���QXR+
M�JP-�EL��V.�r�3�����8���IٰuȲg���o�O�Ś7��f1���2�O�d#���xS�Z��<k�����B�<_ϫRdIke������Z2سm`�wяv_�N�8P@��Λ#P�χ�@/x����xv�>:�cv���5������S0�'��[��L�U�~�f�djbs��vH�7>'��m�A53I�w*t�])��!��/��Y�iP�{skQm];�b?;�!4y����u5.�Z��eu�>5 �$٨T����ua���mm�fv|��i�����0_��u��"E�%�5�>죥_�/Nx���-��#��FrwN�C��cl��`���V��sv\����(����b���n���yu�Yu��>��X�������O��0|��Z��#1�o�Md�EB�8F 2�����3�K�m��Dd>�Ee$��BY��7<�n!�Q��ίI��$a��i��-�AXW���P�J5�ܕ�A���L�Z��6�T{�}��E8W�:���{'��LG�B�����j��A'�hgP6h�k���]�M���Uz���3���KT}R�+IO�q�=�e^��J]6%E�����a�Yӳ�d���e�Ngf��r�<��V��=`!+=?L�?�k2��!/���RɅ�-����8���\M��&H��O�i,7�Z���m�k�$��< ���!n��b a�4��)�mT�3��Y�"6I܇B�5,�V�T{��V%�:	�j���&�>6�3D��2�.�c�7 �֮g)�A$(��|����ؕ+A�o�$*��K��"fi�T��оV�3��ul�\O�̍�� Ȉn��Cp���[s�BOxpQ�Xs~�����ej�+���l[`Ϻ�C�Ɲ>��(>��Ɗ�m�\0�,��!�B��]�Ćӻ~�.{��^�o�o��߽�\;�BHu����{g:�^�Ll!O_�������jS�9��V�([mI�B�A��;zȼ(}�:-?���3}n��b��awwl6�0�>�q�gM-+A�����/�<���|TJ-�Mʐ��ߚL4� �ۯqov!ep1KZ�����l�X������a
�t#�5�ܓ��}卽�Rԫw��7�Y��cW[�_�i��M9M��B�s	����'��}�U;j-A%���6���/4����G���.�X7������U����&.�����1l�����!��1OH�Sr�g�-��X�����#�؟/�y�ƑbB�������`pic�}��ĆM������:zn"��k��q 2si��!|T~_�3p�_1,�\�ϳ���)�#���b�EC�DJ�4ӷ{z)�Q�a�0{�����yiп���
~����`υ����"e5Q�N�6;���N����� !���~�]�!4薡?��)��z����ΡM�*��}�?�&=*�[��{���E�@��#	�;2�4!�Fū�p-�&� ��$��U[׹(�e�,Ы��(n�>8�F��x�̀�.@4:_�8���&�`�1H �,b��9'�\�"��Z�^���ږd�[��<��J8Sڤ��P@��de���FA�u�ȳ�-6�O��+SO���\1�P���	� G9d���
�r�UA���`J	�˗k�m�N~�,�'-�pY�2��Ir�i�k�K6#vô^�����,�ynH�Z�zp�coDK4e9q�6�6���啍�	�!��7Z
��{���!Z(s�x#��+Q�n�����0v����P�ܳ�=hLn����~{�Q����W��(�!���%�c�WlÛ���|�����J���et�|Q�׶�@}������^5���i�夎�Ss5���|���<lz)�-ޱ4��f3m�i,:�׊/�g��,�+��`Ƣ�m�vr��%@-�e�oHq��z�q?�ER����6�5R�N-���T�6�WTn�K��k�[��D�D�D�%c��_���&`� ���P��|��o���������Iґ�N�c@�3Y�V�j�Ik3�h�t7�v���������������9��͙�A��g����L)��g>���[�&�����j$F�$@<�����U���T��d�@�N$�{�C=O�LG���o�/x߉����H/�8��F/1̻.����L,j=W�i��ĺH�e4MUo ���jh��2jD����C�m�J�r.��A��eF��������W@ˈ�>�i:�z줛oCsV��,n��1l��XH$�L%d ĝlخW'�f���'�'y��k��/�ֵ�P:����I")^A(ڸ�ƊuЅB�6Cez��s��?�l�h��4g�Զ�4�u�Ÿm�%��=�"-"1G���{�Y.TW��/�Ԭy���JD���yV1Z��n�D�g�����0y�'���

�� Z)�'ӣE�N��)gX�s�u�1�ꡘ\����Y���6�+�Z��LG;�����S{��0~�A`il8��2���W����'��F����H��j�
�<�_?����uE���p�1�gM-����O c��F3yQs����	�P>7��]V�˱���y�h`V����,an�bݑ3�z;g��F�sGv�_��T1�6�n-� �CJ~X)���z���3[���RG3���y �s�4Mş�ŋ~9�ٖ;�'ק��I��� �=��KVep�����"��m�����B ���(�j⬍�@��$�qEY_�e��=�}-�)�S��}R��`�E��9�����B���}�r������:ȇ3G��
e"V�|���O�3���-t<�
w4���&��v׏l��{V���1=��3��{`0���U*��~_��қw#������$�\/��0t�	��ʽ�|m5?T��f�/��=~8�W<�N�u���S���24EfX�������s�� �n�]��d�C��ư�YZ����r��*4��GL�����*әz�<�ۉ��P6(��8�'�2��M�eJ�f������1���1�� >�MWC�w���P�H�,���e��M�|�9C�_�rd�M�Ipۻ%yhE�M��'����q�a�z�_yc��V^dܢ�&�,��+K�m���u�
|*�K]����7t\7	w��g�'j�m�ÔR4���1Z�X
��ӕ�Cŋ傖>c�3O]�U<�����(�ڭ���HP֤����
�Ga�S$�˶�ū].L�`��6�j��;Dq.��E����elD��Ae˞4U�����`k���Ʈ��ߕ��mƞ~�y�!�B5sL�.EF:в�o5�R���qnml7��z���#r>Q&Z܈_�L�_���»�S�%�H��;_���.q�ys'�V�c�ݾ����ƨeyNw��zB2C>�P��
��񱣥T�3���?u�ט�-�����~0�@yi<��r�fV(��m}h��~�R�?ꝿi���[MH�֦�4�#ߕy��i$�v.rj�A�a���,��0?�ԁ��k"Z�5�-N����S���jh�{۔3��l������2n��ۑi��Д��.�&?�4�a� ��������i���f]����Z��c�*c��~ɣ=�P�
�C���TG�v�E	�Gvl�Y��^��_G(���ʿ੆N����"�� *����K�����huܰC�1 �Ȋ�M���hUV=�(�&�����zt��#d5����N��'"�Ni�4ϦT_��`��ԉK�7C{�>�>��1e�o������?"
ө}�'}\�(H��2�wc�OJ�Jt��ޭ.	N��k�yb��t&PBZ�KK
����$�7��zJ�
��yA�����:�ح�`o�G���2��PJ��&����h=àl
.�	�W��y�=�l�P�^ �~	YI�G���KD*A��#�7��,��Ǉ
8%s9�^�r]�u�O�6J잀�vݲ`[8�?�(7'��hb�r:�Ź4��u0i����_��j�yR�����/�{
%��-vYG[o���Y��."!-f������?�a6�} W�SN7r���3AQ�Z-�1VeF�s^�VHl"��Zc
�QѴo��?��a9Q2�i};D=?��m@k�|�~Z0�d4�����V�b�
�;��+.�%��r�j��r	��'�����>c'g}����i��}\i}�odL[O�Bط1�ǈ�|�Q�h����bb�e��|�:	�%��߭�6��ံ��_%�y^�Ɋ	��LU�8w�ܱo�c���b��,zǱ�"�K��\�.,m���%ks�S���]�j$��rF$���e����P�vY��W��K�{�m���ԥ�e�f ѕ�)^ҥ�JF����$�2g�w13��H�����Зe�%���M�b?��o�$�E�'I��fve�w�*�\��c���e/�w��Y�w���1R��Z|#��ڧ�F �;QN��!)�f&���[}@�W��3חb���8RlBIz�,O�J�I��W�oy�G8�A��ƿ���o��$y��w�g�9姻��E��M���10��@Y.T}3�a�fQ�����{�mx��P}��z(�GJ;���
�k��"��>��z�h�#�����D�s�Q��V�gu�q�Ez��+B�q�'w>&�,�R���~qt
����,�o�,�����a���#@i��ˀ���&��� �6��V��2�tK"��HҪ�A�J��׃6ح(b��n�-kg�k�M,]��Ĩ�m��ޖF�����-ߵ������y:���@�uAs�q��
;���~X��=d�ټ�3��C�;gJ������Q�� p�G���F��1�EL~�!�n�����ĵ%�KK�A�������w�GdX�� P^U�<uq����#��6�̟tAC�~`,~��X4�h�g�ʓ�ӣ��[;�PU:/��H�bA�<��mw/�h��O��}�;�,*��f�%��@�/������,\;�{:�:��XH�)���u��EK)U��!0���(ӕ���H������t�9��-�l=z�����z�xќ"��k���#��+D8��V�Pp�0)Z*�Up�tZ@�� ��zzjE�	ͧ�gY�y3�yuz��<���5lk=r�NX�U��{��� {r!xH,M��-{f�	�#��p=��S��3�
����e}L4?89�k�h)sU.�?)8d�Q�j�+g������o�(�]-�skw�N6}�d�gv�H�R)��/��]I�n2�ϖc�8=tW��e�v*N�/ ������R�
f����T_\�!�;~I7t4�?y�YMݻ�[đ%��wG�� O	m��""��M�����/�F>��
a��̙�F����Gر���K�"G����g�K����G:}��3]�����$��y�|U�����Gѡ��v�(eWE�4�!��[�@����h_y�nk�_ő˲����<¥��-i�-�JGIh!?%BA���|:1�9�*׳b��|7q��G){��Y#�:�x���pV��|0#�����W�3�w�~�-w��5����L�!2��K*1���������@	����W��=�x�Z,����Ad���aI>5t��=<s���hs�,����	�����:��r�d���@/�ݗ�W̢=P|�0k���	?i�mÕE5��9��;�v�.����3 �x��-�>A3����H�߯��T'ՙ�|Q���v ���V�	})����,.��r��k��z�7������4�4���@2d�9�A�EB� �o8d���d V9���AH��.~5+�F<����� i_��s=ɲP��� v�uh0}@t���[����!����М���ط�P�S�썝i�����龝��4�B�Y៛�g��"�X��|	�f�}��N��F�{�W9��g7���Y�t����r.�bq.A�cV�V46s��x��C-8I^p`� 4�z�:��>�Μ��z2X<w��6��%]$���e��y�,��+����C�.�#��8"��υ���ۋ
�>݋N�Q[�
����e�
����� �x�Gµ^��vt9��}O �4r�m����Os�����	�\��io#��>���?�H#a`���x������\�4Y
�F��(k8��r��܄f^�R��7��Lzo��/�o`����Tq���/�����
)MQJ�=�����صh�4��{>+�i��?�M�Q�����K�7X�
�P�$�h�勪�����7�@�q��׷SY�ԡ�䤷\Hp���,�yL��r殪|��Ǐy��>~���R�"w�H�2!_�X��)�ˍDlPvP����ac���|_PFj}�r�j����t�QD�th���̚%�>�z�N�A��|�k=�\g�Ь�L��a�vÕ`�A���?
��&k{�B5�b�
O�B;n���'�H\�f�{T�M��p+��RR	34u��$M�s�?�y��8{���*8m��x��(�Z1�:Zz�9Bv:�=����[ڠ���^��fi�"�Sg�T�T��7*<Y�]W������J�K/{>���t0h�[n�l*VLh���K�w�� 'QFr���d�@2�Y;Ʀ��*��x�0�|�hԣ0�G�q�����X��Vm�G����������Q_�jŮ_+�-8�n+%w�}�jW�c�pb�c��l�޸'de�4����գ��W�@�N�-��`uP-�_b���a
C�L2��12�dī�)�S��Y���p����C+6tVl�Nj%�c�P�״�nCXQ���6H���i���.�����[��1q���#M닞rb�����)ð����cJ'fu��[��.(�T#1�&���@�D�PD��]�`��	����),3H��0��C�(����i�7d�܀�l�}�(a��.=_�U�F��.�Og����
��� I�%�?c�0�!��QjՂY�')E�P�c�z@�?�W��b�<��sb��<~��2!e"޵7Q{�.�l��ظ3��R�p�;����d3���dڨ����<V'��|��/������܇�n�8uS]_[��+���~mXo'�r��)]	���va�1"]���J��:e�����㩞,��
�֨���p�i%-��� �Y5OR�� d��@
Ea������b�#������~�4�F�e=�_U��'\�>� ��VT)�Wгu��q[��E�����S+��H#WX{��Zn���2�,i'F��1���5�kFO����rp�E��}�#Gx�����m�pCݧd�K�Ab �D����$�N��{���F����y���+W��t�w���*�g����iK�y���V��饦$ ���}�'j�YuQ�[>��F�Ao,>��1�~�KC!�y��f�<kդ��qA3��l�۪���VR��q$�E s�&�B2?�BT{���>N����	���E(^!c~4#�bo銯�S�(� ���Q7^��ggx^���^��o7���3�]Ұ	90�:�<���?PK?3  c w^S�S���'  � H          ��    d5d9210ef49c6780016536b0863cc50f6de03f73e70c2af46cc3cff0e2bf9353.unknown�  AE PK      �   �'   